
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_registerfile_generic_n_bit32_data_bit64 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_registerfile_generic_n_bit32_data_bit64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerfile_generic_n_bit32_data_bit64.all;

entity registerfile_generic_n_bit32_data_bit64 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end registerfile_generic_n_bit32_data_bit64;

architecture SYN_behav of registerfile_generic_n_bit32_data_bit64 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, OUT1_59_port,
      OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, OUT1_54_port, 
      OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, OUT1_49_port, 
      OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, OUT1_44_port, 
      OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, OUT1_39_port, 
      OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, OUT1_34_port, 
      OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, OUT1_29_port, 
      OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, 
      OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, 
      OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, 
      OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, 
      OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, 
      OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, OUT2_63_port, 
      OUT2_62_port, OUT2_61_port, OUT2_60_port, OUT2_59_port, OUT2_58_port, 
      OUT2_57_port, OUT2_56_port, OUT2_55_port, OUT2_54_port, OUT2_53_port, 
      OUT2_52_port, OUT2_51_port, OUT2_50_port, OUT2_49_port, OUT2_48_port, 
      OUT2_47_port, OUT2_46_port, OUT2_45_port, OUT2_44_port, OUT2_43_port, 
      OUT2_42_port, OUT2_41_port, OUT2_40_port, OUT2_39_port, OUT2_38_port, 
      OUT2_37_port, OUT2_36_port, OUT2_35_port, OUT2_34_port, OUT2_33_port, 
      OUT2_32_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port, n4159, n4160, n4161, n4162, n4163,
      n4164, n4165, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
      n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, 
      n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, 
      n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, 
      n4265, n4266, n4267, n4268, n5311, n5312, n5313, n5314, n5315, n5316, 
      n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, 
      n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, 
      n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, 
      n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, 
      n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, 
      n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, 
      n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, 
      n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, 
      n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, 
      n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, 
      n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, 
      n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, 
      n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, 
      n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, 
      n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, 
      n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, 
      n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, 
      n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, 
      n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, 
      n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, 
      n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, 
      n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, 
      n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, 
      n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, 
      n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, 
      n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, 
      n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, 
      n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, 
      n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, 
      n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, 
      n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, 
      n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, 
      n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, 
      n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, 
      n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, 
      n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, 
      n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, 
      n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, 
      n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, 
      n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, 
      n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, 
      n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, 
      n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, 
      n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, 
      n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, 
      n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, 
      n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, 
      n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, 
      n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, 
      n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, 
      n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, 
      n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, 
      n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, 
      n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, 
      n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, 
      n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, 
      n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, 
      n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, 
      n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, 
      n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, 
      n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, 
      n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, 
      n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, 
      n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, 
      n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, 
      n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, 
      n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, 
      n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, 
      n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, 
      n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, 
      n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, 
      n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, 
      n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, 
      n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, 
      n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, 
      n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, 
      n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, 
      n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, 
      n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, 
      n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, 
      n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, 
      n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, 
      n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, 
      n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, 
      n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, 
      n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, 
      n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, 
      n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, 
      n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, 
      n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, 
      n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, 
      n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, 
      n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, 
      n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, 
      n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, 
      n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, 
      n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, 
      n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, 
      n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, 
      n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, 
      n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, 
      n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, 
      n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, 
      n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, 
      n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, 
      n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, 
      n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, 
      n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, 
      n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, 
      n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, 
      n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, 
      n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, 
      n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, 
      n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, 
      n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, 
      n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, 
      n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, 
      n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, 
      n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, 
      n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, 
      n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, 
      n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, 
      n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, 
      n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, 
      n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, 
      n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, 
      n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, 
      n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, 
      n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, 
      n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, 
      n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, 
      n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, 
      n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, 
      n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, 
      n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, 
      n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, 
      n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, 
      n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, 
      n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, 
      n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, 
      n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, 
      n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, 
      n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, 
      n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, 
      n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, 
      n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, 
      n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, 
      n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, 
      n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, 
      n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, 
      n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, 
      n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, 
      n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, 
      n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, 
      n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, 
      n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, 
      n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, 
      n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, 
      n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, 
      n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, 
      n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, 
      n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, 
      n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, 
      n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, 
      n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, 
      n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, 
      n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, 
      n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, 
      n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, 
      n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, 
      n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, 
      n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, 
      n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, 
      n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, 
      n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, 
      n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, 
      n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, 
      n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, 
      n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, 
      n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, 
      n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, 
      n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, 
      n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, 
      n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, 
      n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, 
      n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, 
      n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, 
      n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, 
      n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, 
      n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, 
      n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, 
      n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, 
      n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, 
      n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, 
      n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, 
      n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, 
      n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, 
      n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, 
      n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, 
      n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, 
      n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, 
      n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, 
      n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, 
      n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, 
      n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, 
      n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, 
      n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, 
      n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, 
      n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, 
      n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, 
      n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, 
      n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, 
      n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, 
      n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, 
      n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, 
      n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, 
      n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, 
      n89493, n89496, n89498, n89500, n89965, n89967, n89968, n89969, n90031, 
      n90033, n90034, n90035, n90036, n90037, n90038, n90039, n90040, n90041, 
      n90042, n90043, n90044, n90045, n90046, n90047, n90048, n90049, n90050, 
      n90051, n90052, n90053, n90054, n90055, n90056, n90057, n90058, n90059, 
      n90060, n90061, n90062, n90063, n90064, n90065, n90066, n90067, n90068, 
      n90069, n90070, n90071, n90072, n90073, n90074, n90075, n90076, n90077, 
      n90078, n90079, n90080, n90081, n90082, n90083, n90084, n90085, n90086, 
      n90087, n90088, n90089, n90090, n90091, n90092, n90093, n90094, n90095, 
      n90306, n90308, n90309, n90310, n90311, n90312, n90313, n90314, n90315, 
      n90316, n90317, n90318, n90319, n90320, n90321, n90322, n90323, n90324, 
      n90325, n90326, n90327, n90328, n90329, n90330, n90331, n90332, n90333, 
      n90334, n90335, n90336, n90337, n90338, n90339, n90340, n90341, n90342, 
      n90343, n90344, n90345, n90346, n90347, n90348, n90349, n90350, n90351, 
      n90352, n90353, n90354, n90355, n90356, n90357, n90358, n90359, n90360, 
      n90361, n90362, n90363, n90364, n90365, n90366, n90367, n90368, n90369, 
      n90370, n90373, n90375, n90376, n90377, n90378, n90379, n90380, n90381, 
      n90382, n90383, n90384, n90385, n90386, n90387, n90388, n90389, n90390, 
      n90391, n90392, n90393, n90394, n90395, n90396, n90397, n90398, n90399, 
      n90400, n90401, n90402, n90403, n90404, n90405, n90406, n90407, n90408, 
      n90409, n90410, n90411, n90412, n90413, n90414, n90415, n90416, n90417, 
      n90418, n90419, n90420, n90421, n90422, n90423, n90424, n90425, n90426, 
      n90427, n90428, n90429, n90430, n90431, n90432, n90433, n90434, n90435, 
      n90436, n90437, n90512, n90514, n90515, n90516, n90517, n90518, n90519, 
      n90520, n90521, n90522, n90523, n90524, n90525, n90526, n90527, n90528, 
      n90529, n90530, n90531, n90532, n90533, n90534, n90535, n90536, n90537, 
      n90538, n90539, n90540, n90541, n90542, n90543, n90544, n90545, n90546, 
      n90547, n90548, n90549, n90550, n90551, n90552, n90553, n90554, n90555, 
      n90556, n90557, n90711, n90713, n90714, n90715, n90716, n90717, n90718, 
      n90719, n90720, n90721, n90722, n90723, n90724, n90725, n90726, n90727, 
      n90728, n90729, n90730, n90731, n90732, n90733, n90734, n90735, n90736, 
      n90737, n90738, n90739, n90740, n90741, n90742, n90743, n90744, n90745, 
      n90746, n90747, n90748, n90749, n90750, n90751, n90752, n90753, n90754, 
      n90755, n90756, n90757, n90758, n90759, n90760, n90761, n90762, n90763, 
      n90764, n90765, n90766, n90767, n90768, n90769, n90770, n90771, n90772, 
      n90773, n90774, n90775, n94636, n94637, n94638, n94639, n95429, n95430, 
      n95431, n95432, n95433, n95434, n95435, n95436, n95437, n95438, n95439, 
      n95440, n95441, n95442, n95443, n95444, n95445, n95446, n95447, n95448, 
      n95449, n95450, n95451, n95452, n95453, n95454, n95455, n95456, n95457, 
      n95458, n95459, n95460, n95461, n95462, n95463, n95464, n95465, n95466, 
      n95467, n95468, n95469, n95470, n95471, n95472, n95473, n95474, n95475, 
      n95476, n95477, n95478, n95479, n95480, n95481, n95482, n95483, n95484, 
      n95485, n95486, n95487, n95488, n95525, n95526, n95527, n95528, n98523, 
      n98524, n98525, n98526, n98527, n98528, n98529, n98530, n98531, n98532, 
      n98533, n98534, n98535, n98536, n98537, n98538, n98539, n98540, n98541, 
      n98542, n98543, n98544, n98545, n98546, n98547, n98548, n98549, n98550, 
      n98551, n98552, n98553, n98554, n98555, n98556, n98557, n98558, n98559, 
      n98560, n98561, n98562, n98563, n98564, n98565, n98566, n98567, n98568, 
      n98569, n98570, n98571, n98572, n98573, n98574, n98575, n98576, n98577, 
      n98578, n98579, n98580, n98581, n98582, n98586, n98587, n98588, n98589, 
      n98590, n98591, n98592, n98593, n98594, n98595, n98596, n98597, n98598, 
      n98599, n98600, n98601, n98602, n98603, n98604, n98605, n98606, n98607, 
      n98608, n98609, n98610, n98611, n98612, n98613, n98614, n98615, n98616, 
      n98617, n98618, n98619, n98620, n98621, n98622, n98623, n98624, n98625, 
      n98626, n98627, n98628, n98629, n98630, n98631, n98632, n98633, n98634, 
      n98635, n98636, n98637, n98638, n98639, n98640, n98641, n98642, n98643, 
      n98644, n98645, n98648, n98650, n98651, n98652, n98653, n98654, n98655, 
      n98656, n98657, n98658, n98659, n98660, n98661, n98662, n98663, n98664, 
      n98665, n98666, n98667, n98668, n98669, n98670, n98671, n98672, n98673, 
      n98674, n98675, n98676, n98677, n98678, n98679, n98680, n98681, n98682, 
      n98683, n98684, n98685, n98686, n98687, n98688, n98689, n98690, n98691, 
      n98692, n98693, n98694, n98695, n98696, n98697, n98698, n98699, n98700, 
      n98701, n98702, n98703, n98704, n98705, n98706, n98707, n98708, n98709, 
      n98710, n98711, n98712, n98714, n98716, n98717, n98718, n98719, n98720, 
      n98721, n98722, n98723, n98724, n98725, n98726, n98727, n98728, n98729, 
      n98730, n98731, n98732, n98733, n98734, n98735, n98736, n98737, n98738, 
      n98739, n98740, n98741, n98742, n98743, n98744, n98745, n98746, n98747, 
      n98748, n98749, n98750, n98751, n98752, n98753, n98754, n98755, n98756, 
      n98757, n98758, n98759, n98760, n98761, n98762, n98763, n98764, n98765, 
      n98766, n98767, n98768, n98769, n98770, n98771, n98772, n98773, n98774, 
      n98775, n98776, n98777, n98778, n98848, n98849, n98850, n98851, n98852, 
      n98853, n98854, n98855, n98856, n98857, n98858, n98859, n98860, n98861, 
      n98862, n98863, n98864, n98865, n98866, n98867, n98868, n98869, n98870, 
      n98871, n98872, n98873, n98874, n98875, n98876, n98877, n98878, n98879, 
      n98880, n98881, n98882, n98883, n98884, n98885, n98886, n98887, n98888, 
      n98889, n98890, n98891, n98892, n98893, n98894, n98895, n98896, n98897, 
      n98898, n98899, n98900, n98901, n98902, n98903, n98904, n98905, n98906, 
      n98907, n98986, n98987, n98988, n98989, n98990, n98991, n98992, n98993, 
      n98994, n98995, n98996, n98997, n98998, n98999, n99000, n99001, n99002, 
      n99003, n99004, n99005, n99006, n99007, n99008, n99009, n99010, n99011, 
      n99012, n99013, n99014, n99015, n99016, n99017, n99018, n99019, n99020, 
      n99021, n99022, n99023, n99024, n99025, n99026, n99027, n99028, n99029, 
      n99030, n99031, n99032, n99033, n99034, n99035, n99036, n99037, n99038, 
      n99039, n99040, n99041, n99042, n99043, n99044, n99045, n99047, n99049, 
      n99050, n99051, n99052, n99053, n99054, n99055, n99056, n99057, n99058, 
      n99059, n99060, n99061, n99062, n99063, n99064, n99065, n99066, n99067, 
      n99068, n99069, n99070, n99071, n99072, n99073, n99074, n99075, n99076, 
      n99077, n99078, n99079, n99080, n99081, n99082, n99083, n99084, n99085, 
      n99086, n99087, n99088, n99089, n99090, n99091, n99092, n99093, n99094, 
      n99095, n99096, n99097, n99098, n99099, n99100, n99101, n99102, n99103, 
      n99104, n99105, n99106, n99107, n99108, n99109, n99110, n99111, n99113, 
      n99115, n99116, n99117, n99118, n99119, n99120, n99121, n99122, n99123, 
      n99124, n99125, n99126, n99127, n99128, n99129, n99130, n99131, n99132, 
      n99133, n99134, n99135, n99136, n99137, n99138, n99139, n99140, n99141, 
      n99142, n99143, n99144, n99145, n99146, n99147, n99148, n99149, n99150, 
      n99151, n99152, n99153, n99154, n99155, n99156, n99157, n99158, n99159, 
      n99160, n99161, n99162, n99163, n99164, n99165, n99166, n99167, n99168, 
      n99169, n99170, n99171, n99172, n99173, n99174, n99175, n99176, n99177, 
      n99179, n99181, n99182, n99183, n99184, n99185, n99186, n99187, n99188, 
      n99189, n99190, n99191, n99192, n99193, n99194, n99195, n99196, n99197, 
      n99198, n99199, n99200, n99201, n99202, n99203, n99204, n99205, n99206, 
      n99207, n99208, n99209, n99210, n99211, n99212, n99213, n99214, n99215, 
      n99216, n99217, n99218, n99219, n99220, n99221, n99222, n99223, n99224, 
      n99225, n99226, n99227, n99228, n99229, n99230, n99231, n99232, n99233, 
      n99234, n99235, n99236, n99237, n99238, n99239, n99240, n99241, n99242, 
      n99243, n99245, n99247, n99248, n99249, n99250, n99251, n99252, n99253, 
      n99254, n99255, n99256, n99257, n99258, n99259, n99260, n99261, n99262, 
      n99263, n99264, n99265, n99266, n99267, n99268, n99269, n99270, n99271, 
      n99272, n99273, n99274, n99275, n99276, n99277, n99278, n99279, n99280, 
      n99281, n99282, n99283, n99284, n99285, n99286, n99287, n99288, n99289, 
      n99290, n99291, n99292, n99293, n99294, n99295, n99296, n99297, n99298, 
      n99299, n99300, n99301, n99302, n99303, n99304, n99305, n99306, n99307, 
      n99308, n99309, n99311, n99313, n99314, n99315, n99316, n99317, n99318, 
      n99319, n99320, n99321, n99322, n99323, n99324, n99325, n99326, n99327, 
      n99328, n99329, n99330, n99331, n99332, n99333, n99334, n99335, n99336, 
      n99337, n99338, n99339, n99340, n99341, n99342, n99343, n99344, n99345, 
      n99346, n99347, n99348, n99349, n99350, n99351, n99352, n99353, n99354, 
      n99355, n99356, n99357, n99358, n99359, n99360, n99361, n99362, n99363, 
      n99364, n99365, n99366, n99367, n99368, n99369, n99370, n99371, n99372, 
      n99373, n99374, n99375, n99446, n99448, n99449, n99450, n99451, n99452, 
      n99453, n99454, n99455, n99456, n99457, n99458, n99459, n99460, n99461, 
      n99462, n99463, n99464, n99465, n99466, n99467, n99468, n99469, n99470, 
      n99471, n99472, n99473, n99474, n99475, n99476, n99477, n99478, n99479, 
      n99480, n99481, n99482, n99483, n99484, n99485, n99486, n99487, n99488, 
      n99489, n99490, n99491, n99492, n99493, n99494, n99495, n99496, n99497, 
      n99498, n99499, n99500, n99501, n99502, n99503, n99504, n99505, n99506, 
      n99507, n99508, n99509, n99510, n99580, n99582, n99583, n99584, n99585, 
      n99586, n99587, n99588, n99589, n99590, n99591, n99592, n99593, n99594, 
      n99595, n99596, n99597, n99598, n99599, n99600, n99601, n99602, n99603, 
      n99604, n99605, n99606, n99607, n99608, n99609, n99610, n99611, n99612, 
      n99613, n99614, n99615, n99616, n99617, n99618, n99619, n99620, n99621, 
      n99622, n99623, n99624, n99625, n99626, n99627, n99628, n99629, n99630, 
      n99631, n99632, n99633, n99634, n99635, n99636, n99637, n99638, n99639, 
      n99640, n99641, n99642, n99643, n99644, n99716, n99718, n99719, n99720, 
      n99721, n99722, n99723, n99724, n99725, n99726, n99727, n99728, n99729, 
      n99730, n99731, n99732, n99733, n99734, n99735, n99736, n99737, n99738, 
      n99739, n99740, n99741, n99742, n99743, n99744, n99745, n99746, n99747, 
      n99748, n99749, n99750, n99751, n99752, n99753, n99754, n99755, n99756, 
      n99757, n99758, n99759, n99760, n99761, n99762, n99763, n99764, n99765, 
      n99766, n99767, n99768, n99769, n99770, n99771, n99772, n99773, n99774, 
      n99775, n99776, n99777, n99778, n99779, n99780, n99914, n99916, n99917, 
      n99918, n99919, n99920, n99921, n99922, n99923, n99924, n99925, n99926, 
      n99927, n99928, n99929, n99930, n99931, n99932, n99933, n99934, n99935, 
      n99936, n99937, n99938, n99939, n99940, n99941, n99942, n99943, n99944, 
      n99945, n99946, n99947, n99948, n99949, n99950, n99951, n99952, n99953, 
      n99954, n99955, n99956, n99957, n99958, n99959, n99960, n99961, n99962, 
      n99963, n99964, n99965, n99966, n99967, n99968, n99969, n99970, n99971, 
      n99972, n99973, n99974, n99975, n99976, n99977, n99978, n103034, n103035,
      n103036, n103037, n103038, n103039, n103040, n103041, n103042, n103043, 
      n103044, n103045, n103046, n103047, n103048, n103049, n103050, n103051, 
      n103552, n103553, n103554, n103555, n103556, n103557, n103558, n103559, 
      n103560, n103561, n103562, n103563, n103564, n103565, n103566, n103567, 
      n103568, n103569, n103570, n103571, n103572, n103573, n103574, n103575, 
      n103576, n103577, n103578, n103579, n103580, n103581, n103582, n103583, 
      n103584, n103585, n103586, n103587, n103588, n103589, n103590, n103591, 
      n103592, n103593, n103594, n103595, n103596, n103597, n103598, n103599, 
      n103600, n103601, n103602, n103603, n103604, n103605, n103606, n103607, 
      n103608, n103609, n103610, n103611, n103736, n103737, n103738, n103739, 
      n109895, n109896, n109897, n109898, n109903, n109904, n109905, n109906, 
      n109979, n109980, n109981, n109982, n109983, n109984, n109985, n109986, 
      n109987, n109988, n109989, n109990, n109991, n109992, n109993, n109994, 
      n109995, n109996, n109997, n110107, n110108, n110109, n110110, n110171, 
      n110172, n110173, n110174, n110175, n110176, n110177, n110178, n110179, 
      n110180, n110181, n110182, n110183, n110184, n110185, n110186, n110187, 
      n110188, n110189, n110190, n110191, n110192, n110193, n110194, n110195, 
      n110196, n110197, n110198, n110199, n110200, n110201, n110202, n110203, 
      n110204, n110205, n110206, n110207, n110208, n110209, n110210, n110211, 
      n110212, n110213, n110214, n110215, n110216, n110217, n110218, n110219, 
      n110220, n110221, n110222, n110223, n110224, n110225, n110226, n110227, 
      n110228, n110229, n110230, n110231, n110232, n110233, n110234, n110363, 
      n110364, n110365, n110366, n110431, n110432, n110433, n110434, n110435, 
      n110436, n110437, n110438, n110439, n110440, n110441, n110442, n110443, 
      n110444, n110445, n110446, n110447, n110448, n110449, n110450, n110451, 
      n110452, n110453, n110454, n110455, n110456, n110457, n110458, n110459, 
      n110460, n110461, n110462, n110463, n110464, n110465, n110466, n110467, 
      n110468, n110469, n110470, n110471, n110472, n110473, n110474, n110475, 
      n110476, n110477, n110478, n110479, n110480, n110481, n110482, n110483, 
      n110484, n110485, n110486, n110487, n110488, n110489, n110490, n110491, 
      n110492, n110493, n110494, n110495, n110496, n110497, n110498, n110499, 
      n110500, n110501, n110502, n110503, n110504, n110505, n110506, n110507, 
      n110508, n110509, n110510, n110511, n110512, n110513, n110514, n110515, 
      n110516, n110517, n110518, n110519, n110520, n110521, n110522, n110523, 
      n110524, n110525, n110526, n110527, n110528, n110529, n110530, n110531, 
      n110532, n110533, n110534, n110535, n110536, n110537, n110538, n110539, 
      n110540, n110541, n110542, n110543, n110544, n110545, n110546, n110547, 
      n110548, n110549, n110550, n110551, n110552, n110553, n110554, n110555, 
      n110556, n110557, n110558, n110559, n110560, n110561, n110562, n110563, 
      n110564, n110565, n110566, n110567, n110568, n110569, n110570, n110571, 
      n110572, n110573, n110574, n110575, n110576, n110577, n110578, n110579, 
      n110580, n110581, n110582, n110583, n110584, n110585, n110586, n110587, 
      n110588, n110589, n110590, n110591, n110592, n110593, n110594, n110595, 
      n110596, n110597, n110598, n110599, n110600, n110601, n110602, n110603, 
      n110604, n110605, n110606, n110607, n110608, n110609, n110610, n110611, 
      n110612, n110613, n110614, n110615, n110616, n110617, n110618, n110619, 
      n110620, n110621, n110622, n110811, n110812, n110813, n110814, n110815, 
      n110816, n110817, n110818, n110819, n110820, n110821, n110822, n110823, 
      n110824, n110825, n110826, n110827, n110828, n110829, n110830, n110831, 
      n110832, n110833, n110834, n110835, n110836, n110837, n110838, n110839, 
      n110840, n110841, n110842, n110843, n110844, n110845, n110846, n110847, 
      n110848, n110849, n110850, n110851, n110852, n110853, n110854, n110855, 
      n110856, n110857, n110858, n110859, n110860, n110861, n110862, n110863, 
      n110864, n110865, n110866, n110867, n110868, n110869, n110870, n110871, 
      n110872, n110873, n110874, n110939, n110940, n110941, n110942, n110943, 
      n110944, n110945, n110946, n110947, n110948, n110949, n110950, n110951, 
      n110952, n110953, n110954, n110955, n110956, n110957, n110996, n110997, 
      n110998, n110999, n111000, n111001, n111002, n111003, n111004, n111005, 
      n111006, n111007, n111008, n111009, n111010, n111011, n111012, n111013, 
      n111014, n111015, n111016, n111017, n111018, n111019, n111020, n111021, 
      n111022, n111023, n111024, n111025, n111026, n111027, n111028, n111029, 
      n111030, n111031, n111032, n111033, n111034, n111035, n111036, n111037, 
      n111038, n111039, n111040, n111041, n111042, n111043, n111044, n111045, 
      n111046, n111047, n111048, n113766, n113767, n113768, n113769, n113770, 
      n113771, n113772, n113773, n113774, n113775, n113776, n113777, n113778, 
      n113779, n113780, n113781, n113782, n113783, n113784, n113785, n113786, 
      n113787, n113788, n113789, n113790, n113791, n113792, n113793, n113794, 
      n113795, n113796, n113797, n113798, n113799, n113800, n113801, n113802, 
      n113803, n113804, n113805, n113806, n113807, n113808, n113809, n113810, 
      n113811, n113812, n113813, n113814, n113815, n113816, n113817, n113818, 
      n113819, n113820, n113821, n113822, n113823, n113824, n113825, n113826, 
      n113827, n113828, n113829, n113830, n113831, n113832, n113833, n113834, 
      n113835, n113836, n113837, n113838, n113839, n113840, n113841, n113842, 
      n113843, n113844, n113845, n113846, n113847, n113848, n113849, n113850, 
      n113851, n113852, n113853, n113854, n113855, n113856, n113857, n113858, 
      n113859, n113860, n113861, n113862, n113863, n113864, n113865, n113866, 
      n113867, n113868, n113869, n113870, n113871, n113872, n113873, n113874, 
      n113875, n113876, n113877, n113878, n113879, n113880, n113881, n113882, 
      n113883, n113884, n113885, n113886, n113887, n113888, n113889, n113890, 
      n113891, n113892, n113893, n113894, n113895, n113896, n113897, n113898, 
      n113899, n113900, n113901, n113902, n113903, n113904, n113905, n113906, 
      n113907, n113908, n113909, n113910, n113911, n113912, n113913, n113914, 
      n113915, n113916, n113917, n113918, n113919, n113920, n113921, n113922, 
      n113923, n113924, n113925, n113926, n113927, n113928, n113929, n113930, 
      n113931, n113932, n113933, n113934, n113935, n113936, n113937, n113938, 
      n113939, n113940, n113941, n113942, n113943, n113944, n113945, n113946, 
      n113947, n113948, n113949, n113950, n113951, n113952, n113953, n113954, 
      n113955, n113956, n113957, n113958, n113959, n113960, n113961, n113962, 
      n113963, n113964, n113965, n113966, n113967, n113968, n113969, n113970, 
      n113971, n113972, n113973, n113974, n113975, n113976, n113977, n113978, 
      n113979, n113980, n113981, n113982, n113983, n113984, n113985, n113986, 
      n113987, n113988, n113989, n113990, n113991, n113992, n113993, n113994, 
      n113995, n113996, n113997, n113998, n113999, n114000, n114001, n114002, 
      n114003, n114004, n114005, n114006, n114007, n114008, n114009, n114010, 
      n114011, n114012, n114013, n114014, n114015, n114016, n114017, n114018, 
      n114019, n114020, n114021, n114022, n114023, n114024, n114025, n114026, 
      n114027, n114028, n114029, n114030, n114031, n114032, n114033, n114034, 
      n114035, n114036, n114037, n114038, n114039, n114040, n114041, n114042, 
      n114043, n114044, n114045, n114046, n114047, n114048, n114049, n114050, 
      n114051, n114052, n114053, n114054, n114055, n114056, n114057, n114058, 
      n114059, n114060, n114061, n114062, n114063, n114064, n114065, n114066, 
      n114067, n114068, n114069, n114070, n114071, n114072, n114073, n114074, 
      n114075, n114076, n114077, n114078, n114079, n114080, n114081, n114082, 
      n114083, n114084, n114085, n114086, n114087, n114088, n114089, n114090, 
      n114091, n114092, n114093, n114094, n114095, n114096, n114097, n114098, 
      n114099, n114100, n114101, n114102, n114103, n114104, n114105, n114106, 
      n114107, n114108, n114109, n114110, n114111, n114112, n114113, n114114, 
      n114115, n114116, n114117, n114118, n114119, n114120, n114121, n114122, 
      n114123, n114124, n114125, n114126, n114127, n114128, n114129, n114130, 
      n114131, n114132, n114133, n114134, n114135, n114136, n114137, n114138, 
      n114139, n114140, n114141, n114142, n114143, n114144, n114145, n114146, 
      n114147, n114148, n114149, n114150, n114151, n114152, n114153, n114154, 
      n114155, n114156, n114157, n114158, n114159, n114160, n114161, n114162, 
      n114163, n114164, n114165, n114166, n114167, n114168, n114169, n114170, 
      n114171, n114172, n114173, n114174, n114175, n114176, n114177, n114178, 
      n114179, n114180, n114181, n114182, n114183, n114184, n114185, n114186, 
      n114187, n114188, n114189, n114190, n114191, n114192, n114193, n114194, 
      n114195, n114196, n114197, n114198, n114199, n114200, n114201, n114202, 
      n114203, n114204, n114205, n114206, n114207, n114208, n114209, n114210, 
      n114211, n114212, n114213, n114214, n114215, n114216, n114217, n114218, 
      n114219, n114220, n114221, n114222, n114223, n114224, n114225, n114226, 
      n114227, n114228, n114229, n114230, n114231, n114232, n114233, n114234, 
      n114235, n114236, n114237, n114238, n114239, n114240, n114241, n114242, 
      n114243, n114244, n114245, n114246, n114247, n114248, n114249, n114250, 
      n114251, n114252, n114253, n114254, n114255, n114256, n114257, n114258, 
      n114259, n114260, n114261, n114262, n114263, n114264, n114265, n114266, 
      n114267, n114268, n114269, n114270, n114271, n114272, n114273, n114274, 
      n114275, n114276, n114277, n114278, n114279, n114280, n114281, n114282, 
      n114283, n114284, n114285, n114286, n114287, n114288, n114289, n114290, 
      n114291, n114292, n114293, n114294, n114295, n114296, n114297, n114298, 
      n114299, n114300, n114301, n114302, n114303, n114304, n114305, n114306, 
      n114307, n114308, n114309, n114310, n114311, n114312, n114313, n114314, 
      n114315, n114316, n114317, n114318, n114319, n114320, n114321, n114322, 
      n114323, n114324, n114325, n114326, n114327, n114328, n114329, n114330, 
      n114331, n114332, n114333, n114334, n114335, n114336, n114337, n114338, 
      n114339, n114340, n114341, n114342, n114343, n114344, n114345, n114346, 
      n114347, n114348, n114349, n114350, n114351, n114352, n114353, n114354, 
      n114355, n114356, n114357, n114358, n114359, n114360, n114361, n114362, 
      n114363, n114364, n114365, n114366, n114367, n114368, n114369, n114370, 
      n114371, n114372, n114373, n114374, n114375, n114376, n114377, n114378, 
      n114379, n114380, n114381, n114382, n114383, n114384, n114385, n114386, 
      n114387, n114388, n114389, n114390, n114391, n114392, n114393, n114394, 
      n114395, n114396, n114397, n114398, n114399, n114400, n114401, n114402, 
      n114403, n114404, n114405, n114406, n114407, n114408, n114409, n114410, 
      n114411, n114412, n114413, n114414, n114415, n114416, n114417, n114418, 
      n114419, n114420, n114421, n114422, n114423, n114424, n114425, n114426, 
      n114427, n114428, n114429, n114430, n114431, n114432, n114433, n114434, 
      n114435, n114436, n114437, n114438, n114439, n114440, n114441, n114442, 
      n114443, n114444, n114445, n114446, n114447, n114448, n114449, n114450, 
      n114451, n114452, n114453, n114454, n114455, n114456, n114457, n114458, 
      n114459, n114460, n114461, n114462, n114463, n114464, n114465, n114466, 
      n114467, n114468, n114469, n114470, n114471, n114472, n114473, n114474, 
      n114475, n114476, n114477, n114478, n114479, n114480, n114481, n114482, 
      n114483, n114484, n114485, n114486, n114487, n114488, n114489, n114490, 
      n114491, n114492, n114493, n114494, n114495, n114496, n114497, n114498, 
      n114499, n114500, n114501, n114502, n114503, n114504, n114505, n114506, 
      n114507, n114508, n114509, n114510, n114511, n114512, n114513, n114514, 
      n114515, n114516, n114517, n114518, n114519, n114520, n114521, n114522, 
      n114523, n114524, n114525, n114526, n114527, n114528, n114529, n114530, 
      n114531, n114532, n114533, n114534, n114535, n114536, n114537, n114538, 
      n114539, n114540, n114541, n114542, n114543, n114544, n114545, n114546, 
      n114547, n114548, n114549, n114550, n114551, n114552, n114553, n114554, 
      n114555, n114556, n114557, n114558, n114559, n114560, n114561, n114562, 
      n114563, n114564, n114565, n114566, n114567, n114568, n114569, n114570, 
      n114571, n114572, n114573, n114574, n114575, n114576, n114577, n114578, 
      n114579, n114580, n114581, n114582, n114583, n114584, n114585, n114586, 
      n114587, n114588, n114589, n114590, n114591, n114592, n114593, n114594, 
      n114595, n114596, n114597, n114598, n114599, n114600, n114601, n114602, 
      n114603, n114604, n114605, n114606, n114607, n114608, n114609, n114610, 
      n114611, n114612, n114613, n114614, n114615, n114616, n114617, n114618, 
      n114619, n114620, n114621, n114622, n114623, n114624, n114625, n114626, 
      n114627, n114628, n114629, n114630, n114631, n114632, n114633, n114634, 
      n114635, n114636, n114637, n114638, n114639, n114640, n114641, n114642, 
      n114643, n114644, n114645, n114646, n114647, n114648, n114649, n114650, 
      n114651, n114652, n114653, n114654, n114655, n114656, n114657, n114658, 
      n114659, n114660, n114661, n114662, n114664, n114666, n114667, n114668, 
      n114669, n114670, n114672, n114673, n114674, n114675, n114676, n114678, 
      n114679, n114680, n114681, n114682, n114683, n114684, n114685, n114686, 
      n114687, n114688, n114689, n114690, n114691, n114693, n114695, n114696, 
      n114697, n114698, n114700, n114701, n114702, n114703, n114704, n114705, 
      n114706, n114707, n114708, n114709, n114710, n114711, n114712, n114713, 
      n114714, n114717, n114719, n114721, n114722, n114723, n114724, n114727, 
      n114729, n114730, n114731, n114732, n114733, n114734, n114735, n114736, 
      n114737, n114738, n114739, n114740, n114743, n114745, n114747, n114748, 
      n114749, n114750, n114753, n114755, n114756, n114757, n114758, n114759, 
      n114760, n114761, n114762, n114763, n114764, n114765, n114766, n114769, 
      n114771, n114773, n114774, n114775, n114776, n114779, n114781, n114782, 
      n114783, n114784, n114785, n114786, n114787, n114788, n114789, n114790, 
      n114791, n114793, n114796, n114798, n114801, n114802, n114803, n114804, 
      n114807, n114809, n114810, n114811, n114812, n114813, n114814, n114815, 
      n114816, n114817, n114818, n114819, n114821, n114824, n114826, n114829, 
      n114830, n114831, n114832, n114835, n114837, n114838, n114839, n114840, 
      n114841, n114842, n114843, n114844, n114845, n114846, n114847, n114849, 
      n114852, n114854, n114857, n114858, n114859, n114860, n114863, n114865, 
      n114866, n114867, n114868, n114869, n114870, n114871, n114872, n114873, 
      n114874, n114875, n114877, n114880, n114882, n114885, n114886, n114887, 
      n114888, n114891, n114893, n114894, n114895, n114896, n114897, n114898, 
      n114899, n114900, n114901, n114902, n114903, n114905, n114908, n114910, 
      n114913, n114914, n114915, n114916, n114919, n114921, n114922, n114923, 
      n114924, n114925, n114926, n114927, n114928, n114929, n114930, n114931, 
      n114933, n114936, n114938, n114941, n114942, n114943, n114944, n114947, 
      n114949, n114950, n114951, n114952, n114953, n114954, n114955, n114956, 
      n114957, n114958, n114959, n114961, n114964, n114966, n114969, n114970, 
      n114971, n114972, n114975, n114977, n114978, n114979, n114980, n114981, 
      n114982, n114983, n114984, n114985, n114986, n114987, n114989, n114992, 
      n114994, n114997, n114998, n114999, n115000, n115003, n115005, n115006, 
      n115007, n115008, n115009, n115010, n115011, n115012, n115013, n115014, 
      n115015, n115017, n115020, n115022, n115025, n115026, n115027, n115028, 
      n115031, n115033, n115034, n115035, n115036, n115037, n115038, n115039, 
      n115040, n115041, n115042, n115043, n115045, n115048, n115050, n115053, 
      n115054, n115055, n115056, n115059, n115061, n115062, n115063, n115064, 
      n115065, n115066, n115067, n115068, n115069, n115070, n115071, n115073, 
      n115076, n115078, n115081, n115082, n115083, n115084, n115087, n115089, 
      n115090, n115091, n115092, n115093, n115094, n115095, n115096, n115097, 
      n115098, n115099, n115101, n115104, n115106, n115109, n115110, n115111, 
      n115112, n115115, n115117, n115118, n115119, n115120, n115121, n115122, 
      n115123, n115124, n115125, n115126, n115127, n115129, n115132, n115134, 
      n115137, n115138, n115139, n115140, n115143, n115145, n115146, n115147, 
      n115148, n115149, n115150, n115151, n115152, n115153, n115154, n115155, 
      n115157, n115160, n115162, n115165, n115166, n115167, n115168, n115171, 
      n115173, n115174, n115175, n115176, n115177, n115178, n115179, n115180, 
      n115181, n115182, n115183, n115185, n115188, n115190, n115193, n115194, 
      n115195, n115196, n115199, n115201, n115202, n115203, n115204, n115205, 
      n115206, n115207, n115208, n115209, n115210, n115211, n115213, n115216, 
      n115218, n115221, n115222, n115223, n115224, n115227, n115229, n115230, 
      n115231, n115232, n115233, n115234, n115235, n115236, n115237, n115238, 
      n115239, n115241, n115244, n115246, n115249, n115250, n115251, n115252, 
      n115255, n115257, n115258, n115259, n115260, n115261, n115262, n115263, 
      n115264, n115265, n115266, n115267, n115269, n115272, n115274, n115277, 
      n115278, n115279, n115280, n115283, n115285, n115286, n115287, n115288, 
      n115289, n115290, n115291, n115292, n115293, n115294, n115295, n115297, 
      n115300, n115302, n115305, n115306, n115307, n115308, n115311, n115313, 
      n115314, n115315, n115316, n115317, n115318, n115319, n115320, n115321, 
      n115322, n115323, n115325, n115328, n115330, n115333, n115334, n115335, 
      n115336, n115339, n115341, n115342, n115343, n115344, n115345, n115346, 
      n115347, n115348, n115349, n115350, n115351, n115353, n115356, n115358, 
      n115361, n115362, n115363, n115364, n115367, n115369, n115370, n115371, 
      n115372, n115373, n115374, n115375, n115376, n115377, n115378, n115379, 
      n115381, n115384, n115386, n115389, n115390, n115391, n115392, n115395, 
      n115397, n115398, n115399, n115400, n115401, n115402, n115403, n115404, 
      n115405, n115406, n115407, n115409, n115412, n115414, n115417, n115418, 
      n115419, n115420, n115423, n115425, n115426, n115427, n115428, n115429, 
      n115430, n115431, n115432, n115433, n115434, n115435, n115437, n115440, 
      n115442, n115445, n115446, n115447, n115448, n115451, n115453, n115454, 
      n115455, n115456, n115457, n115458, n115459, n115460, n115461, n115462, 
      n115463, n115465, n115468, n115470, n115473, n115474, n115475, n115476, 
      n115479, n115481, n115482, n115483, n115484, n115485, n115486, n115487, 
      n115488, n115489, n115490, n115491, n115493, n115496, n115498, n115501, 
      n115502, n115503, n115504, n115507, n115509, n115510, n115511, n115512, 
      n115513, n115514, n115515, n115516, n115517, n115518, n115519, n115521, 
      n115524, n115526, n115529, n115530, n115531, n115532, n115535, n115537, 
      n115538, n115539, n115540, n115541, n115542, n115543, n115544, n115545, 
      n115546, n115547, n115549, n115552, n115554, n115557, n115558, n115559, 
      n115560, n115563, n115565, n115566, n115567, n115568, n115569, n115570, 
      n115571, n115572, n115573, n115574, n115575, n115577, n115580, n115582, 
      n115585, n115586, n115587, n115588, n115591, n115593, n115594, n115595, 
      n115596, n115597, n115598, n115599, n115600, n115601, n115602, n115603, 
      n115605, n115608, n115610, n115613, n115614, n115615, n115616, n115619, 
      n115621, n115622, n115623, n115624, n115625, n115626, n115627, n115628, 
      n115629, n115630, n115631, n115633, n115636, n115638, n115641, n115642, 
      n115643, n115644, n115647, n115649, n115650, n115651, n115652, n115653, 
      n115654, n115655, n115656, n115657, n115658, n115659, n115661, n115664, 
      n115666, n115669, n115670, n115671, n115672, n115675, n115677, n115678, 
      n115679, n115680, n115681, n115682, n115683, n115684, n115685, n115686, 
      n115687, n115689, n115692, n115694, n115697, n115698, n115699, n115700, 
      n115703, n115705, n115706, n115707, n115708, n115709, n115710, n115711, 
      n115712, n115713, n115714, n115715, n115717, n115720, n115722, n115725, 
      n115726, n115727, n115728, n115731, n115733, n115734, n115735, n115736, 
      n115737, n115738, n115739, n115740, n115741, n115742, n115743, n115745, 
      n115748, n115750, n115753, n115754, n115755, n115756, n115759, n115761, 
      n115762, n115763, n115764, n115765, n115766, n115767, n115768, n115769, 
      n115770, n115771, n115773, n115776, n115778, n115781, n115782, n115783, 
      n115784, n115787, n115789, n115790, n115791, n115792, n115793, n115794, 
      n115795, n115796, n115797, n115798, n115799, n115801, n115804, n115806, 
      n115809, n115810, n115811, n115812, n115815, n115817, n115818, n115819, 
      n115820, n115821, n115822, n115823, n115824, n115825, n115826, n115827, 
      n115829, n115832, n115834, n115837, n115838, n115839, n115840, n115843, 
      n115845, n115846, n115847, n115848, n115849, n115850, n115851, n115852, 
      n115853, n115854, n115855, n115857, n115860, n115862, n115865, n115866, 
      n115867, n115868, n115871, n115873, n115874, n115875, n115876, n115877, 
      n115878, n115879, n115880, n115881, n115882, n115883, n115885, n115888, 
      n115890, n115893, n115894, n115895, n115896, n115899, n115901, n115902, 
      n115903, n115904, n115905, n115906, n115907, n115908, n115909, n115910, 
      n115911, n115913, n115916, n115918, n115921, n115922, n115923, n115924, 
      n115927, n115929, n115930, n115931, n115932, n115933, n115934, n115935, 
      n115936, n115937, n115938, n115939, n115941, n115944, n115946, n115949, 
      n115950, n115951, n115952, n115955, n115957, n115958, n115959, n115960, 
      n115961, n115962, n115963, n115964, n115965, n115966, n115967, n115969, 
      n115972, n115974, n115977, n115978, n115979, n115980, n115983, n115985, 
      n115986, n115987, n115988, n115989, n115990, n115991, n115992, n115993, 
      n115994, n115995, n115997, n116000, n116002, n116005, n116006, n116007, 
      n116008, n116011, n116013, n116014, n116015, n116016, n116017, n116018, 
      n116019, n116020, n116021, n116022, n116023, n116025, n116028, n116030, 
      n116033, n116034, n116035, n116036, n116039, n116041, n116042, n116043, 
      n116044, n116045, n116046, n116047, n116048, n116049, n116050, n116051, 
      n116053, n116056, n116058, n116061, n116062, n116063, n116064, n116067, 
      n116069, n116070, n116071, n116072, n116073, n116074, n116075, n116076, 
      n116077, n116078, n116079, n116081, n116084, n116086, n116089, n116090, 
      n116091, n116092, n116095, n116097, n116098, n116099, n116100, n116101, 
      n116102, n116103, n116104, n116105, n116106, n116107, n116109, n116112, 
      n116114, n116117, n116118, n116119, n116120, n116123, n116125, n116126, 
      n116127, n116128, n116129, n116130, n116131, n116132, n116133, n116134, 
      n116135, n116137, n116140, n116142, n116145, n116146, n116147, n116148, 
      n116151, n116153, n116154, n116155, n116156, n116157, n116158, n116159, 
      n116160, n116161, n116162, n116163, n116165, n116168, n116170, n116173, 
      n116174, n116175, n116176, n116179, n116181, n116182, n116183, n116184, 
      n116185, n116186, n116187, n116188, n116189, n116190, n116191, n116193, 
      n116196, n116198, n116201, n116202, n116203, n116204, n116207, n116209, 
      n116210, n116211, n116212, n116213, n116214, n116215, n116216, n116217, 
      n116218, n116219, n116221, n116224, n116226, n116229, n116230, n116231, 
      n116232, n116235, n116237, n116238, n116239, n116240, n116241, n116242, 
      n116243, n116244, n116245, n116246, n116247, n116249, n116252, n116254, 
      n116257, n116258, n116259, n116260, n116263, n116265, n116266, n116267, 
      n116268, n116269, n116270, n116271, n116272, n116273, n116274, n116275, 
      n116277, n116280, n116282, n116285, n116286, n116287, n116288, n116291, 
      n116293, n116294, n116295, n116296, n116297, n116298, n116299, n116300, 
      n116301, n116302, n116303, n116305, n116308, n116310, n116313, n116314, 
      n116315, n116316, n116319, n116321, n116322, n116323, n116324, n116325, 
      n116326, n116327, n116328, n116329, n116330, n116331, n116333, n116336, 
      n116338, n116341, n116342, n116343, n116344, n116347, n116349, n116350, 
      n116351, n116352, n116353, n116354, n116355, n116356, n116357, n116358, 
      n116359, n116361, n116364, n116366, n116369, n116370, n116371, n116372, 
      n116375, n116377, n116378, n116379, n116380, n116381, n116382, n116383, 
      n116384, n116385, n116386, n116387, n116389, n116392, n116394, n116397, 
      n116398, n116399, n116400, n116403, n116405, n116406, n116407, n116408, 
      n116409, n116410, n116411, n116412, n116413, n116414, n116415, n116417, 
      n116420, n116422, n116425, n116426, n116427, n116428, n116431, n116433, 
      n116434, n116435, n116436, n116437, n116438, n116439, n116440, n116441, 
      n116442, n116443, n116445, n116446, n116447, n116448, n116449, n116452, 
      n116453, n116454, n116455, n116457, n116458, n116459, n116460, n116463, 
      n116464, n116465, n116466, n116467, n116468, n116469, n116470, n116471, 
      n116474, n116475, n116477, n116478, n116479, n116480, n116481, n116482, 
      n116483, n116484, n116485, n116486, n116487, n116488, n116489, n116490, 
      n116491, n116492, n116493, n116494, n116495, n116497, n116499, n116500, 
      n116501, n116502, n116503, n116504, n116505, n116506, n116507, n116508, 
      n116509, n116510, n116511, n116512, n116513, n116514, n116515, n116516, 
      n116517, n116518, n116519, n116520, n116521, n116522, n116523, n116525, 
      n116526, n116527, n116528, n116529, n116530, n116531, n116532, n116533, 
      n116534, n116535, n116536, n116537, n116538, n116539, n116540, n116541, 
      n116542, n116545, n116546, n116547, n116548, n116549, n116550, n116552, 
      n116553, n116554, n116555, n116556, n116557, n116558, n116559, n116560, 
      n116561, n116562, n116563, n116566, n116567, n116568, n116569, n116570, 
      n116571, n116573, n116574, n116575, n116576, n116577, n116578, n116579, 
      n116580, n116581, n116582, n116583, n116584, n116587, n116588, n116589, 
      n116590, n116591, n116592, n116594, n116595, n116596, n116597, n116598, 
      n116599, n116600, n116601, n116602, n116603, n116604, n116606, n116609, 
      n116611, n116612, n116613, n116614, n116615, n116617, n116618, n116619, 
      n116620, n116621, n116622, n116623, n116624, n116625, n116626, n116627, 
      n116629, n116632, n116634, n116635, n116636, n116637, n116638, n116640, 
      n116641, n116642, n116643, n116644, n116645, n116646, n116647, n116648, 
      n116649, n116650, n116652, n116655, n116657, n116658, n116659, n116660, 
      n116661, n116663, n116664, n116665, n116666, n116667, n116668, n116669, 
      n116670, n116671, n116672, n116673, n116675, n116678, n116680, n116681, 
      n116682, n116683, n116684, n116686, n116687, n116688, n116689, n116690, 
      n116691, n116692, n116693, n116694, n116695, n116696, n116698, n116701, 
      n116703, n116704, n116705, n116706, n116707, n116709, n116710, n116711, 
      n116712, n116713, n116714, n116715, n116716, n116717, n116718, n116719, 
      n116721, n116724, n116726, n116727, n116728, n116729, n116730, n116732, 
      n116733, n116734, n116735, n116736, n116737, n116738, n116739, n116740, 
      n116741, n116742, n116744, n116747, n116749, n116750, n116751, n116752, 
      n116753, n116755, n116756, n116757, n116758, n116759, n116760, n116761, 
      n116762, n116763, n116764, n116765, n116767, n116770, n116772, n116773, 
      n116774, n116775, n116776, n116778, n116779, n116780, n116781, n116782, 
      n116783, n116784, n116785, n116786, n116787, n116788, n116790, n116793, 
      n116795, n116796, n116797, n116798, n116799, n116801, n116802, n116803, 
      n116804, n116805, n116806, n116807, n116808, n116809, n116810, n116811, 
      n116813, n116816, n116818, n116819, n116820, n116821, n116822, n116824, 
      n116825, n116826, n116827, n116828, n116829, n116830, n116831, n116832, 
      n116833, n116834, n116836, n116839, n116841, n116842, n116843, n116844, 
      n116845, n116847, n116848, n116849, n116850, n116851, n116852, n116853, 
      n116854, n116855, n116856, n116857, n116859, n116862, n116864, n116865, 
      n116866, n116867, n116868, n116870, n116871, n116872, n116873, n116874, 
      n116875, n116876, n116877, n116878, n116879, n116880, n116882, n116885, 
      n116887, n116888, n116889, n116890, n116891, n116893, n116894, n116895, 
      n116896, n116897, n116898, n116899, n116900, n116901, n116902, n116903, 
      n116905, n116908, n116910, n116911, n116912, n116913, n116914, n116916, 
      n116917, n116918, n116919, n116920, n116921, n116922, n116923, n116924, 
      n116925, n116926, n116928, n116931, n116933, n116934, n116935, n116936, 
      n116937, n116939, n116940, n116941, n116942, n116943, n116944, n116945, 
      n116946, n116947, n116948, n116949, n116951, n116954, n116956, n116957, 
      n116958, n116959, n116960, n116962, n116963, n116964, n116965, n116966, 
      n116967, n116968, n116969, n116970, n116971, n116972, n116974, n116977, 
      n116979, n116980, n116981, n116982, n116983, n116985, n116986, n116987, 
      n116988, n116989, n116990, n116991, n116992, n116993, n116994, n116995, 
      n116997, n117000, n117002, n117003, n117004, n117005, n117006, n117008, 
      n117009, n117010, n117011, n117012, n117013, n117014, n117015, n117016, 
      n117017, n117018, n117020, n117023, n117025, n117026, n117027, n117028, 
      n117029, n117031, n117032, n117033, n117034, n117035, n117036, n117037, 
      n117038, n117039, n117040, n117041, n117043, n117046, n117048, n117049, 
      n117050, n117051, n117052, n117054, n117055, n117056, n117057, n117058, 
      n117059, n117060, n117061, n117062, n117063, n117064, n117066, n117069, 
      n117071, n117072, n117073, n117074, n117075, n117077, n117078, n117079, 
      n117080, n117081, n117082, n117083, n117084, n117085, n117086, n117087, 
      n117089, n117092, n117094, n117095, n117096, n117097, n117098, n117100, 
      n117101, n117102, n117103, n117104, n117105, n117106, n117107, n117108, 
      n117109, n117110, n117112, n117115, n117117, n117118, n117119, n117120, 
      n117121, n117123, n117124, n117125, n117126, n117127, n117128, n117129, 
      n117130, n117131, n117132, n117133, n117135, n117138, n117140, n117141, 
      n117142, n117143, n117144, n117146, n117147, n117148, n117149, n117150, 
      n117151, n117152, n117153, n117154, n117155, n117156, n117158, n117161, 
      n117163, n117164, n117165, n117166, n117167, n117169, n117170, n117171, 
      n117172, n117173, n117174, n117175, n117176, n117177, n117178, n117179, 
      n117181, n117184, n117186, n117187, n117188, n117189, n117190, n117192, 
      n117193, n117194, n117195, n117196, n117197, n117198, n117199, n117200, 
      n117201, n117202, n117204, n117207, n117209, n117210, n117211, n117212, 
      n117213, n117215, n117216, n117217, n117218, n117219, n117220, n117221, 
      n117222, n117223, n117224, n117225, n117227, n117230, n117232, n117233, 
      n117234, n117235, n117236, n117238, n117239, n117240, n117241, n117242, 
      n117243, n117244, n117245, n117246, n117247, n117248, n117250, n117253, 
      n117255, n117256, n117257, n117258, n117259, n117261, n117262, n117263, 
      n117264, n117265, n117266, n117267, n117268, n117269, n117270, n117271, 
      n117273, n117276, n117278, n117279, n117280, n117281, n117282, n117284, 
      n117285, n117286, n117287, n117288, n117289, n117290, n117291, n117292, 
      n117293, n117294, n117296, n117299, n117301, n117302, n117303, n117304, 
      n117305, n117307, n117308, n117309, n117310, n117311, n117312, n117313, 
      n117314, n117315, n117316, n117317, n117319, n117322, n117324, n117325, 
      n117326, n117327, n117328, n117330, n117331, n117332, n117333, n117334, 
      n117335, n117336, n117337, n117338, n117339, n117340, n117342, n117345, 
      n117347, n117348, n117349, n117350, n117351, n117353, n117354, n117355, 
      n117356, n117357, n117358, n117359, n117360, n117361, n117362, n117363, 
      n117365, n117368, n117370, n117371, n117372, n117373, n117374, n117376, 
      n117377, n117378, n117379, n117380, n117381, n117382, n117383, n117384, 
      n117385, n117386, n117388, n117391, n117393, n117394, n117395, n117396, 
      n117397, n117399, n117400, n117401, n117402, n117403, n117404, n117405, 
      n117406, n117407, n117408, n117409, n117411, n117414, n117416, n117417, 
      n117418, n117419, n117420, n117422, n117423, n117424, n117425, n117426, 
      n117427, n117428, n117429, n117430, n117431, n117432, n117434, n117437, 
      n117439, n117440, n117441, n117442, n117443, n117445, n117446, n117447, 
      n117448, n117449, n117450, n117451, n117452, n117453, n117454, n117455, 
      n117457, n117460, n117462, n117463, n117464, n117465, n117466, n117468, 
      n117469, n117470, n117471, n117472, n117473, n117474, n117475, n117476, 
      n117477, n117478, n117480, n117483, n117485, n117486, n117487, n117488, 
      n117489, n117491, n117492, n117493, n117494, n117495, n117496, n117497, 
      n117498, n117499, n117500, n117501, n117503, n117506, n117508, n117509, 
      n117510, n117511, n117512, n117514, n117515, n117516, n117517, n117518, 
      n117519, n117520, n117521, n117522, n117523, n117524, n117526, n117529, 
      n117531, n117532, n117533, n117534, n117535, n117537, n117538, n117539, 
      n117540, n117541, n117542, n117543, n117544, n117545, n117546, n117547, 
      n117549, n117552, n117554, n117555, n117556, n117557, n117558, n117559, 
      n117560, n117561, n117562, n117563, n117564, n117565, n117566, n117567, 
      n117568, n117569, n117571, n117574, n117576, n117577, n117578, n117579, 
      n117580, n117581, n117582, n117583, n117584, n117585, n117586, n117587, 
      n117588, n117589, n117590, n117591, n117593, n117596, n117598, n117599, 
      n117600, n117601, n117602, n117603, n117604, n117605, n117606, n117607, 
      n117608, n117609, n117610, n117611, n117612, n117613, n117615, n117618, 
      n117620, n117621, n117622, n117623, n117624, n117625, n117626, n117627, 
      n117628, n117629, n117630, n117631, n117632, n117633, n117634, n117635, 
      n117637, n117640, n117642, n117643, n117644, n117645, n117646, n117647, 
      n117648, n117649, n117650, n117651, n117652, n117653, n117654, n117655, 
      n117656, n117657, n117659, n117662, n117664, n117665, n117666, n117667, 
      n117668, n117669, n117670, n117671, n117672, n117673, n117674, n117675, 
      n117676, n117677, n117678, n117679, n117681, n117684, n117686, n117687, 
      n117688, n117689, n117690, n117691, n117692, n117693, n117694, n117695, 
      n117696, n117697, n117698, n117699, n117700, n117701, n117703, n117706, 
      n117708, n117709, n117710, n117711, n117712, n117713, n117714, n117715, 
      n117716, n117717, n117718, n117719, n117720, n117721, n117722, n117723, 
      n117725, n117728, n117730, n117731, n117732, n117733, n117734, n117735, 
      n117736, n117737, n117738, n117739, n117740, n117741, n117742, n117743, 
      n117744, n117745, n117747, n117750, n117752, n117753, n117754, n117755, 
      n117756, n117757, n117758, n117759, n117760, n117761, n117762, n117763, 
      n117764, n117765, n117766, n117767, n117769, n117772, n117774, n117775, 
      n117776, n117777, n117778, n117779, n117780, n117781, n117782, n117783, 
      n117784, n117785, n117786, n117787, n117788, n117789, n117791, n117794, 
      n117796, n117797, n117798, n117799, n117800, n117801, n117802, n117803, 
      n117804, n117805, n117806, n117807, n117808, n117809, n117810, n117811, 
      n117813, n117816, n117818, n117819, n117820, n117821, n117822, n117823, 
      n117824, n117825, n117826, n117827, n117828, n117829, n117830, n117831, 
      n117832, n117833, n117835, n117838, n117840, n117841, n117842, n117843, 
      n117844, n117845, n117846, n117847, n117848, n117849, n117850, n117851, 
      n117852, n117853, n117854, n117855, n117857, n117860, n117862, n117863, 
      n117864, n117865, n117866, n117867, n117868, n117869, n117870, n117871, 
      n117872, n117873, n117874, n117875, n117876, n117877, n117879, n117882, 
      n117884, n117885, n117886, n117887, n117888, n117889, n117890, n117891, 
      n117892, n117893, n117894, n117895, n117896, n117897, n117898, n117899, 
      n117901, n117904, n117906, n117907, n117908, n117909, n117910, n117911, 
      n117912, n117913, n117914, n117915, n117916, n117917, n117918, n117919, 
      n117920, n117921, n117923, n117926, n117928, n117929, n117930, n117931, 
      n117932, n117933, n117934, n117935, n117936, n117937, n117938, n117939, 
      n117940, n117941, n117942, n117943, n117945, n117946, n117947, n117948, 
      n117949, n117950, n117953, n117954, n117955, n117956, n117958, n117959, 
      n117960, n117961, n117962, n117963, n117964, n117965, n117966, n117967, 
      n117968, n117969, n117970, n117971, n117972, n117973, n117974, n117975, 
      n117976, n117977, n117981, n117982, n117983, n117984, n117985, n117986, 
      n117987, n117988, n117993, n117994, n117995, n117996, n118070, n118071, 
      n118072, n118073, n118074, n118075, n118076, n118077, n118078, n118079, 
      n118080, n118081, n118082, n118083, n118084, n118205, n118206, n118207, 
      n118208, n118209, n118210, n118211, n118212, n118213, n118214, n118215, 
      n118216, n118217, n118218, n118219, n118220, n118221, n118222, n118223, 
      n118224, n118225, n118226, n118227, n118228, n118229, n118230, n118231, 
      n118232, n118233, n118234, n118235, n118236, n118237, n118238, n118239, 
      n118240, n118241, n118242, n118243, n118244, n118245, n118246, n118247, 
      n118248, n118249, n118250, n118251, n118252, n118253, n118254, n118255, 
      n118256, n118257, n118258, n118259, n118260, n118261, n118262, n118263, 
      n118264, n118325, n118326, n118327, n118328, n118329, n118330, n118331, 
      n118332, n118333, n118334, n118335, n118336, n118337, n118338, n118339, 
      n118340, n118341, n118342, n118343, n118344, n118345, n118346, n118347, 
      n118348, n118349, n118350, n118351, n118352, n118353, n118354, n118355, 
      n118356, n118357, n118358, n118359, n118360, n118361, n118362, n118363, 
      n118364, n118365, n118366, n118367, n118368, n118369, n118370, n118371, 
      n118372, n118373, n118374, n118375, n118376, n118377, n118378, n118379, 
      n118380, n118381, n118382, n118383, n118384, n118385, n118386, n118387, 
      n118388, n118389, n118390, n118391, n118392, n118393, n118394, n118395, 
      n118396, n118397, n118398, n118399, n118400, n118401, n118402, n118403, 
      n118404, n118405, n118406, n118407, n118408, n118409, n118410, n118411, 
      n118412, n118413, n118414, n118415, n118416, n118417, n118418, n118419, 
      n118420, n118421, n118422, n118423, n118424, n118425, n118426, n118427, 
      n118428, n118429, n118430, n118431, n118432, n118433, n118434, n118435, 
      n118436, n118437, n118438, n118439, n118440, n118441, n118442, n118443, 
      n118444, n118505, n118506, n118507, n118508, n118509, n118510, n118511, 
      n118512, n118513, n118514, n118515, n118516, n118517, n118518, n118519, 
      n118520, n118521, n118522, n118523, n118524, n118525, n118526, n118527, 
      n118528, n118529, n118530, n118531, n118532, n118533, n118534, n118535, 
      n118536, n118537, n118538, n118539, n118540, n118541, n118542, n118543, 
      n118544, n118545, n118546, n118547, n118548, n118549, n118550, n118551, 
      n118552, n118553, n118554, n118555, n118556, n118557, n118558, n118559, 
      n118560, n118561, n118562, n118563, n118564, n118565, n118566, n118567, 
      n118568, n118569, n118570, n118571, n118572, n118573, n118574, n118575, 
      n118576, n118577, n118578, n118579, n118580, n118581, n118582, n118583, 
      n118584, n118585, n118586, n118587, n118588, n118589, n118590, n118591, 
      n118592, n118593, n118594, n118595, n118596, n118597, n118598, n118599, 
      n118600, n118601, n118602, n118603, n118604, n118605, n118606, n118607, 
      n118608, n118609, n118610, n118611, n118612, n118613, n118614, n118615, 
      n118616, n118617, n118618, n118619, n118620, n118621, n118622, n118623, 
      n118624, n118625, n118626, n118627, n118628, n118629, n118630, n118631, 
      n118632, n118633, n118634, n118635, n118636, n118637, n118638, n118639, 
      n118640, n118641, n118642, n118643, n118644, n118645, n118646, n118647, 
      n118648, n118649, n118650, n118651, n118652, n118653, n118654, n118655, 
      n118656, n118657, n118658, n118659, n118660, n118661, n118662, n118663, 
      n118664, n118665, n118666, n118667, n118668, n118669, n118670, n118671, 
      n118672, n118673, n118674, n118675, n118676, n118677, n118678, n118679, 
      n118680, n118681, n118682, n118683, n118684, n118685, n118686, n118687, 
      n118688, n118689, n118690, n118691, n118692, n118693, n118694, n118695, 
      n118696, n118697, n118698, n118699, n118700, n118701, n118702, n118703, 
      n118704, n118705, n118706, n118707, n118708, n118709, n118710, n118711, 
      n118712, n118713, n118714, n118715, n118716, n118717, n118718, n118719, 
      n118720, n118721, n118722, n118723, n118724, n118725, n118726, n118727, 
      n118728, n118729, n118730, n118731, n118732, n118733, n118734, n118735, 
      n118736, n118737, n118738, n118739, n118740, n118741, n118742, n118743, 
      n118744, n118745, n118746, n118747, n118748, n118749, n118750, n118751, 
      n118752, n118753, n118754, n118755, n118756, n118757, n118758, n118759, 
      n118760, n118761, n118762, n118763, n118764, n118765, n118766, n118767, 
      n118768, n118769, n118770, n118771, n118772, n118773, n118774, n118775, 
      n118776, n118777, n118778, n118779, n118780, n118781, n118782, n118783, 
      n118784, n118785, n118786, n118787, n118788, n118789, n118790, n118791, 
      n118792, n118793, n118794, n118795, n118796, n118797, n118798, n118799, 
      n118800, n118801, n118802, n118803, n118804, n118805, n118806, n118807, 
      n118808, n118809, n118810, n118811, n118812, n118813, n118814, n118815, 
      n118816, n118817, n118818, n118819, n118820, n118821, n118822, n118823, 
      n118824, n118825, n118826, n118827, n118828, n118829, n118830, n118831, 
      n118832, n118833, n118834, n118835, n118836, n118837, n118838, n118839, 
      n118840, n118841, n118842, n118843, n118844, n118845, n118846, n118847, 
      n118848, n118849, n118850, n118851, n118852, n118853, n118854, n118855, 
      n118856, n118857, n118858, n118859, n118860, n118861, n118862, n118863, 
      n118864, n118865, n118866, n118867, n118868, n118869, n118870, n118871, 
      n118872, n118873, n118874, n118875, n118876, n118877, n118878, n118879, 
      n118880, n118881, n118882, n118883, n118884, n118885, n118886, n118887, 
      n118888, n118889, n118890, n118891, n118892, n118893, n118894, n118895, 
      n118896, n118897, n118898, n118899, n118900, n118901, n118902, n118903, 
      n118904, n118905, n118906, n118907, n118908, n118909, n118910, n118911, 
      n118912, n118913, n118914, n118915, n118916, n118917, n118918, n118919, 
      n118920, n118921, n118922, n118923, n118924, n118925, n118926, n118927, 
      n118928, n118929, n118930, n118931, n118932, n118933, n118934, n118935, 
      n118936, n118937, n118938, n118939, n118940, n118941, n118942, n118943, 
      n118944, n118945, n118946, n118947, n118948, n118949, n118950, n118951, 
      n118952, n118953, n118954, n118955, n118956, n118957, n118958, n118959, 
      n118960, n118961, n118962, n118963, n118964, n118965, n118966, n118967, 
      n118968, n118969, n118970, n118971, n118972, n118973, n118974, n118975, 
      n118976, n118977, n118978, n118979, n118980, n118981, n118982, n118983, 
      n118984, n118985, n118986, n118987, n118988, n118989, n118990, n118991, 
      n118992, n118993, n118994, n118995, n118996, n118997, n118998, n118999, 
      n119000, n119001, n119002, n119003, n119004, n119005, n119006, n119007, 
      n119008, n119009, n119010, n119011, n119012, n119013, n119014, n119015, 
      n119016, n119017, n119018, n119019, n119020, n119021, n119022, n119023, 
      n119024, n119025, n119026, n119027, n119028, n119029, n119030, n119031, 
      n119032, n119033, n119034, n119035, n119036, n119037, n119038, n119039, 
      n119040, n119041, n119042, n119043, n119044, n119045, n119046, n119047, 
      n119048, n119049, n119050, n119051, n119052, n119053, n119054, n119055, 
      n119056, n119057, n119058, n119059, n119060, n119061, n119062, n119063, 
      n119064, n119065, n119066, n119067, n119068, n119069, n119070, n119071, 
      n119072, n119073, n119074, n119075, n119076, n119077, n119078, n119079, 
      n119080, n119081, n119082, n119083, n119084, n119085, n119086, n119087, 
      n119088, n119089, n119090, n119091, n119092, n119093, n119094, n119095, 
      n119096, n119097, n119098, n119099, n119100, n119101, n119102, n119103, 
      n119104, n119105, n119106, n119107, n119108, n119109, n119110, n119111, 
      n119112, n119113, n119114, n119115, n119116, n119117, n119118, n119119, 
      n119120, n119121, n119122, n119123, n119124, n119125, n119126, n119127, 
      n119128, n119129, n119130, n119131, n119132, n119133, n119134, n119135, 
      n119136, n119137, n119138, n119139, n119140, n119141, n119142, n119143, 
      n119144, n119145, n119146, n119147, n119148, n119149, n119150, n119151, 
      n119152, n119153, n119154, n119155, n119156, n119157, n119158, n119159, 
      n119160, n119161, n119162, n119163, n119164, n119165, n119166, n119167, 
      n119168, n119169, n119170, n119171, n119172, n119173, n119174, n119175, 
      n119176, n119177, n119178, n119179, n119180, n119181, n119182, n119183, 
      n119184, n119185, n119186, n119187, n119188, n119189, n119190, n119191, 
      n119192, n119193, n119194, n119195, n119196, n119197, n119198, n119199, 
      n119200, n119201, n119202, n119203, n119204, n119205, n119206, n119207, 
      n119208, n119209, n119210, n119211, n119212, n119213, n119214, n119215, 
      n119216, n119217, n119218, n119219, n119220, n119221, n119222, n119223, 
      n119224, n119225, n119226, n119227, n119228, n119229, n119230, n119231, 
      n119232, n119233, n119234, n119235, n119236, n119237, n119238, n119239, 
      n119240, n119241, n119242, n119243, n119244, n119245, n119246, n119247, 
      n119248, n119249, n119250, n119251, n119252, n119253, n119254, n119255, 
      n119256, n119257, n119258, n119259, n119260, n119261, n119262, n119263, 
      n119264, n119265, n119266, n119267, n119268, n119269, n119270, n119271, 
      n119272, n119273, n119274, n119275, n119276, n119277, n119278, n119279, 
      n119280, n119281, n119282, n119283, n119284, n119285, n119286, n119287, 
      n119288, n119289, n119290, n119291, n119292, n119293, n119294, n119295, 
      n119296, n119297, n119298, n119299, n119300, n119301, n119302, n119303, 
      n119304, n119305, n119306, n119307, n119308, n119309, n119310, n119311, 
      n119312, n119313, n119314, n119315, n119316, n119317, n119318, n119319, 
      n119320, n119321, n119322, n119323, n119324, n119325, n119326, n119327, 
      n119328, n119329, n119330, n119331, n119332, n119333, n119334, n119335, 
      n119336, n119337, n119338, n119339, n119340, n119341, n119342, n119343, 
      n119344, n119345, n119346, n119347, n119348, n119349, n119350, n119351, 
      n119352, n119353, n119354, n119355, n119356, n119357, n119358, n119359, 
      n119360, n119361, n119362, n119363, n119364, n119365, n119366, n119367, 
      n119368, n119369, n119370, n119371, n119372, n119373, n119374, n119375, 
      n119376, n119377, n119378, n119379, n119380, n119381, n119382, n119383, 
      n119384, n119385, n119386, n119387, n119388, n119389, n119390, n119391, 
      n119392, n119393, n119394, n119395, n119396, n119397, n119398, n119399, 
      n119400, n119401, n119402, n119403, n119404, n119405, n119406, n119407, 
      n119408, n119409, n119410, n119411, n119412, n119413, n119414, n119415, 
      n119416, n119417, n119418, n119419, n119420, n119421, n119422, n119423, 
      n119424, n119425, n119426, n119427, n119428, n119429, n119430, n119431, 
      n119432, n119433, n119434, n119435, n119436, n119437, n119438, n119439, 
      n119440, n119441, n119442, n119443, n119444, n119445, n119446, n119447, 
      n119448, n119449, n119450, n119451, n119452, n119453, n119454, n119455, 
      n119456, n119457, n119458, n119459, n119460, n119461, n119462, n119463, 
      n119464, n119465, n119466, n119467, n119468, n119469, n119470, n119471, 
      n119472, n119473, n119474, n119475, n119476, n119477, n119478, n119479, 
      n119480, n119481, n119482, n119483, n119484, n119485, n119486, n119487, 
      n119488, n119489, n119490, n119491, n119492, n119493, n119494, n119495, 
      n119496, n119497, n119498, n119499, n119500, n119501, n119502, n119503, 
      n119504, n119505, n119506, n119507, n119508, n119509, n119510, n119511, 
      n119512, n119513, n119514, n119515, n119516, n119517, n119518, n119519, 
      n119520, n119521, n119522, n119523, n119524, n119525, n119526, n119527, 
      n119528, n119529, n119530, n119531, n119532, n119533, n119534, n119535, 
      n119536, n119537, n119538, n119539, n119540, n119541, n119542, n119543, 
      n119544, n119545, n119546, n119547, n119548, n119549, n119550, n119551, 
      n119552, n119553, n119554, n119555, n119556, n119557, n119558, n119559, 
      n119560, n119561, n119562, n119563, n119564, n119565, n119566, n119567, 
      n119568, n119569, n119570, n119571, n119572, n119573, n119574, n119575, 
      n119576, n119577, n119578, n119579, n119580, n119581, n119582, n119583, 
      n119584, n119585, n119586, n119587, n119588, n119589, n119590, n119591, 
      n119592, n119593, n119594, n119595, n119596, n119597, n119598, n119599, 
      n119600, n119601, n119602, n119603, n119604, n119605, n119606, n119607, 
      n119608, n119609, n119610, n119611, n119612, n119613, n119614, n119615, 
      n119616, n119617, n119618, n119619, n119620, n119621, n119622, n119623, 
      n119624, n119625, n119626, n119627, n119628, n119629, n119630, n119631, 
      n119632, n119633, n119634, n119635, n119636, n119637, n119638, n119639, 
      n119640, n119641, n119642, n119643, n119644, n119645, n119646, n119647, 
      n119648, n119649, n119650, n119651, n119652, n119653, n119654, n119655, 
      n119656, n119657, n119658, n119659, n119660, n119661, n119662, n119663, 
      n119664, n119665, n119666, n119667, n119668, n119669, n119670, n119671, 
      n119672, n119673, n119674, n119675, n119676, n119677, n119678, n119679, 
      n119680, n119681, n119682, n119683, n119684, n119685, n119686, n119687, 
      n119688, n119689, n119690, n119691, n119692, n119693, n119694, n119695, 
      n119696, n119697, n119698, n119699, n119700, n119701, n119702, n119703, 
      n119704, n119705, n119706, n119707, n119708, n119709, n119710, n119711, 
      n119712, n119713, n119714, n119715, n119716, n119717, n119718, n119719, 
      n119720, n119721, n119722, n119723, n119724, n119725, n119726, n119727, 
      n119728, n119729, n119730, n119731, n119732, n119733, n119734, n119735, 
      n119736, n119737, n119738, n119739, n119740, n119741, n119742, n119743, 
      n119744, n119745, n119746, n119747, n119748, n119749, n119750, n119751, 
      n119752, n119753, n119754, n119755, n119756, n119757, n119758, n119759, 
      n119760, n119761, n119762, n119763, n119764, n119765, n119766, n119767, 
      n119768, n119769, n119770, n119771, n119772, n119773, n119774, n119775, 
      n119776, n119777, n119778, n119779, n119780, n119781, n119782, n119783, 
      n119784, n119785, n119786, n119787, n119788, n119789, n119790, n119791, 
      n119792, n119793, n119794, n119795, n119796, n119797, n119798, n119799, 
      n119800, n119801, n119802, n119803, n119804, n119805, n119806, n119807, 
      n119808, n119809, n119810, n119811, n119812, n119813, n119814, n119815, 
      n119816, n119817, n119818, n119819, n119820, n119821, n119822, n119823, 
      n119824, n119825, n119826, n119827, n119828, n119829, n119830, n119831, 
      n119832, n119833, n119834, n119835, n119836, n119837, n119838, n119839, 
      n119840, n119841, n119842, n119843, n119844, n119845, n119846, n119847, 
      n119848, n119849, n119850, n119851, n119852, n119853, n119854, n119855, 
      n119856, n119857, n119858, n119859, n119860, n119861, n119862, n119863, 
      n119864, n119865, n119866, n119867, n119868, n119869, n119870, n119871, 
      n119872, n119873, n119874, n119875, n119876, n119877, n119878, n119879, 
      n119880, n119881, n119882, n119883, n119884, n119885, n119886, n119887, 
      n119888, n119889, n119890, n119891, n119892, n119893, n119894, n119895, 
      n119896, n119897, n119898, n119899, n119900, n119901, n119902, n119903, 
      n119904, n119905, n119906, n119907, n119908, n119909, n119910, n119911, 
      n119912, n119913, n119914, n119915, n119916, n119917, n119918, n119919, 
      n119920, n119921, n119922, n119923, n119924, n119925, n119926, n119927, 
      n119928, n119929, n119930, n119931, n119932, n119933, n119934, n119935, 
      n119936, n119937, n119938, n119939, n119940, n119941, n119942, n119943, 
      n119944, n119945, n119946, n119947, n119948, n119949, n119950, n119951, 
      n119952, n119953, n119954, n119955, n119956, n119957, n119958, n119959, 
      n119960, n119961, n119962, n119963, n119964, n119965, n119966, n119967, 
      n119968, n119969, n119970, n119971, n119972, n119973, n119974, n119975, 
      n119976, n119977, n119978, n119979, n119980, n119981, n119982, n119983, 
      n119984, n119985, n119986, n119987, n119988, n119989, n119990, n119991, 
      n119992, n119993, n119994, n119995, n119996, n119997, n119998, n119999, 
      n120000, n120001, n120002, n120003, n120004, n120005, n120006, n120007, 
      n120008, n120009, n120010, n120011, n120012, n120013, n120014, n120015, 
      n120016, n120017, n120018, n120019, n120020, n120021, n120022, n120023, 
      n120024, n120025, n120026, n120027, n120028, n120029, n120030, n120031, 
      n120032, n120033, n120034, n120035, n120036, n120037, n120038, n120039, 
      n120040, n120041, n120042, n120043, n120044, n120045, n120046, n120047, 
      n120048, n120049, n120050, n120051, n120052, n120053, n120054, n120055, 
      n120056, n120057, n120058, n120059, n120060, n120061, n120062, n120063, 
      n120064, n120065, n120066, n120067, n120068, n120069, n120070, n120071, 
      n120072, n120073, n120074, n120075, n120076, n120077, n120078, n120079, 
      n120080, n120081, n120082, n120083, n120084, n120085, n120086, n120087, 
      n120088, n120089, n120090, n120091, n120092, n120093, n120094, n120095, 
      n120096, n120097, n120098, n120099, n120100, n120101, n120102, n120103, 
      n120104, n120105, n120106, n120107, n120108, n120109, n120110, n120111, 
      n120112, n120113, n120114, n120115, n120116, n120117, n120118, n120119, 
      n120120, n120121, n120122, n120123, n120124, n120125, n120126, n120127, 
      n120128, n120129, n120130, n120131, n120132, n120133, n120134, n120135, 
      n120136, n120137, n120138, n120139, n120140, n120141, n120142, n120143, 
      n120144, n120145, n120146, n120147, n120148, n120149, n120150, n120151, 
      n120152, n120153, n120154, n120155, n120156, n120157, n120158, n120159, 
      n120160, n120161, n120162, n120163, n120164, n120165, n120166, n120167, 
      n120168, n120169, n120170, n120171, n120172, n120173, n120174, n120175, 
      n120176, n120177, n120178, n120179, n120180, n120181, n120182, n120183, 
      n120184, n120185, n120186, n120187, n120188, n120189, n120190, n120191, 
      n120192, n120193, n120194, n120195, n120196, n120197, n120198, n120199, 
      n120200, n120201, n120202, n120203, n120204, n120205, n120206, n120207, 
      n120208, n120209, n120210, n120211, n120212, n120213, n120214, n120215, 
      n120216, n120217, n120218, n120219, n120220, n120221, n120222, n120223, 
      n120224, n120225, n120226, n120227, n120228, n120229, n120230, n120231, 
      n120232, n120233, n120234, n120235, n120236, n120237, n120238, n120239, 
      n120240, n120241, n120242, n120243, n120244, n120245, n120246, n120247, 
      n120248, n120249, n120250, n120251, n120252, n120253, n120254, n120255, 
      n120256, n120257, n120258, n120259, n120260, n120261, n120262, n120263, 
      n120264, n120265, n120266, n120267, n120268, n120269, n120270, n120271, 
      n120272, n120273, n120274, n120275, n120276, n120277, n120278, n120279, 
      n120280, n120281, n120282, n120283, n120284, n120285, n120286, n120287, 
      n120288, n120289, n120290, n120291, n120292, n120293, n120294, n120295, 
      n120296, n120297, n120298, n120299, n120300, n120301, n120302, n120303, 
      n120304, n120305, n120306, n120307, n120308, n120309, n120310, n120311, 
      n120312, n120313, n120314, n120315, n120316, n120317, n120318, n120319, 
      n120320, n120321, n120322, n120323, n120324, n120325, n120326, n120327, 
      n120328, n120329, n120330, n120331, n120332, n120333, n120334, n120335, 
      n120336, n120337, n120338, n120339, n120340, n120341, n120342, n120343, 
      n120344, n120345, n120346, n120347, n120348, n120349, n120350, n120351, 
      n120352, n120353, n120354, n120355, n120356, n120357, n120358, n120359, 
      n120360, n120361, n120362, n120363, n120364, n120365, n120366, n120367, 
      n120368, n120369, n120370, n120371, n120372, n120373, n120374, n120375, 
      n120376, n120377, n120378, n120379, n120380, n120381, n120382, n120383, 
      n120384, n120385, n120386, n120387, n120388, n120389, n120390, n120391, 
      n120392, n120393, n120394, n120395, n120396, n120397, n120398, n120399, 
      n120400, n120401, n120402, n120403, n120404, n120405, n120406, n120407, 
      n120408, n120409, n120410, n120411, n120412, n120413, n120414, n120415, 
      n120416, n120417, n120418, n120419, n120420, n120421, n120422, n120423, 
      n120424, n120425, n120426, n120427, n120428, n120429, n120430, n120431, 
      n120432, n120433, n120434, n120435, n120436, n120437, n120438, n120439, 
      n120440, n120441, n120442, n120443, n120444, n120445, n120446, n120447, 
      n120448, n120449, n120450, n120451, n120452, n120453, n120454, n120455, 
      n120456, n120457, n120458, n120459, n120460, n120461, n120462, n120463, 
      n120464, n120465, n120466, n120467, n120468, n120469, n120470, n120471, 
      n120472, n120473, n120474, n120475, n120476, n120477, n120478, n120479, 
      n120480, n120481, n120482, n120483, n120484, n120485, n120486, n120487, 
      n120488, n120489, n120490, n120491, n120492, n120493, n120494, n120495, 
      n120496, n120497, n120498, n120499, n120500, n120501, n120502, n120503, 
      n120504, n120505, n120506, n120507, n120508, n120509, n120510, n120511, 
      n120512, n120513, n120514, n120515, n120516, n120517, n120518, n120519, 
      n120520, n120521, n120522, n120523, n120524, n120525, n120526, n120527, 
      n120528, n120529, n120530, n120531, n120532, n120533, n120534, n120535, 
      n120536, n120537, n120538, n120539, n120540, n120541, n120542, n120543, 
      n120544, n120545, n120546, n120547, n120548, n120549, n120550, n120551, 
      n120552, n120553, n120554, n120555, n120556, n120557, n120558, n120559, 
      n120560, n120561, n120562, n120563, n120564, n120565, n120566, n120567, 
      n120568, n120569, n120570, n120571, n120572, n120573, n120574, n120575, 
      n120576, n120577, n120578, n120579, n120580, n120581, n120582, n120583, 
      n120584, n120585, n120586, n120587, n120588, n120589, n120590, n120591, 
      n120592, n120593, n120594, n120595, n120596, n120597, n120598, n120599, 
      n120600, n120601, n120602, n120603, n120604, n120605, n120606, n120607, 
      n120608, n120609, n120610, n120611, n120612, n120613, n120614, n120615, 
      n120616, n120617, n120618, n120619, n120620, n120621, n120622, n120623, 
      n120624, n120625, n120626, n120627, n120628, n120629, n120630, n120631, 
      n120632, n120633, n120634, n120635, n120636, n120637, n120638, n120639, 
      n120640, n120641, n120642, n120643, n120644, n120645, n120646, n120647, 
      n120648, n120649, n120650, n120651, n120652, n120653, n120654, n120655, 
      n120656, n120657, n120658, n120659, n120660, n120661, n120662, n120663, 
      n120664, n120665, n120666, n120667, n120668, n120669, n120670, n120671, 
      n120672, n120673, n120674, n120675, n120676, n120677, n120678, n120679, 
      n120680, n120681, n120682, n120683, n120684, n120685, n120686, n120687, 
      n120688, n120689, n120690, n120691, n120692, n120693, n120694, n120695, 
      n120696, n120697, n120698, n120699, n120700, n120701, n120702, n120703, 
      n120704, n120705, n120706, n120707, n120708, n120709, n120710, n120711, 
      n120712, n120713, n120714, n120715, n120716, n120717, n120718, n120719, 
      n120720, n120721, n120722, n120723, n120724, n120725, n120726, n120727, 
      n120728, n120729, n120730, n120731, n120732, n120733, n120734, n120735, 
      n120736, n120737, n120738, n120739, n120740, n120741, n120742, n120743, 
      n120744, n120745, n120746, n120747, n120748, n120749, n120750, n120751, 
      n120752, n120753, n120754, n120755, n120756, n120757, n120758, n120759, 
      n120760, n120761, n120762, n120763, n120764, n120765, n120766, n120767, 
      n120768, n120769, n120770, n120771, n120772, n120773, n120774, n120775, 
      n120776, n120777, n120778, n120779, n120780, n120781, n120782, n120783, 
      n120784, n120785, n120786, n120787, n120788, n120789, n120790, n120791, 
      n120792, n120793, n120794, n120795, n120796, n120797, n120798, n120799, 
      n120800, n120801, n120802, n120803, n120804, n120805, n120806, n120807, 
      n120808, n120809, n120810, n120811, n120812, n120813, n120814, n120815, 
      n120816, n120817, n120818, n120819, n120820, n120821, n120822, n120823, 
      n120824, n120825, n120826, n120827, n120828, n120829, n120830, n120831, 
      n120832, n120833 : std_logic;

begin
   OUT1 <= ( OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, 
      OUT1_59_port, OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, 
      OUT1_54_port, OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, 
      OUT1_49_port, OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, 
      OUT1_44_port, OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, 
      OUT1_39_port, OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, 
      OUT1_34_port, OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, 
      OUT1_29_port, OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, 
      OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, 
      OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, 
      OUT1_14_port, OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, 
      OUT1_9_port, OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, 
      OUT1_4_port, OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_63_port, OUT2_62_port, OUT2_61_port, OUT2_60_port, 
      OUT2_59_port, OUT2_58_port, OUT2_57_port, OUT2_56_port, OUT2_55_port, 
      OUT2_54_port, OUT2_53_port, OUT2_52_port, OUT2_51_port, OUT2_50_port, 
      OUT2_49_port, OUT2_48_port, OUT2_47_port, OUT2_46_port, OUT2_45_port, 
      OUT2_44_port, OUT2_43_port, OUT2_42_port, OUT2_41_port, OUT2_40_port, 
      OUT2_39_port, OUT2_38_port, OUT2_37_port, OUT2_36_port, OUT2_35_port, 
      OUT2_34_port, OUT2_33_port, OUT2_32_port, OUT2_31_port, OUT2_30_port, 
      OUT2_29_port, OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, 
      OUT2_24_port, OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, 
      OUT2_19_port, OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, 
      OUT2_14_port, OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, 
      OUT2_9_port, OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, 
      OUT2_4_port, OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   OUT1_reg_45_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => OUT1_45_port
                           , QN => n4268);
   OUT1_reg_44_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => OUT1_44_port
                           , QN => n4267);
   OUT1_reg_43_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => OUT1_43_port
                           , QN => n4266);
   OUT1_reg_42_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => OUT1_42_port
                           , QN => n4265);
   OUT1_reg_41_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => OUT1_41_port
                           , QN => n4264);
   OUT1_reg_40_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => OUT1_40_port
                           , QN => n4263);
   OUT1_reg_39_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => OUT1_39_port
                           , QN => n4262);
   OUT1_reg_38_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => OUT1_38_port
                           , QN => n4261);
   OUT1_reg_37_inst : DFF_X1 port map( D => n5449, CK => CLK, Q => OUT1_37_port
                           , QN => n4260);
   OUT1_reg_36_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => OUT1_36_port
                           , QN => n4259);
   OUT1_reg_35_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => OUT1_35_port
                           , QN => n4258);
   OUT1_reg_34_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => OUT1_34_port
                           , QN => n4257);
   OUT1_reg_33_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => OUT1_33_port
                           , QN => n4256);
   OUT1_reg_32_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => OUT1_32_port
                           , QN => n4255);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => OUT1_31_port
                           , QN => n4254);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => OUT1_30_port
                           , QN => n4253);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => OUT1_29_port
                           , QN => n4252);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => OUT1_28_port
                           , QN => n4251);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => OUT1_27_port
                           , QN => n4250);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => OUT1_26_port
                           , QN => n4249);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => OUT1_25_port
                           , QN => n4248);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => OUT1_24_port
                           , QN => n4247);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => OUT1_23_port
                           , QN => n4246);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => OUT1_22_port
                           , QN => n4245);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5417, CK => CLK, Q => OUT1_21_port
                           , QN => n4244);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5415, CK => CLK, Q => OUT1_20_port
                           , QN => n4243);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => OUT1_19_port
                           , QN => n4242);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => OUT1_18_port
                           , QN => n4241);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => OUT1_17_port
                           , QN => n4240);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => OUT1_16_port
                           , QN => n4239);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => OUT1_15_port
                           , QN => n4238);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => OUT1_14_port
                           , QN => n4237);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => OUT1_13_port
                           , QN => n4236);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => OUT1_12_port
                           , QN => n4235);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => OUT1_11_port
                           , QN => n4234);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => OUT1_10_port
                           , QN => n4233);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => OUT1_9_port, 
                           QN => n4232);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => OUT1_8_port, 
                           QN => n4231);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => OUT1_7_port, 
                           QN => n4230);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => OUT1_6_port, 
                           QN => n4229);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => OUT1_5_port, 
                           QN => n4228);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => OUT1_4_port, 
                           QN => n4227);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5317, CK => CLK, Q => OUT2_6_port, 
                           QN => n4165);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5316, CK => CLK, Q => OUT2_5_port, 
                           QN => n4164);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5315, CK => CLK, Q => OUT2_4_port, 
                           QN => n4163);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5314, CK => CLK, Q => OUT2_3_port, 
                           QN => n4162);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5313, CK => CLK, Q => OUT2_2_port, 
                           QN => n4161);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5312, CK => CLK, Q => OUT2_1_port, 
                           QN => n4160);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5311, CK => CLK, Q => OUT2_0_port, 
                           QN => n4159);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n118718, QN => n90036);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n118717, QN => n90037);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n118716, QN => n90038);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n118715, QN => n90039);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n118714, QN => n90040);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n118713, QN => n90041);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n118712, QN => n90042);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n118711, QN => n90043);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n118710, QN => n90044);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n118709, QN => n90045);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n118708, QN => n90046);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n118707, QN => n90047);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n118706, QN => n90048);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n118705, QN => n90049);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n118704, QN => n90050);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n118703, QN => n90051);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n118702, QN => n90052);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n118701, QN => n90053);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n118700, QN => n90054);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n118699, QN => n90055);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n118698, QN => n90056);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n118697, QN => n90057);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n118696, QN => n90058);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n118695, QN => n90059);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n118694, QN => n90060);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n118693, QN => n90061);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n118692, QN => n90062);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n118691, QN => n90063);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n118690, QN => n90064);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n118689, QN => n90065);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n118688, QN => n90066);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n118687, QN => n90067);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n118686, QN => n90068);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n118685, QN => n90069);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n118684, QN => n90070);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n118683, QN => n90071);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n118682, QN => n90072);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n118681, QN => n90073);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n118680, QN => n90074);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n118679, QN => n90075);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n118678, QN => n90076);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n118677, QN => n90077);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n118676, QN => n90078);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n118675, QN => n90079);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n118674, QN => n90080);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n118673, QN => n90081);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n118672, QN => n90082);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n118671, QN => n90083);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n118670, QN => n90084);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n118730, QN => n90085);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => 
                           n118729, QN => n90086);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => 
                           n118728, QN => n90087);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => 
                           n118727, QN => n90088);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => 
                           n118737, QN => n90089);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => 
                           n118736, QN => n90090);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => 
                           n118735, QN => n90091);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => 
                           n118734, QN => n90092);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => 
                           n118733, QN => n90093);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => 
                           n118732, QN => n90094);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => 
                           n118731, QN => n90095);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5321, CK => CLK, Q => OUT2_10_port
                           , QN => n94639);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5320, CK => CLK, Q => OUT2_9_port, 
                           QN => n94638);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5319, CK => CLK, Q => OUT2_8_port, 
                           QN => n94637);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5318, CK => CLK, Q => OUT2_7_port, 
                           QN => n94636);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => 
                           n118985, QN => n90711);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n118984, QN => n90713);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n118983, QN => n90714);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n118982, QN => n90715);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => 
                           n118549, QN => n90373);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n118548, QN => n90375);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n118547, QN => n90376);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n118546, QN => n90377);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => 
                           n110482, QN => n90306);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n110481, QN => n90308);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n110480, QN => n90309);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n110479, QN => n90310);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => 
                           n118861, QN => n90512);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n118860, QN => n90514);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n118859, QN => n90515);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n118858, QN => n90516);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7486, CK => CLK, Q => 
                           n110110, QN => n89493);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7485, CK => CLK, Q => 
                           n110109, QN => n89496);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7484, CK => CLK, Q => 
                           n110108, QN => n89498);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7483, CK => CLK, Q => 
                           n110107, QN => n89500);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => 
                           n110366, QN => n89965);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => 
                           n110365, QN => n89967);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n110364, QN => n89968);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n110363, QN => n89969);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => 
                           n118726, QN => n90031);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n118725, QN => n90033);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n118724, QN => n90034);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n118723, QN => n90035);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n118999, QN => n90716);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n118998, QN => n90717);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n118997, QN => n90718);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n118996, QN => n90719);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n118995, QN => n90720);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n118994, QN => n90721);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n118993, QN => n90722);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n118992, QN => n90723);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n118991, QN => n90724);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n118990, QN => n90725);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n118989, QN => n90726);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n118988, QN => n90727);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n118987, QN => n90728);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n118986, QN => n90729);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n119045, QN => n90730);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n119044, QN => n90731);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n119043, QN => n90732);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n119042, QN => n90733);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n119041, QN => n90734);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => 
                           n119040, QN => n90735);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => 
                           n119039, QN => n90736);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => 
                           n119038, QN => n90737);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => 
                           n119037, QN => n90738);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => 
                           n119036, QN => n90739);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => 
                           n119035, QN => n90740);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => 
                           n119034, QN => n90741);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => 
                           n119033, QN => n90742);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => 
                           n119032, QN => n90743);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => 
                           n119031, QN => n90744);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n119030, QN => n90745);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n119029, QN => n90746);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n119028, QN => n90747);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n119027, QN => n90748);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n119026, QN => n90749);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n119025, QN => n90750);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n119024, QN => n90751);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n119023, QN => n90752);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n119022, QN => n90753);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n119021, QN => n90754);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n119020, QN => n90755);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n119019, QN => n90756);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n119018, QN => n90757);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n119017, QN => n90758);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n119016, QN => n90759);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n119015, QN => n90760);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n119014, QN => n90761);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n119013, QN => n90762);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n119012, QN => n90763);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n119011, QN => n90764);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n119010, QN => n90765);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n119009, QN => n90766);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => 
                           n119008, QN => n90767);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => 
                           n119007, QN => n90768);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => 
                           n119006, QN => n90769);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => 
                           n119005, QN => n90770);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => 
                           n119004, QN => n90771);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => 
                           n119003, QN => n90772);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => 
                           n119002, QN => n90773);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => 
                           n119001, QN => n90774);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => 
                           n119000, QN => n90775);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n118563, QN => n90378);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n118562, QN => n90379);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n118561, QN => n90380);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n118560, QN => n90381);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n118559, QN => n90382);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n118558, QN => n90383);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n118557, QN => n90384);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n118556, QN => n90385);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n118555, QN => n90386);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n118554, QN => n90387);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n118553, QN => n90388);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n118552, QN => n90389);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n118551, QN => n90390);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n118550, QN => n90391);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n118609, QN => n90392);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n118608, QN => n90393);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n118607, QN => n90394);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n118606, QN => n90395);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n118605, QN => n90396);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n118604, QN => n90397);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n118603, QN => n90398);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n118602, QN => n90399);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n118601, QN => n90400);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n118600, QN => n90401);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n118599, QN => n90402);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n118598, QN => n90403);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n118597, QN => n90404);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n118596, QN => n90405);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n118595, QN => n90406);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n118594, QN => n90407);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n118593, QN => n90408);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n118592, QN => n90409);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n118591, QN => n90410);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n118590, QN => n90411);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n118589, QN => n90412);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n118588, QN => n90413);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n118587, QN => n90414);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n118586, QN => n90415);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n118585, QN => n90416);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n118584, QN => n90417);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n118583, QN => n90418);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n118582, QN => n90419);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n118581, QN => n90420);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n118580, QN => n90421);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n118579, QN => n90422);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n118578, QN => n90423);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n118577, QN => n90424);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n118576, QN => n90425);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n118575, QN => n90426);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n118574, QN => n90427);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n118573, QN => n90428);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n118572, QN => n90429);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n118571, QN => n90430);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n118570, QN => n90431);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n118569, QN => n90432);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n118568, QN => n90433);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n118567, QN => n90434);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n118566, QN => n90435);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n118565, QN => n90436);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n118564, QN => n90437);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n110478, QN => n90311);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n110477, QN => n90312);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n110476, QN => n90313);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n110475, QN => n90314);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n110474, QN => n90315);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n110473, QN => n90316);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n110472, QN => n90317);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n110471, QN => n90318);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n110470, QN => n90319);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n110469, QN => n90320);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n110468, QN => n90321);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n110467, QN => n90322);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n110466, QN => n90323);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n110465, QN => n90324);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n110464, QN => n90325);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n110463, QN => n90326);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n110462, QN => n90327);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n110461, QN => n90328);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n110460, QN => n90329);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n110459, QN => n90330);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n110458, QN => n90331);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n110457, QN => n90332);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n110456, QN => n90333);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n110455, QN => n90334);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n110454, QN => n90335);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n110453, QN => n90336);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n110452, QN => n90337);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n110451, QN => n90338);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n110450, QN => n90339);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n110449, QN => n90340);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n110448, QN => n90341);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n110447, QN => n90342);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n110446, QN => n90343);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n110445, QN => n90344);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n110444, QN => n90345);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n110443, QN => n90346);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n110442, QN => n90347);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n110441, QN => n90348);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n110440, QN => n90349);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n110439, QN => n90350);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n110438, QN => n90351);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n110437, QN => n90352);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n110436, QN => n90353);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n110435, QN => n90354);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n110434, QN => n90355);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n110433, QN => n90356);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n110432, QN => n90357);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n110431, QN => n90358);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n110491, QN => n90359);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n110490, QN => n90360);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n110489, QN => n90361);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => 
                           n110488, QN => n90362);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => 
                           n110487, QN => n90363);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => 
                           n110546, QN => n90364);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => 
                           n110545, QN => n90365);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => 
                           n110544, QN => n90366);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => 
                           n110543, QN => n90367);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => 
                           n110542, QN => n90368);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => 
                           n110541, QN => n90369);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => 
                           n110540, QN => n90370);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n118857, QN => n90517);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n118856, QN => n90518);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n118855, QN => n90519);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n118854, QN => n90520);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n118853, QN => n90521);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n118852, QN => n90522);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n118851, QN => n90523);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n118850, QN => n90524);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n118849, QN => n90525);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n118848, QN => n90526);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n118847, QN => n90527);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n118846, QN => n90528);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n118845, QN => n90529);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n118844, QN => n90530);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n118843, QN => n90531);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n118842, QN => n90532);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n118841, QN => n90533);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n118840, QN => n90534);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n118839, QN => n90535);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n118838, QN => n90536);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n118837, QN => n90537);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n118836, QN => n90538);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n118835, QN => n90539);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n118834, QN => n90540);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n118833, QN => n90541);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n118832, QN => n90542);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n118831, QN => n90543);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n118830, QN => n90544);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n118829, QN => n90545);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n118828, QN => n90546);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n118827, QN => n90547);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n118826, QN => n90548);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n118825, QN => n90549);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n118824, QN => n90550);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n118823, QN => n90551);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n118822, QN => n90552);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n118821, QN => n90553);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n118820, QN => n90554);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n118819, QN => n90555);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n118818, QN => n90556);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n118817, QN => n90557);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => 
                           n110874, QN => n99914);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => 
                           n110873, QN => n99916);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => 
                           n110872, QN => n99917);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => 
                           n110871, QN => n99918);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => 
                           n119049, QN => n99716);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => 
                           n119048, QN => n99718);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n119047, QN => n99719);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => 
                           n119046, QN => n99720);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n118722, QN => n99446);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n118721, QN => n99448);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n118720, QN => n99449);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n118719, QN => n99450);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n103739, QN => n99580);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n103738, QN => n99582);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n103737, QN => n99583);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n103736, QN => n99584);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => 
                           n110192, QN => n98648);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => 
                           n110191, QN => n98650);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => 
                           n110190, QN => n98651);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => 
                           n110189, QN => n98652);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => 
                           n110486, QN => n98714);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => 
                           n110485, QN => n98716);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => 
                           n110484, QN => n98717);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => 
                           n110483, QN => n98718);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => 
                           n119177, QN => n99245);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n119176, QN => n99247);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n119175, QN => n99248);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n119174, QN => n99249);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => 
                           n119354, QN => n99113);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n119353, QN => n99115);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n119352, QN => n99116);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n119351, QN => n99117);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => 
                           n110863, QN => n99919);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => 
                           n110862, QN => n99920);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => 
                           n110861, QN => n99921);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => 
                           n110860, QN => n99922);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => 
                           n110859, QN => n99923);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => 
                           n110858, QN => n99924);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => 
                           n110857, QN => n99925);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => 
                           n110856, QN => n99926);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => 
                           n110855, QN => n99927);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => 
                           n110854, QN => n99928);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => 
                           n110853, QN => n99929);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => 
                           n110852, QN => n99930);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => 
                           n110851, QN => n99931);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => 
                           n110850, QN => n99932);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => 
                           n110849, QN => n99933);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => 
                           n110848, QN => n99934);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => 
                           n110847, QN => n99935);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => 
                           n110846, QN => n99936);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n5608, CK => CLK, Q => 
                           n110845, QN => n99937);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n5607, CK => CLK, Q => 
                           n110844, QN => n99938);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n5606, CK => CLK, Q => 
                           n110843, QN => n99939);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n5605, CK => CLK, Q => 
                           n110842, QN => n99940);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n5604, CK => CLK, Q => 
                           n110841, QN => n99941);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n5603, CK => CLK, Q => 
                           n110840, QN => n99942);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n5602, CK => CLK, Q => 
                           n110839, QN => n99943);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n5601, CK => CLK, Q => 
                           n110838, QN => n99944);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n5600, CK => CLK, Q => 
                           n110837, QN => n99945);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n5599, CK => CLK, Q => 
                           n110836, QN => n99946);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n5598, CK => CLK, Q => 
                           n110835, QN => n99947);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n5597, CK => CLK, Q => 
                           n110834, QN => n99948);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n5596, CK => CLK, Q => 
                           n110833, QN => n99949);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n5595, CK => CLK, Q => 
                           n110832, QN => n99950);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n5594, CK => CLK, Q => 
                           n110831, QN => n99951);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n5593, CK => CLK, Q => 
                           n110830, QN => n99952);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n5592, CK => CLK, Q => 
                           n110829, QN => n99953);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n5591, CK => CLK, Q => 
                           n110828, QN => n99954);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n5590, CK => CLK, Q => 
                           n110827, QN => n99955);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n5589, CK => CLK, Q => 
                           n110826, QN => n99956);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n5588, CK => CLK, Q => 
                           n110825, QN => n99957);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n5587, CK => CLK, Q => 
                           n110824, QN => n99958);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n5586, CK => CLK, Q => 
                           n110823, QN => n99959);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n5585, CK => CLK, Q => 
                           n110822, QN => n99960);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n5584, CK => CLK, Q => 
                           n110821, QN => n99961);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n5583, CK => CLK, Q => 
                           n110820, QN => n99962);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n5582, CK => CLK, Q => 
                           n110819, QN => n99963);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n5581, CK => CLK, Q => 
                           n110818, QN => n99964);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n5580, CK => CLK, Q => 
                           n110817, QN => n99965);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n5579, CK => CLK, Q => 
                           n110816, QN => n99966);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n5578, CK => CLK, Q => 
                           n110815, QN => n99967);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n5577, CK => CLK, Q => 
                           n110814, QN => n99968);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n5576, CK => CLK, Q => 
                           n110813, QN => n99969);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n5575, CK => CLK, Q => 
                           n110812, QN => n99970);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n5574, CK => CLK, Q => 
                           n110811, QN => n99971);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n5573, CK => CLK, Q => 
                           n110870, QN => n99972);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n5572, CK => CLK, Q => 
                           n110869, QN => n99973);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n5571, CK => CLK, Q => 
                           n110868, QN => n99974);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n5570, CK => CLK, Q => 
                           n110867, QN => n99975);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n5569, CK => CLK, Q => 
                           n110866, QN => n99976);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n5568, CK => CLK, Q => 
                           n110865, QN => n99977);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n5567, CK => CLK, Q => 
                           n110864, QN => n99978);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n119063, QN => n99721);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => 
                           n119062, QN => n99722);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n119061, QN => n99723);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => 
                           n119060, QN => n99724);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n119059, QN => n99725);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => 
                           n119058, QN => n99726);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n119057, QN => n99727);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => 
                           n119056, QN => n99728);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n119055, QN => n99729);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => 
                           n119054, QN => n99730);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n119053, QN => n99731);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => 
                           n119052, QN => n99732);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n119051, QN => n99733);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => 
                           n119050, QN => n99734);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n119109, QN => n99735);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => 
                           n119108, QN => n99736);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n119107, QN => n99737);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => 
                           n119106, QN => n99738);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n119105, QN => n99739);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => 
                           n119104, QN => n99740);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n119103, QN => n99741);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => 
                           n119102, QN => n99742);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n119101, QN => n99743);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => 
                           n119100, QN => n99744);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n119099, QN => n99745);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => 
                           n119098, QN => n99746);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n119097, QN => n99747);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => 
                           n119096, QN => n99748);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n119095, QN => n99749);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => 
                           n119094, QN => n99750);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n119093, QN => n99751);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => 
                           n119092, QN => n99752);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n119091, QN => n99753);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => 
                           n119090, QN => n99754);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n119089, QN => n99755);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => 
                           n119088, QN => n99756);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n119087, QN => n99757);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => 
                           n119086, QN => n99758);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n119085, QN => n99759);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => 
                           n119084, QN => n99760);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n119083, QN => n99761);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => 
                           n119082, QN => n99762);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n119081, QN => n99763);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => 
                           n119080, QN => n99764);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n119079, QN => n99765);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => 
                           n119078, QN => n99766);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n119077, QN => n99767);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => 
                           n119076, QN => n99768);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n119075, QN => n99769);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => 
                           n119074, QN => n99770);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => 
                           n119073, QN => n99771);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => 
                           n119072, QN => n99772);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => 
                           n119071, QN => n99773);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => 
                           n119070, QN => n99774);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => 
                           n119069, QN => n99775);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => 
                           n119068, QN => n99776);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => 
                           n119067, QN => n99777);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => 
                           n119066, QN => n99778);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => 
                           n119065, QN => n99779);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => 
                           n119064, QN => n99780);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n118623, QN => n99451);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n118622, QN => n99452);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n118621, QN => n99453);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n118620, QN => n99454);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n118619, QN => n99455);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n118618, QN => n99456);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n118617, QN => n99457);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n118616, QN => n99458);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n118615, QN => n99459);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n118614, QN => n99460);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n118613, QN => n99461);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n118612, QN => n99462);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n118611, QN => n99463);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n118610, QN => n99464);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n118657, QN => n99465);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n118656, QN => n99466);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n118655, QN => n99467);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n118654, QN => n99468);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n118653, QN => n99469);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n118652, QN => n99470);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n118651, QN => n99471);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n118650, QN => n99472);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n118649, QN => n99473);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n118648, QN => n99474);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n118647, QN => n99475);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n118646, QN => n99476);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n118645, QN => n99477);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n118644, QN => n99478);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n118643, QN => n99479);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n118642, QN => n99480);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n118641, QN => n99481);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n118640, QN => n99482);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n118639, QN => n99483);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n118638, QN => n99484);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n118637, QN => n99485);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n118636, QN => n99486);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n118635, QN => n99487);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n118634, QN => n99488);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n118633, QN => n99489);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n118632, QN => n99490);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n118631, QN => n99491);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n118630, QN => n99492);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n118629, QN => n99493);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n118628, QN => n99494);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n118627, QN => n99495);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n118626, QN => n99496);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n118625, QN => n99497);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n118624, QN => n99498);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n118669, QN => n99499);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n118668, QN => n99500);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n118667, QN => n99501);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => 
                           n118666, QN => n99502);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => 
                           n118665, QN => n99503);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => 
                           n118664, QN => n99504);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => 
                           n118663, QN => n99505);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => 
                           n118662, QN => n99506);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => 
                           n118661, QN => n99507);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => 
                           n118660, QN => n99508);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => 
                           n118659, QN => n99509);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => 
                           n118658, QN => n99510);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n103611, QN => n99585);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n103610, QN => n99586);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n103609, QN => n99587);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n103608, QN => n99588);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n103607, QN => n99589);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n103606, QN => n99590);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n103605, QN => n99591);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n103604, QN => n99592);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n103603, QN => n99593);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n103602, QN => n99594);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n103601, QN => n99595);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n103600, QN => n99596);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n103599, QN => n99597);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n103598, QN => n99598);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n103597, QN => n99599);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n103596, QN => n99600);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n103595, QN => n99601);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n103594, QN => n99602);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n103593, QN => n99603);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n103592, QN => n99604);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n103591, QN => n99605);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n103590, QN => n99606);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n103589, QN => n99607);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n103588, QN => n99608);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n103587, QN => n99609);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n103586, QN => n99610);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n103585, QN => n99611);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n103584, QN => n99612);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n103583, QN => n99613);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n103582, QN => n99614);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n103581, QN => n99615);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n103580, QN => n99616);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n103579, QN => n99617);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n103578, QN => n99618);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n103577, QN => n99619);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n103576, QN => n99620);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n103575, QN => n99621);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n103574, QN => n99622);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n103573, QN => n99623);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n103572, QN => n99624);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n103571, QN => n99625);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n103570, QN => n99626);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n103569, QN => n99627);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n103568, QN => n99628);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n103567, QN => n99629);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n103566, QN => n99630);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n103565, QN => n99631);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n103564, QN => n99632);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n103563, QN => n99633);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n103562, QN => n99634);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n103561, QN => n99635);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => 
                           n103560, QN => n99636);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => 
                           n103559, QN => n99637);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => 
                           n103558, QN => n99638);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => 
                           n103557, QN => n99639);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n103556, QN => n99640);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n103555, QN => n99641);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => 
                           n103554, QN => n99642);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => 
                           n103553, QN => n99643);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => 
                           n103552, QN => n99644);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => 
                           n110580, QN => n99047);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n110579, QN => n99049);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n110578, QN => n99050);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n110577, QN => n99051);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => 
                           n119301, QN => n99311);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n119300, QN => n99313);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n119299, QN => n99314);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n119298, QN => n99315);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n119113, QN => n99179);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n119112, QN => n99181);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n119111, QN => n99182);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n119110, QN => n99183);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => 
                           n118910, QN => n98586);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => 
                           n118909, QN => n98587);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => 
                           n118908, QN => n98588);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => 
                           n118907, QN => n98589);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => 
                           n118906, QN => n98590);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => 
                           n118905, QN => n98591);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => 
                           n118904, QN => n98592);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => 
                           n118903, QN => n98593);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => 
                           n118902, QN => n98594);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => 
                           n118901, QN => n98595);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => 
                           n118900, QN => n98596);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => 
                           n118899, QN => n98597);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => 
                           n118898, QN => n98598);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => 
                           n118897, QN => n98599);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => 
                           n118896, QN => n98600);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => 
                           n118895, QN => n98601);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => 
                           n118894, QN => n98602);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => 
                           n118893, QN => n98603);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => 
                           n118892, QN => n98604);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => 
                           n118891, QN => n98605);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => 
                           n118890, QN => n98606);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => 
                           n118889, QN => n98607);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => 
                           n118888, QN => n98608);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => 
                           n118887, QN => n98609);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => 
                           n118886, QN => n98610);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => 
                           n118885, QN => n98611);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => 
                           n118884, QN => n98612);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => 
                           n118883, QN => n98613);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => 
                           n118882, QN => n98614);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => 
                           n118881, QN => n98615);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => 
                           n118880, QN => n98616);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => 
                           n118879, QN => n98617);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => 
                           n118878, QN => n98618);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => 
                           n118877, QN => n98619);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => 
                           n118876, QN => n98620);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => 
                           n118875, QN => n98621);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => 
                           n118874, QN => n98622);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => 
                           n118873, QN => n98623);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => 
                           n118872, QN => n98624);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => 
                           n118871, QN => n98625);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => 
                           n118870, QN => n98626);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => 
                           n118869, QN => n98627);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => 
                           n118868, QN => n98628);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => 
                           n118867, QN => n98629);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => 
                           n118866, QN => n98630);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => 
                           n118865, QN => n98631);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => 
                           n118864, QN => n98632);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => 
                           n118863, QN => n98633);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => 
                           n118862, QN => n98634);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => 
                           n118914, QN => n98635);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => 
                           n118913, QN => n98636);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => 
                           n118912, QN => n98637);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => 
                           n118911, QN => n98638);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => 
                           n118921, QN => n98639);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => 
                           n118920, QN => n98640);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => 
                           n118919, QN => n98641);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => 
                           n118918, QN => n98642);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => 
                           n118917, QN => n98643);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => 
                           n118916, QN => n98644);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => 
                           n118915, QN => n98645);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => 
                           n110184, QN => n98653);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => 
                           n110183, QN => n98654);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => 
                           n110182, QN => n98655);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => 
                           n110181, QN => n98656);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => 
                           n110180, QN => n98657);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => 
                           n110179, QN => n98658);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => 
                           n110178, QN => n98659);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => 
                           n110177, QN => n98660);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => 
                           n110176, QN => n98661);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => 
                           n110175, QN => n98662);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => 
                           n110174, QN => n98663);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => 
                           n110173, QN => n98664);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => 
                           n110172, QN => n98665);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => 
                           n110171, QN => n98666);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => 
                           n110234, QN => n98667);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => 
                           n110233, QN => n98668);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => 
                           n110232, QN => n98669);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => 
                           n110231, QN => n98670);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => 
                           n110230, QN => n98671);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => 
                           n110229, QN => n98672);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => 
                           n110228, QN => n98673);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => 
                           n110227, QN => n98674);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => 
                           n110226, QN => n98675);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => 
                           n110225, QN => n98676);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => 
                           n110224, QN => n98677);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => 
                           n110223, QN => n98678);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => 
                           n110222, QN => n98679);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => 
                           n110221, QN => n98680);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => 
                           n110220, QN => n98681);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => 
                           n110219, QN => n98682);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => 
                           n110218, QN => n98683);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => 
                           n110217, QN => n98684);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => 
                           n110216, QN => n98685);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => 
                           n110215, QN => n98686);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => 
                           n110214, QN => n98687);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => 
                           n110213, QN => n98688);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => 
                           n110212, QN => n98689);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => 
                           n110211, QN => n98690);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => 
                           n110210, QN => n98691);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => 
                           n110209, QN => n98692);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => 
                           n110208, QN => n98693);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => 
                           n110207, QN => n98694);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => 
                           n110206, QN => n98695);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => 
                           n110205, QN => n98696);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => 
                           n110204, QN => n98697);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => 
                           n110203, QN => n98698);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => 
                           n110202, QN => n98699);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => 
                           n110201, QN => n98700);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => 
                           n110200, QN => n98701);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => 
                           n110199, QN => n98702);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => 
                           n110198, QN => n98703);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => 
                           n110197, QN => n98704);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => 
                           n110196, QN => n98705);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => 
                           n110195, QN => n98706);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => 
                           n110194, QN => n98707);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => 
                           n110193, QN => n98708);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => 
                           n110188, QN => n98709);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => 
                           n110187, QN => n98710);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => 
                           n110186, QN => n98711);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => 
                           n110185, QN => n98712);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => 
                           n118545, QN => n98523);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => 
                           n118544, QN => n98524);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => 
                           n118543, QN => n98525);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => 
                           n118542, QN => n98526);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => 
                           n118541, QN => n98527);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => 
                           n118540, QN => n98528);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => 
                           n118539, QN => n98529);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => 
                           n118538, QN => n98530);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => 
                           n118537, QN => n98531);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => 
                           n118536, QN => n98532);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => 
                           n118535, QN => n98533);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => 
                           n118534, QN => n98534);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => 
                           n118533, QN => n98535);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => 
                           n118532, QN => n98536);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => 
                           n118531, QN => n98537);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => 
                           n118530, QN => n98538);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => 
                           n118529, QN => n98539);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => 
                           n118528, QN => n98540);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => 
                           n118527, QN => n98541);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => 
                           n118526, QN => n98542);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => 
                           n118525, QN => n98543);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => 
                           n118524, QN => n98544);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => 
                           n118523, QN => n98545);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => 
                           n118522, QN => n98546);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => 
                           n118521, QN => n98547);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => 
                           n118520, QN => n98548);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => 
                           n118519, QN => n98549);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => 
                           n118518, QN => n98550);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => 
                           n118517, QN => n98551);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => 
                           n118516, QN => n98552);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => 
                           n118515, QN => n98553);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => 
                           n118514, QN => n98554);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => 
                           n118513, QN => n98555);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => 
                           n118512, QN => n98556);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => 
                           n118511, QN => n98557);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => 
                           n118510, QN => n98558);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => 
                           n118509, QN => n98559);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => 
                           n118508, QN => n98560);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => 
                           n118507, QN => n98561);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => 
                           n118506, QN => n98562);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => 
                           n118505, QN => n98563);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => 
                           n118805, QN => n98564);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => 
                           n118804, QN => n98565);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => 
                           n118803, QN => n98566);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => 
                           n118802, QN => n98567);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => 
                           n118801, QN => n98568);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => 
                           n118800, QN => n98569);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => 
                           n118799, QN => n98570);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => 
                           n118798, QN => n98571);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => 
                           n118809, QN => n98572);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => 
                           n118808, QN => n98573);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => 
                           n118807, QN => n98574);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => 
                           n118806, QN => n98575);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => 
                           n118816, QN => n98576);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => 
                           n118815, QN => n98577);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => 
                           n118814, QN => n98578);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => 
                           n118813, QN => n98579);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => 
                           n118812, QN => n98580);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => 
                           n118811, QN => n98581);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => 
                           n118810, QN => n98582);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n118751, QN => n98848);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n118750, QN => n98849);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n118749, QN => n98850);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n118748, QN => n98851);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n118747, QN => n98852);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n118746, QN => n98853);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n118745, QN => n98854);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n118744, QN => n98855);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n118743, QN => n98856);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n118742, QN => n98857);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n118741, QN => n98858);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n118740, QN => n98859);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n118739, QN => n98860);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n118738, QN => n98861);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n118797, QN => n98862);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n118796, QN => n98863);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n118795, QN => n98864);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n118794, QN => n98865);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n118793, QN => n98866);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n118792, QN => n98867);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           n118791, QN => n98868);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           n118790, QN => n98869);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           n118789, QN => n98870);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           n118788, QN => n98871);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           n118787, QN => n98872);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => 
                           n118786, QN => n98873);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           n118785, QN => n98874);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           n118784, QN => n98875);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => 
                           n118783, QN => n98876);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n118782, QN => n98877);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n118781, QN => n98878);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n118780, QN => n98879);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n118779, QN => n98880);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n118778, QN => n98881);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n118777, QN => n98882);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n118776, QN => n98883);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n118775, QN => n98884);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n118774, QN => n98885);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n118773, QN => n98886);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n118772, QN => n98887);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => 
                           n118771, QN => n98888);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => 
                           n118770, QN => n98889);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => 
                           n118769, QN => n98890);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => 
                           n118768, QN => n98891);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => 
                           n118767, QN => n98892);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => 
                           n118766, QN => n98893);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => 
                           n118765, QN => n98894);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => 
                           n118764, QN => n98895);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => 
                           n118763, QN => n98896);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => 
                           n118762, QN => n98897);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => 
                           n118761, QN => n98898);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => 
                           n118760, QN => n98899);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => 
                           n118759, QN => n98900);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => 
                           n118758, QN => n98901);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => 
                           n118757, QN => n98902);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => 
                           n118756, QN => n98903);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => 
                           n118755, QN => n98904);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => 
                           n118754, QN => n98905);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => 
                           n118753, QN => n98906);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => 
                           n118752, QN => n98907);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => 
                           n118970, QN => n98986);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => 
                           n118969, QN => n98987);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => 
                           n118968, QN => n98988);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => 
                           n118967, QN => n98989);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => 
                           n118966, QN => n98990);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => 
                           n118965, QN => n98991);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => 
                           n118964, QN => n98992);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => 
                           n118963, QN => n98993);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => 
                           n118962, QN => n98994);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => 
                           n118961, QN => n98995);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => 
                           n118960, QN => n98996);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => 
                           n118959, QN => n98997);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => 
                           n118958, QN => n98998);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => 
                           n118957, QN => n98999);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => 
                           n118956, QN => n99000);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => 
                           n118955, QN => n99001);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => 
                           n118954, QN => n99002);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => 
                           n118953, QN => n99003);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => 
                           n118952, QN => n99004);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => 
                           n118951, QN => n99005);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => 
                           n118950, QN => n99006);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => 
                           n118949, QN => n99007);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => 
                           n118948, QN => n99008);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => 
                           n118947, QN => n99009);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => 
                           n118946, QN => n99010);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => 
                           n118945, QN => n99011);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => 
                           n118944, QN => n99012);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => 
                           n118943, QN => n99013);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => 
                           n118942, QN => n99014);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => 
                           n118941, QN => n99015);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => 
                           n118940, QN => n99016);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => 
                           n118939, QN => n99017);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => 
                           n118938, QN => n99018);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => 
                           n118937, QN => n99019);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => 
                           n118936, QN => n99020);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => 
                           n118935, QN => n99021);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => 
                           n118934, QN => n99022);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => 
                           n118933, QN => n99023);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => 
                           n118932, QN => n99024);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => 
                           n118931, QN => n99025);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => 
                           n118930, QN => n99026);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => 
                           n118929, QN => n99027);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => 
                           n118928, QN => n99028);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => 
                           n118927, QN => n99029);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => 
                           n118926, QN => n99030);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => 
                           n118925, QN => n99031);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => 
                           n118924, QN => n99032);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => 
                           n118923, QN => n99033);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => 
                           n118922, QN => n99034);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => 
                           n118974, QN => n99035);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => 
                           n118973, QN => n99036);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => 
                           n118972, QN => n99037);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => 
                           n118971, QN => n99038);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => 
                           n118981, QN => n99039);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => 
                           n118980, QN => n99040);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => 
                           n118979, QN => n99041);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => 
                           n118978, QN => n99042);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => 
                           n118977, QN => n99043);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => 
                           n118976, QN => n99044);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => 
                           n118975, QN => n99045);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => 
                           n110539, QN => n98719);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => 
                           n110538, QN => n98720);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => 
                           n110537, QN => n98721);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => 
                           n110536, QN => n98722);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => 
                           n110535, QN => n98723);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => 
                           n110534, QN => n98724);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => 
                           n110533, QN => n98725);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => 
                           n110532, QN => n98726);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => 
                           n110531, QN => n98727);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => 
                           n110530, QN => n98728);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => 
                           n110529, QN => n98729);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => 
                           n110528, QN => n98730);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => 
                           n110527, QN => n98731);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => 
                           n110526, QN => n98732);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => 
                           n110525, QN => n98733);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => 
                           n110524, QN => n98734);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => 
                           n110523, QN => n98735);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => 
                           n110522, QN => n98736);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => 
                           n110521, QN => n98737);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => 
                           n110520, QN => n98738);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => 
                           n110519, QN => n98739);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => 
                           n110518, QN => n98740);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => 
                           n110517, QN => n98741);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => 
                           n110516, QN => n98742);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n7202, CK => CLK, Q => 
                           n110515, QN => n98743);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => 
                           n110514, QN => n98744);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => 
                           n110513, QN => n98745);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => 
                           n110512, QN => n98746);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => 
                           n110511, QN => n98747);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => 
                           n110510, QN => n98748);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => 
                           n110509, QN => n98749);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => 
                           n110508, QN => n98750);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => 
                           n110507, QN => n98751);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => 
                           n110506, QN => n98752);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => 
                           n110505, QN => n98753);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => 
                           n110504, QN => n98754);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => 
                           n110503, QN => n98755);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => 
                           n110502, QN => n98756);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => 
                           n110501, QN => n98757);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => 
                           n110500, QN => n98758);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => 
                           n110499, QN => n98759);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => 
                           n110498, QN => n98760);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => 
                           n110497, QN => n98761);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => 
                           n110496, QN => n98762);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => 
                           n110495, QN => n98763);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => 
                           n110494, QN => n98764);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => 
                           n110493, QN => n98765);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => 
                           n110492, QN => n98766);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => 
                           n110551, QN => n98767);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => 
                           n110550, QN => n98768);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => 
                           n110549, QN => n98769);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => 
                           n110548, QN => n98770);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => 
                           n110547, QN => n98771);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => 
                           n110558, QN => n98772);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => 
                           n110557, QN => n98773);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => 
                           n110556, QN => n98774);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => 
                           n110555, QN => n98775);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => 
                           n110554, QN => n98776);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => 
                           n110553, QN => n98777);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => 
                           n110552, QN => n98778);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n119191, QN => n99250);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n119190, QN => n99251);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n119189, QN => n99252);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n119188, QN => n99253);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n119187, QN => n99254);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n119186, QN => n99255);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n119185, QN => n99256);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n119184, QN => n99257);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n119183, QN => n99258);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n119182, QN => n99259);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n119181, QN => n99260);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n119180, QN => n99261);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n119179, QN => n99262);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n119178, QN => n99263);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n119237, QN => n99264);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n119236, QN => n99265);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n119235, QN => n99266);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n119234, QN => n99267);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n119233, QN => n99268);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => 
                           n119232, QN => n99269);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => 
                           n119231, QN => n99270);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => 
                           n119230, QN => n99271);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => 
                           n119229, QN => n99272);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => 
                           n119228, QN => n99273);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => 
                           n119227, QN => n99274);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => 
                           n119226, QN => n99275);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => 
                           n119225, QN => n99276);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => 
                           n119224, QN => n99277);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => 
                           n119223, QN => n99278);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n119222, QN => n99279);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n119221, QN => n99280);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n119220, QN => n99281);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n119219, QN => n99282);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n119218, QN => n99283);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n119217, QN => n99284);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n119216, QN => n99285);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n119215, QN => n99286);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n119214, QN => n99287);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n119213, QN => n99288);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n119212, QN => n99289);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n119211, QN => n99290);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n119210, QN => n99291);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n119209, QN => n99292);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n119208, QN => n99293);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n119207, QN => n99294);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n119206, QN => n99295);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n119205, QN => n99296);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n119204, QN => n99297);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n119203, QN => n99298);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n119202, QN => n99299);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n119201, QN => n99300);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => 
                           n119200, QN => n99301);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => 
                           n119199, QN => n99302);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => 
                           n119198, QN => n99303);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => 
                           n119197, QN => n99304);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => 
                           n119196, QN => n99305);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => 
                           n119195, QN => n99306);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => 
                           n119194, QN => n99307);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => 
                           n119193, QN => n99308);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => 
                           n119192, QN => n99309);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n119350, QN => n99118);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n119349, QN => n99119);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n119348, QN => n99120);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n119347, QN => n99121);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n119346, QN => n99122);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n119345, QN => n99123);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n119344, QN => n99124);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n119343, QN => n99125);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n119342, QN => n99126);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n119341, QN => n99127);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n119340, QN => n99128);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n119339, QN => n99129);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n119338, QN => n99130);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n119337, QN => n99131);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n119336, QN => n99132);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n119335, QN => n99133);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n119334, QN => n99134);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n119333, QN => n99135);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n119332, QN => n99136);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n119331, QN => n99137);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n119330, QN => n99138);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n119329, QN => n99139);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n119328, QN => n99140);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n119327, QN => n99141);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n119326, QN => n99142);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n119325, QN => n99143);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n119324, QN => n99144);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n119323, QN => n99145);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n119322, QN => n99146);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n119321, QN => n99147);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n119320, QN => n99148);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n119319, QN => n99149);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n119318, QN => n99150);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n119317, QN => n99151);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n119316, QN => n99152);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n119315, QN => n99153);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n119314, QN => n99154);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n119313, QN => n99155);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n119312, QN => n99156);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n119311, QN => n99157);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n119310, QN => n99158);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n119309, QN => n99159);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n119308, QN => n99160);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n119307, QN => n99161);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n119306, QN => n99162);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n119305, QN => n99163);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n119304, QN => n99164);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n119303, QN => n99165);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n119302, QN => n99166);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n119358, QN => n99167);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n119357, QN => n99168);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => 
                           n119356, QN => n99169);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => 
                           n119355, QN => n99170);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => 
                           n119365, QN => n99171);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => 
                           n119364, QN => n99172);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n119363, QN => n99173);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n119362, QN => n99174);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n119361, QN => n99175);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n119360, QN => n99176);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n119359, QN => n99177);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n110572, QN => n99052);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n110571, QN => n99053);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n110570, QN => n99054);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n110569, QN => n99055);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n110568, QN => n99056);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n110567, QN => n99057);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n110566, QN => n99058);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n110565, QN => n99059);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n110564, QN => n99060);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n110563, QN => n99061);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n110562, QN => n99062);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n110561, QN => n99063);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n110560, QN => n99064);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n110559, QN => n99065);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n110622, QN => n99066);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n110621, QN => n99067);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n110620, QN => n99068);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n110619, QN => n99069);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n110618, QN => n99070);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n110617, QN => n99071);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n110616, QN => n99072);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n110615, QN => n99073);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n110614, QN => n99074);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n110613, QN => n99075);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n110612, QN => n99076);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n110611, QN => n99077);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n110610, QN => n99078);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n110609, QN => n99079);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n110608, QN => n99080);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n110607, QN => n99081);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n110606, QN => n99082);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n110605, QN => n99083);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n110604, QN => n99084);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n110603, QN => n99085);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n110602, QN => n99086);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n110601, QN => n99087);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n110600, QN => n99088);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n110599, QN => n99089);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n110598, QN => n99090);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n110597, QN => n99091);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n110596, QN => n99092);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n110595, QN => n99093);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n110594, QN => n99094);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n110593, QN => n99095);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n110592, QN => n99096);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n110591, QN => n99097);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n110590, QN => n99098);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n110589, QN => n99099);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n110588, QN => n99100);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n110587, QN => n99101);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n110586, QN => n99102);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => 
                           n110585, QN => n99103);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => 
                           n110584, QN => n99104);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => 
                           n110583, QN => n99105);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => 
                           n110582, QN => n99106);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => 
                           n110581, QN => n99107);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => 
                           n110576, QN => n99108);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => 
                           n110575, QN => n99109);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => 
                           n110574, QN => n99110);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => 
                           n110573, QN => n99111);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n119251, QN => n99316);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n119250, QN => n99317);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n119249, QN => n99318);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n119248, QN => n99319);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n119247, QN => n99320);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n119246, QN => n99321);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n119245, QN => n99322);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n119244, QN => n99323);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n119243, QN => n99324);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n119242, QN => n99325);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n119241, QN => n99326);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n119240, QN => n99327);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n119239, QN => n99328);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n119238, QN => n99329);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n119285, QN => n99330);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n119284, QN => n99331);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n119283, QN => n99332);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n119282, QN => n99333);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n119281, QN => n99334);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n119280, QN => n99335);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n119279, QN => n99336);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n119278, QN => n99337);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n119277, QN => n99338);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n119276, QN => n99339);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n119275, QN => n99340);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n119274, QN => n99341);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n119273, QN => n99342);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n119272, QN => n99343);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n119271, QN => n99344);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n119270, QN => n99345);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n119269, QN => n99346);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n119268, QN => n99347);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n119267, QN => n99348);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n119266, QN => n99349);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n119265, QN => n99350);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n119264, QN => n99351);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n119263, QN => n99352);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n119262, QN => n99353);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n119261, QN => n99354);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n119260, QN => n99355);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n119259, QN => n99356);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n119258, QN => n99357);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n119257, QN => n99358);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n119256, QN => n99359);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n119255, QN => n99360);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n119254, QN => n99361);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n119253, QN => n99362);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n119252, QN => n99363);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n119297, QN => n99364);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n119296, QN => n99365);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n119295, QN => n99366);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => 
                           n119294, QN => n99367);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => 
                           n119293, QN => n99368);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => 
                           n119292, QN => n99369);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => 
                           n119291, QN => n99370);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => 
                           n119290, QN => n99371);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => 
                           n119289, QN => n99372);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => 
                           n119288, QN => n99373);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => 
                           n119287, QN => n99374);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => 
                           n119286, QN => n99375);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n119127, QN => n99184);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n119126, QN => n99185);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n119125, QN => n99186);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n119124, QN => n99187);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n119123, QN => n99188);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n119122, QN => n99189);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n119121, QN => n99190);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n119120, QN => n99191);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n119119, QN => n99192);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n119118, QN => n99193);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n119117, QN => n99194);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n119116, QN => n99195);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n119115, QN => n99196);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n119114, QN => n99197);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n119173, QN => n99198);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n119172, QN => n99199);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n119171, QN => n99200);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n119170, QN => n99201);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n119169, QN => n99202);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n119168, QN => n99203);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n119167, QN => n99204);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n119166, QN => n99205);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n119165, QN => n99206);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n119164, QN => n99207);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n119163, QN => n99208);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n119162, QN => n99209);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n119161, QN => n99210);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n119160, QN => n99211);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n119159, QN => n99212);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n119158, QN => n99213);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n119157, QN => n99214);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n119156, QN => n99215);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n119155, QN => n99216);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n119154, QN => n99217);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n119153, QN => n99218);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n119152, QN => n99219);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n119151, QN => n99220);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n119150, QN => n99221);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n119149, QN => n99222);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n119148, QN => n99223);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n119147, QN => n99224);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n119146, QN => n99225);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n119145, QN => n99226);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n119144, QN => n99227);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n119143, QN => n99228);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n119142, QN => n99229);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n119141, QN => n99230);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n119140, QN => n99231);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n119139, QN => n99232);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n119138, QN => n99233);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n119137, QN => n99234);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => 
                           n119136, QN => n99235);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => 
                           n119135, QN => n99236);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => 
                           n119134, QN => n99237);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => 
                           n119133, QN => n99238);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => 
                           n119132, QN => n99239);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => 
                           n119131, QN => n99240);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => 
                           n119130, QN => n99241);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => 
                           n119129, QN => n99242);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => 
                           n119128, QN => n99243);
   OUT1_reg_3_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => OUT1_3_port, 
                           QN => n103051);
   OUT1_reg_2_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => OUT1_2_port, 
                           QN => n103050);
   OUT1_reg_1_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => OUT1_1_port, 
                           QN => n103049);
   OUT1_reg_0_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => OUT1_0_port, 
                           QN => n103048);
   OUT1_reg_59_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => OUT1_59_port
                           , QN => n103047);
   OUT1_reg_58_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => OUT1_58_port
                           , QN => n103046);
   OUT1_reg_57_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => OUT1_57_port
                           , QN => n103045);
   OUT1_reg_56_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => OUT1_56_port
                           , QN => n103044);
   OUT1_reg_55_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => OUT1_55_port
                           , QN => n103043);
   OUT1_reg_54_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => OUT1_54_port
                           , QN => n103042);
   OUT1_reg_53_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => OUT1_53_port
                           , QN => n103041);
   OUT1_reg_52_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => OUT1_52_port
                           , QN => n103040);
   OUT1_reg_51_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => OUT1_51_port
                           , QN => n103039);
   OUT1_reg_50_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => OUT1_50_port
                           , QN => n103038);
   OUT1_reg_49_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => OUT1_49_port
                           , QN => n103037);
   OUT1_reg_48_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => OUT1_48_port
                           , QN => n103036);
   OUT1_reg_47_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => OUT1_47_port
                           , QN => n103035);
   OUT1_reg_46_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => OUT1_46_port
                           , QN => n103034);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5340, CK => CLK, Q => OUT2_29_port
                           , QN => n110957);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5339, CK => CLK, Q => OUT2_28_port
                           , QN => n110956);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5338, CK => CLK, Q => OUT2_27_port
                           , QN => n110955);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5337, CK => CLK, Q => OUT2_26_port
                           , QN => n110954);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5336, CK => CLK, Q => OUT2_25_port
                           , QN => n110953);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5335, CK => CLK, Q => OUT2_24_port
                           , QN => n110952);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5334, CK => CLK, Q => OUT2_23_port
                           , QN => n110951);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5333, CK => CLK, Q => OUT2_22_port
                           , QN => n110950);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5332, CK => CLK, Q => OUT2_21_port
                           , QN => n110949);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5331, CK => CLK, Q => OUT2_20_port
                           , QN => n110948);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5330, CK => CLK, Q => OUT2_19_port
                           , QN => n110947);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5329, CK => CLK, Q => OUT2_18_port
                           , QN => n110946);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5328, CK => CLK, Q => OUT2_17_port
                           , QN => n110945);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5327, CK => CLK, Q => OUT2_16_port
                           , QN => n110944);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5326, CK => CLK, Q => OUT2_15_port
                           , QN => n110943);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5325, CK => CLK, Q => OUT2_14_port
                           , QN => n110942);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5324, CK => CLK, Q => OUT2_13_port
                           , QN => n110941);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5323, CK => CLK, Q => OUT2_12_port
                           , QN => n110940);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5322, CK => CLK, Q => OUT2_11_port
                           , QN => n110939);
   U81228 : NOR3_X2 port map( A1 => n120216, A2 => ADD_RD1(1), A3 => n116475, 
                           ZN => n116457);
   U81241 : NOR3_X2 port map( A1 => n120216, A2 => ADD_RD1(2), A3 => n116478, 
                           ZN => n116453);
   U83316 : NAND3_X1 port map( A1 => n113987, A2 => n113988, A3 => n113989, ZN 
                           => n113893);
   U83317 : NAND3_X1 port map( A1 => n113989, A2 => n113988, A3 => ADD_WR(0), 
                           ZN => n113901);
   U83318 : NAND3_X1 port map( A1 => n113989, A2 => n113987, A3 => ADD_WR(3), 
                           ZN => n114054);
   U83319 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n113989, A3 => ADD_WR(3),
                           ZN => n114121);
   U83320 : NAND3_X1 port map( A1 => n113987, A2 => n113988, A3 => n114302, ZN 
                           => n114141);
   U83321 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n113988, A3 => n114302, 
                           ZN => n114144);
   U83322 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n113987, A3 => n114302, 
                           ZN => n114371);
   U83323 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(0), A3 => n114302,
                           ZN => n114374);
   U83324 : NAND3_X1 port map( A1 => ENABLE, A2 => n120628, A3 => RD1, ZN => 
                           n114658);
   U83325 : NAND3_X1 port map( A1 => ENABLE, A2 => n120628, A3 => RD2, ZN => 
                           n116491);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => 
                           n95528, QN => n114644);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => 
                           n95527, QN => n114704);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => 
                           n95526, QN => n114730);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => 
                           n95525, QN => n114756);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n5566, CK => CLK, Q => 
                           n117996, QN => n114578);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n5565, CK => CLK, Q => 
                           n117995, QN => n114580);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n5564, CK => CLK, Q => 
                           n117994, QN => n114581);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n5563, CK => CLK, Q => 
                           n117993, QN => n114582);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => 
                           n119843, QN => n114510);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n119842, QN => n114512);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => 
                           n119841, QN => n114513);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n119840, QN => n114514);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => 
                           n119839, QN => n114444);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => 
                           n119838, QN => n114446);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => 
                           n119837, QN => n114447);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n119836, QN => n114448);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => 
                           n119835, QN => n114378);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => 
                           n119834, QN => n114380);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n119833, QN => n114381);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => 
                           n119832, QN => n114382);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => 
                           n117988, QN => n114306);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n117987, QN => n114308);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n117986, QN => n114309);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n117985, QN => n114310);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n117984, QN => n114235);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n117983, QN => n114237);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n117982, QN => n114238);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n117981, QN => n114239);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n119831, QN => n114146);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n119830, QN => n114148);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n119829, QN => n114149);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n119828, QN => n114150);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => 
                           n109906, QN => n113903);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => 
                           n109905, QN => n113905);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => 
                           n109904, QN => n113906);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => 
                           n109903, QN => n113907);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => 
                           n111048, QN => n113981);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => 
                           n111047, QN => n113983);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n111046, QN => n113984);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n111045, QN => n113985);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n7422, CK => CLK, Q => 
                           n109898, QN => n113896);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n7421, CK => CLK, Q => 
                           n109897, QN => n113898);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => 
                           n109896, QN => n113899);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => 
                           n109895, QN => n113900);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => 
                           n111044, QN => n114123);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => 
                           n111043, QN => n114125);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => 
                           n111042, QN => n114126);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => 
                           n111041, QN => n114127);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n109997, QN => n114215);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n109996, QN => n114216);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n109995, QN => n114217);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n109994, QN => n114218);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n109993, QN => n114219);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n109992, QN => n114220);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => 
                           n109991, QN => n114221);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => 
                           n109990, QN => n114222);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => 
                           n109989, QN => n114223);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n109988, QN => n114224);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n109987, QN => n114225);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n109986, QN => n114226);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n109985, QN => n114227);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n109984, QN => n114228);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n109983, QN => n114229);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n109982, QN => n114230);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n109981, QN => n114231);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n109980, QN => n114232);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n109979, QN => n114233);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => 
                           n119827, QN => n113915);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => 
                           n119826, QN => n113917);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => 
                           n119825, QN => n113918);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => 
                           n119824, QN => n113919);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => 
                           n95488, QN => n114782);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => 
                           n95487, QN => n114810);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => 
                           n95486, QN => n114838);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => 
                           n95485, QN => n114866);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => 
                           n95484, QN => n114894);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => 
                           n95483, QN => n114922);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => 
                           n95482, QN => n114950);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => 
                           n95481, QN => n114978);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => 
                           n95480, QN => n115006);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => 
                           n95479, QN => n115034);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => 
                           n95478, QN => n115062);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => 
                           n95477, QN => n115090);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => 
                           n95476, QN => n115118);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => 
                           n95475, QN => n115146);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => 
                           n95474, QN => n115174);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => 
                           n95473, QN => n115202);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => 
                           n95472, QN => n115230);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => 
                           n95471, QN => n115258);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => 
                           n95470, QN => n115286);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => 
                           n95469, QN => n115314);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => 
                           n95468, QN => n115342);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => 
                           n95467, QN => n115370);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => 
                           n95466, QN => n115398);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => 
                           n95465, QN => n115426);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => 
                           n95464, QN => n115454);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => 
                           n95463, QN => n115482);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => 
                           n95462, QN => n115510);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => 
                           n95461, QN => n115538);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => 
                           n95460, QN => n115566);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => 
                           n95459, QN => n115594);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => 
                           n95458, QN => n115622);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => 
                           n95457, QN => n115650);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => 
                           n95456, QN => n115678);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => 
                           n95455, QN => n115706);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => 
                           n95454, QN => n115734);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => 
                           n95453, QN => n115762);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => 
                           n95452, QN => n115790);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => 
                           n95451, QN => n115818);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => 
                           n95450, QN => n115846);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => 
                           n95449, QN => n115874);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => 
                           n95448, QN => n115902);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => 
                           n95447, QN => n115930);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => 
                           n95446, QN => n115958);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => 
                           n95445, QN => n115986);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => 
                           n95444, QN => n116014);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => 
                           n95443, QN => n116042);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => 
                           n95442, QN => n116070);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => 
                           n95441, QN => n116098);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => 
                           n95440, QN => n116126);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => 
                           n95439, QN => n116154);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => 
                           n95438, QN => n116182);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => 
                           n95437, QN => n116210);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => 
                           n95436, QN => n116238);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => 
                           n95435, QN => n116266);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => 
                           n95434, QN => n116294);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => 
                           n95433, QN => n116322);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => 
                           n95432, QN => n116350);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => 
                           n95431, QN => n116378);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => 
                           n95430, QN => n116406);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => 
                           n95429, QN => n116434);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n5562, CK => CLK, Q => 
                           n118084, QN => n114583);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n5561, CK => CLK, Q => 
                           n118083, QN => n114584);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n5560, CK => CLK, Q => 
                           n118082, QN => n114585);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n5559, CK => CLK, Q => 
                           n118081, QN => n114586);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n5558, CK => CLK, Q => 
                           n118080, QN => n114587);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n5557, CK => CLK, Q => 
                           n118079, QN => n114588);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n5556, CK => CLK, Q => 
                           n118078, QN => n114589);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n5555, CK => CLK, Q => 
                           n118077, QN => n114590);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n5554, CK => CLK, Q => 
                           n118076, QN => n114591);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n5553, CK => CLK, Q => 
                           n118075, QN => n114592);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n5552, CK => CLK, Q => 
                           n118074, QN => n114593);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n5551, CK => CLK, Q => 
                           n118073, QN => n114594);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n5550, CK => CLK, Q => 
                           n118072, QN => n114595);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n5549, CK => CLK, Q => 
                           n118071, QN => n114596);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n5548, CK => CLK, Q => 
                           n118070, QN => n114597);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n5547, CK => CLK, Q => 
                           n111040, QN => n114598);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n5546, CK => CLK, Q => 
                           n111039, QN => n114599);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n5545, CK => CLK, Q => 
                           n111038, QN => n114600);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n5544, CK => CLK, Q => 
                           n111037, QN => n114601);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n5543, CK => CLK, Q => 
                           n111036, QN => n114602);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n5542, CK => CLK, Q => 
                           n111035, QN => n114603);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n5541, CK => CLK, Q => 
                           n111034, QN => n114604);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n5540, CK => CLK, Q => 
                           n111033, QN => n114605);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n5539, CK => CLK, Q => 
                           n111032, QN => n114606);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n5538, CK => CLK, Q => 
                           n111031, QN => n114607);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n5537, CK => CLK, Q => 
                           n111030, QN => n114608);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n5536, CK => CLK, Q => 
                           n111029, QN => n114609);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n5535, CK => CLK, Q => 
                           n111028, QN => n114610);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n5534, CK => CLK, Q => 
                           n111027, QN => n114611);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n5533, CK => CLK, Q => 
                           n111026, QN => n114612);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n5532, CK => CLK, Q => 
                           n111025, QN => n114613);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n5531, CK => CLK, Q => 
                           n111024, QN => n114614);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n5530, CK => CLK, Q => 
                           n111023, QN => n114615);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n5529, CK => CLK, Q => 
                           n111022, QN => n114616);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n5528, CK => CLK, Q => 
                           n111021, QN => n114617);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n5527, CK => CLK, Q => 
                           n111020, QN => n114618);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n5526, CK => CLK, Q => 
                           n111019, QN => n114619);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n5525, CK => CLK, Q => 
                           n111018, QN => n114620);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n5524, CK => CLK, Q => 
                           n111017, QN => n114621);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n5523, CK => CLK, Q => 
                           n111016, QN => n114622);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n5522, CK => CLK, Q => 
                           n111015, QN => n114623);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n5521, CK => CLK, Q => 
                           n111014, QN => n114624);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n5520, CK => CLK, Q => 
                           n111013, QN => n114625);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n5519, CK => CLK, Q => 
                           n111012, QN => n114626);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n5518, CK => CLK, Q => 
                           n111011, QN => n114627);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n5517, CK => CLK, Q => 
                           n111010, QN => n114628);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n5516, CK => CLK, Q => 
                           n111009, QN => n114629);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n5515, CK => CLK, Q => 
                           n111008, QN => n114630);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n5514, CK => CLK, Q => 
                           n111007, QN => n114631);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => 
                           n111006, QN => n114632);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => 
                           n111005, QN => n114633);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => 
                           n111004, QN => n114634);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => 
                           n111003, QN => n114635);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => 
                           n111002, QN => n114636);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => 
                           n111001, QN => n114637);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => 
                           n111000, QN => n114638);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => 
                           n110999, QN => n114639);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => 
                           n110998, QN => n114640);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => 
                           n110997, QN => n114641);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => 
                           n110996, QN => n114642);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => 
                           n119823, QN => n114515);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n119822, QN => n114516);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => 
                           n119821, QN => n114517);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n119820, QN => n114518);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => 
                           n119819, QN => n114519);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n119818, QN => n114520);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => 
                           n119817, QN => n114521);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n119816, QN => n114522);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => 
                           n119815, QN => n114523);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n119814, QN => n114524);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => 
                           n119813, QN => n114525);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n119812, QN => n114526);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => 
                           n119811, QN => n114527);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n119810, QN => n114528);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => 
                           n119809, QN => n114529);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n119808, QN => n114530);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => 
                           n119807, QN => n114531);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n119806, QN => n114532);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => 
                           n119805, QN => n114533);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => 
                           n119804, QN => n114534);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => 
                           n119803, QN => n114535);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => 
                           n119802, QN => n114536);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => 
                           n119801, QN => n114537);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => 
                           n119800, QN => n114538);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => 
                           n119799, QN => n114539);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => 
                           n119798, QN => n114540);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => 
                           n119797, QN => n114541);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => 
                           n119796, QN => n114542);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => 
                           n119795, QN => n114543);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n119794, QN => n114544);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => 
                           n119793, QN => n114545);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n119792, QN => n114546);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => 
                           n119791, QN => n114547);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n119790, QN => n114548);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => 
                           n119789, QN => n114549);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n119788, QN => n114550);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => 
                           n119787, QN => n114551);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n119786, QN => n114552);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => 
                           n119785, QN => n114553);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n119784, QN => n114554);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => 
                           n119783, QN => n114555);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n119782, QN => n114556);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => 
                           n119781, QN => n114557);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n119780, QN => n114558);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => 
                           n119779, QN => n114559);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n119778, QN => n114560);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => 
                           n119777, QN => n114561);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n119776, QN => n114562);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => 
                           n119775, QN => n114563);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n119774, QN => n114564);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n5640, CK => CLK, Q => 
                           n119773, QN => n114565);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => 
                           n119772, QN => n114566);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => 
                           n119771, QN => n114567);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => 
                           n119770, QN => n114568);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => 
                           n119769, QN => n114569);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => 
                           n119768, QN => n114570);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => 
                           n119767, QN => n114571);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => 
                           n119766, QN => n114572);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => 
                           n119765, QN => n114573);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => 
                           n119764, QN => n114574);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => 
                           n119763, QN => n114449);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n119762, QN => n114450);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => 
                           n119761, QN => n114451);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n119760, QN => n114452);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => 
                           n119759, QN => n114453);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n119758, QN => n114454);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => 
                           n119757, QN => n114455);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n119756, QN => n114456);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => 
                           n119755, QN => n114457);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n119754, QN => n114458);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => 
                           n119753, QN => n114459);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n119752, QN => n114460);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => 
                           n119751, QN => n114461);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n119750, QN => n114462);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => 
                           n119749, QN => n114463);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n119748, QN => n114464);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => 
                           n119747, QN => n114465);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n119746, QN => n114466);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => 
                           n119745, QN => n114467);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n119744, QN => n114468);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => 
                           n119743, QN => n114469);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n119742, QN => n114470);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => 
                           n119741, QN => n114471);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n119740, QN => n114472);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => 
                           n119739, QN => n114473);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n119738, QN => n114474);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => 
                           n119737, QN => n114475);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n119736, QN => n114476);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => 
                           n119735, QN => n114477);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n119734, QN => n114478);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => 
                           n119733, QN => n114479);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n119732, QN => n114480);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => 
                           n119731, QN => n114481);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n119730, QN => n114482);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => 
                           n119729, QN => n114483);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n119728, QN => n114484);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => 
                           n119727, QN => n114485);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n119726, QN => n114486);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => 
                           n119725, QN => n114487);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n119724, QN => n114488);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => 
                           n119723, QN => n114489);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n119722, QN => n114490);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => 
                           n119721, QN => n114491);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n119720, QN => n114492);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => 
                           n119719, QN => n114493);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => 
                           n119718, QN => n114494);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => 
                           n119717, QN => n114495);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => 
                           n119716, QN => n114496);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => 
                           n119715, QN => n114497);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => 
                           n119714, QN => n114498);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => 
                           n119713, QN => n114499);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => 
                           n119712, QN => n114500);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => 
                           n119711, QN => n114501);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => 
                           n119710, QN => n114502);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => 
                           n119709, QN => n114503);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n119708, QN => n114504);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => 
                           n119707, QN => n114505);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n119706, QN => n114506);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => 
                           n119705, QN => n114507);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n119704, QN => n114508);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n119703, QN => n114383);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => 
                           n119702, QN => n114384);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n119701, QN => n114385);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => 
                           n119700, QN => n114386);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n119699, QN => n114387);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => 
                           n119698, QN => n114388);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n119697, QN => n114389);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => 
                           n119696, QN => n114390);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n119695, QN => n114391);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => 
                           n119694, QN => n114392);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n119693, QN => n114393);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => 
                           n119692, QN => n114394);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n119691, QN => n114395);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => 
                           n119690, QN => n114396);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n119689, QN => n114397);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => 
                           n119688, QN => n114398);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n119687, QN => n114399);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => 
                           n119686, QN => n114400);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n119685, QN => n114401);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => 
                           n119684, QN => n114402);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n119683, QN => n114403);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => 
                           n119682, QN => n114404);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n119681, QN => n114405);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => 
                           n119680, QN => n114406);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n119679, QN => n114407);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => 
                           n119678, QN => n114408);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n119677, QN => n114409);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => 
                           n119676, QN => n114410);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n119675, QN => n114411);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => 
                           n119674, QN => n114412);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n119673, QN => n114413);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => 
                           n119672, QN => n114414);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n119671, QN => n114415);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => 
                           n119670, QN => n114416);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n119669, QN => n114417);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => 
                           n119668, QN => n114418);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n119667, QN => n114419);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => 
                           n119666, QN => n114420);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n119665, QN => n114421);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => 
                           n119664, QN => n114422);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n119663, QN => n114423);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => 
                           n119662, QN => n114424);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n119661, QN => n114425);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => 
                           n119660, QN => n114426);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n119659, QN => n114427);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => 
                           n119658, QN => n114428);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n119657, QN => n114429);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => 
                           n119656, QN => n114430);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n119655, QN => n114431);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => 
                           n119654, QN => n114432);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => 
                           n119653, QN => n114433);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => 
                           n119652, QN => n114434);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => 
                           n119651, QN => n114435);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => 
                           n119650, QN => n114436);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => 
                           n119649, QN => n114437);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => 
                           n119648, QN => n114438);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => 
                           n119647, QN => n114439);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => 
                           n119646, QN => n114440);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => 
                           n119645, QN => n114441);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => 
                           n119644, QN => n114442);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n118444, QN => n114311);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n118443, QN => n114312);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n118442, QN => n114313);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n118441, QN => n114314);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n118440, QN => n114315);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n118439, QN => n114316);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n118438, QN => n114317);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n118437, QN => n114318);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n118436, QN => n114319);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n118435, QN => n114320);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n118434, QN => n114321);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n118433, QN => n114322);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n118432, QN => n114323);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n118431, QN => n114324);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n118430, QN => n114325);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n118429, QN => n114326);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n118428, QN => n114327);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n118427, QN => n114328);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n118426, QN => n114329);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n118425, QN => n114330);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n118424, QN => n114331);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n118423, QN => n114332);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n118422, QN => n114333);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n118421, QN => n114334);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n118420, QN => n114335);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n118419, QN => n114336);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n118418, QN => n114337);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n118417, QN => n114338);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n118416, QN => n114339);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n118415, QN => n114340);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n118414, QN => n114341);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n118413, QN => n114342);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n118412, QN => n114343);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n118411, QN => n114344);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n118410, QN => n114345);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n118409, QN => n114346);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n118408, QN => n114347);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n118407, QN => n114348);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n118406, QN => n114349);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n118405, QN => n114350);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n118404, QN => n114351);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n118403, QN => n114352);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n118402, QN => n114353);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n118401, QN => n114354);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n118400, QN => n114355);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n118399, QN => n114356);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n118398, QN => n114357);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n118397, QN => n114358);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n118396, QN => n114359);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n118395, QN => n114360);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n118394, QN => n114361);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => 
                           n118393, QN => n114362);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => 
                           n118392, QN => n114363);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => 
                           n118391, QN => n114364);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => 
                           n118390, QN => n114365);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => 
                           n118389, QN => n114366);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => 
                           n118388, QN => n114367);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => 
                           n118387, QN => n114368);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => 
                           n118386, QN => n114369);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => 
                           n118385, QN => n114370);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n118384, QN => n114240);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n118383, QN => n114241);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n118382, QN => n114242);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n118381, QN => n114243);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n118380, QN => n114244);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n118379, QN => n114245);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n118378, QN => n114246);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n118377, QN => n114247);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n118376, QN => n114248);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n118375, QN => n114249);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n118374, QN => n114250);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n118373, QN => n114251);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n118372, QN => n114252);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n118371, QN => n114253);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n118370, QN => n114254);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n118369, QN => n114255);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n118368, QN => n114256);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n118367, QN => n114257);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n118366, QN => n114258);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n118365, QN => n114259);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n118364, QN => n114260);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n118363, QN => n114261);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n118362, QN => n114262);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n118361, QN => n114263);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n118360, QN => n114264);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n118359, QN => n114265);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n118358, QN => n114266);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n118357, QN => n114267);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n118356, QN => n114268);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n118355, QN => n114269);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n118354, QN => n114270);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n118353, QN => n114271);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n118352, QN => n114272);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n118351, QN => n114273);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n118350, QN => n114274);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n118349, QN => n114275);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n118348, QN => n114276);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n118347, QN => n114277);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n118346, QN => n114278);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n118345, QN => n114279);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n118344, QN => n114280);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n118343, QN => n114281);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n118342, QN => n114282);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n118341, QN => n114283);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n118340, QN => n114284);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n118339, QN => n114285);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n118338, QN => n114286);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n118337, QN => n114287);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n118336, QN => n114288);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n118335, QN => n114289);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n118334, QN => n114290);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n118333, QN => n114291);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n118332, QN => n114292);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n118331, QN => n114293);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n118330, QN => n114294);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n118329, QN => n114295);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n118328, QN => n114296);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n118327, QN => n114297);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n118326, QN => n114298);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n118325, QN => n114299);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n119643, QN => n114151);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n119642, QN => n114152);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n119641, QN => n114153);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n119640, QN => n114154);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n119639, QN => n114155);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n119638, QN => n114156);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n119637, QN => n114157);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n119636, QN => n114158);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n119635, QN => n114159);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n119634, QN => n114160);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n119633, QN => n114161);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n119632, QN => n114162);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n119631, QN => n114163);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n119630, QN => n114164);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n119629, QN => n114165);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n119628, QN => n114166);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n119627, QN => n114167);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n119626, QN => n114168);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n119625, QN => n114169);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n119624, QN => n114170);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n119623, QN => n114171);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n119622, QN => n114172);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n119621, QN => n114173);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n119620, QN => n114174);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n119619, QN => n114175);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n119618, QN => n114176);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n119617, QN => n114177);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n119616, QN => n114178);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n119615, QN => n114179);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n119614, QN => n114180);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n119613, QN => n114181);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n119612, QN => n114182);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n119611, QN => n114183);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n119610, QN => n114184);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n119609, QN => n114185);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n119608, QN => n114186);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n119607, QN => n114187);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n119606, QN => n114188);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n119605, QN => n114189);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n119604, QN => n114190);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n119603, QN => n114191);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n119602, QN => n114192);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n119601, QN => n114193);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n119600, QN => n114194);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n119599, QN => n114195);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n119598, QN => n114196);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n119597, QN => n114197);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n119596, QN => n114198);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n119595, QN => n114199);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n119594, QN => n114200);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n119593, QN => n114201);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n119592, QN => n114202);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n119591, QN => n114203);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n119590, QN => n114204);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n119589, QN => n114205);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n119588, QN => n114206);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n119587, QN => n114207);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n119586, QN => n114208);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n119585, QN => n114209);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n119584, QN => n114210);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => 
                           n117977, QN => n114056);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => 
                           n117976, QN => n114058);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => 
                           n117975, QN => n114059);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => 
                           n117974, QN => n114060);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7482, CK => CLK, Q => 
                           n119583, QN => n113772);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7481, CK => CLK, Q => 
                           n119582, QN => n113774);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7480, CK => CLK, Q => 
                           n119581, QN => n113776);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7479, CK => CLK, Q => 
                           n119580, QN => n113778);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7478, CK => CLK, Q => 
                           n119579, QN => n113780);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7477, CK => CLK, Q => 
                           n119578, QN => n113782);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7476, CK => CLK, Q => 
                           n119577, QN => n113784);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7475, CK => CLK, Q => 
                           n119576, QN => n113786);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7474, CK => CLK, Q => 
                           n119575, QN => n113788);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7473, CK => CLK, Q => 
                           n119574, QN => n113790);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7472, CK => CLK, Q => 
                           n119573, QN => n113792);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7471, CK => CLK, Q => 
                           n119572, QN => n113794);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7470, CK => CLK, Q => 
                           n119571, QN => n113796);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7469, CK => CLK, Q => 
                           n119570, QN => n113798);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7468, CK => CLK, Q => 
                           n119569, QN => n113800);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7467, CK => CLK, Q => 
                           n119568, QN => n113802);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7466, CK => CLK, Q => 
                           n119567, QN => n113804);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7465, CK => CLK, Q => 
                           n119566, QN => n113806);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7464, CK => CLK, Q => 
                           n119565, QN => n113808);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7463, CK => CLK, Q => 
                           n119564, QN => n113810);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7462, CK => CLK, Q => 
                           n119563, QN => n113812);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7461, CK => CLK, Q => 
                           n119562, QN => n113814);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7460, CK => CLK, Q => 
                           n119561, QN => n113816);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7459, CK => CLK, Q => 
                           n119560, QN => n113818);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7458, CK => CLK, Q => 
                           n119559, QN => n113820);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7457, CK => CLK, Q => 
                           n119558, QN => n113822);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7456, CK => CLK, Q => 
                           n119557, QN => n113824);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7455, CK => CLK, Q => 
                           n119556, QN => n113826);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7454, CK => CLK, Q => 
                           n119555, QN => n113828);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7453, CK => CLK, Q => 
                           n119554, QN => n113830);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7452, CK => CLK, Q => 
                           n119553, QN => n113832);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7451, CK => CLK, Q => 
                           n119552, QN => n113834);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7450, CK => CLK, Q => 
                           n119551, QN => n113836);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7449, CK => CLK, Q => 
                           n119550, QN => n113838);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7448, CK => CLK, Q => 
                           n119549, QN => n113840);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7447, CK => CLK, Q => 
                           n119548, QN => n113842);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7446, CK => CLK, Q => 
                           n119547, QN => n113844);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7445, CK => CLK, Q => 
                           n119546, QN => n113846);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7444, CK => CLK, Q => 
                           n119545, QN => n113848);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7443, CK => CLK, Q => 
                           n119544, QN => n113850);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7442, CK => CLK, Q => 
                           n119543, QN => n113852);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7441, CK => CLK, Q => 
                           n119542, QN => n113854);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7440, CK => CLK, Q => 
                           n119541, QN => n113856);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7439, CK => CLK, Q => 
                           n119540, QN => n113858);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7438, CK => CLK, Q => 
                           n119539, QN => n113860);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7437, CK => CLK, Q => 
                           n119538, QN => n113862);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7436, CK => CLK, Q => 
                           n119537, QN => n113864);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7435, CK => CLK, Q => 
                           n119536, QN => n113866);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7434, CK => CLK, Q => 
                           n119535, QN => n113868);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7433, CK => CLK, Q => 
                           n119534, QN => n113870);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7432, CK => CLK, Q => 
                           n119533, QN => n113872);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7431, CK => CLK, Q => 
                           n119532, QN => n113874);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7430, CK => CLK, Q => 
                           n119531, QN => n113876);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7429, CK => CLK, Q => 
                           n119530, QN => n113878);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7428, CK => CLK, Q => 
                           n119529, QN => n113880);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7427, CK => CLK, Q => 
                           n119528, QN => n113882);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7426, CK => CLK, Q => 
                           n119527, QN => n113884);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7425, CK => CLK, Q => 
                           n119526, QN => n113886);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7424, CK => CLK, Q => 
                           n119525, QN => n113888);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7423, CK => CLK, Q => 
                           n119524, QN => n113890);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n119523, QN => n113992);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n119522, QN => n113993);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n119521, QN => n113994);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n119520, QN => n113995);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n119519, QN => n113996);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n119518, QN => n113997);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n119517, QN => n113998);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n119516, QN => n113999);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n119515, QN => n114000);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n119514, QN => n114001);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n119513, QN => n114002);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n119512, QN => n114003);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n119511, QN => n114004);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n119510, QN => n114005);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n119509, QN => n114006);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n119508, QN => n114007);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n119507, QN => n114008);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n119506, QN => n114009);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n119505, QN => n114010);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n119504, QN => n114011);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n119503, QN => n114012);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n119502, QN => n114013);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n119501, QN => n114014);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n119500, QN => n114015);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n119499, QN => n114016);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n119498, QN => n114017);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => 
                           n119497, QN => n114018);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => 
                           n119496, QN => n114019);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => 
                           n119495, QN => n114020);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n119494, QN => n114021);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n119493, QN => n114022);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n119492, QN => n114023);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n119491, QN => n114024);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n119490, QN => n114025);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n119489, QN => n114026);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n119488, QN => n114027);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n119487, QN => n114028);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n119486, QN => n114029);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n119485, QN => n114030);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n119484, QN => n114031);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n119483, QN => n114032);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n119482, QN => n114033);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n119481, QN => n114034);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n119480, QN => n114035);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n119479, QN => n114036);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n119478, QN => n114037);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n119477, QN => n114038);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n119476, QN => n114039);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n119475, QN => n114040);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n119474, QN => n114041);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => 
                           n119473, QN => n114042);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => 
                           n119472, QN => n114043);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => 
                           n119471, QN => n114044);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => 
                           n119470, QN => n114045);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => 
                           n119469, QN => n114046);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => 
                           n119468, QN => n114047);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => 
                           n119467, QN => n114048);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => 
                           n119466, QN => n114049);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => 
                           n119465, QN => n114050);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => 
                           n119464, QN => n114051);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => 
                           n119463, QN => n113920);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => 
                           n119462, QN => n113921);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => 
                           n119461, QN => n113922);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => 
                           n119460, QN => n113923);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => 
                           n119459, QN => n113924);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => 
                           n119458, QN => n113925);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => 
                           n119457, QN => n113926);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => 
                           n119456, QN => n113927);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => 
                           n119455, QN => n113928);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => 
                           n119454, QN => n113929);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => 
                           n119453, QN => n113930);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => 
                           n119452, QN => n113931);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => 
                           n119451, QN => n113932);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => 
                           n119450, QN => n113933);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => 
                           n119449, QN => n113934);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => 
                           n119448, QN => n113935);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => 
                           n119447, QN => n113936);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => 
                           n119446, QN => n113937);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => 
                           n119445, QN => n113938);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => 
                           n119444, QN => n113939);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => 
                           n119443, QN => n113940);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => 
                           n119442, QN => n113941);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => 
                           n119441, QN => n113942);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => 
                           n119440, QN => n113943);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => 
                           n119439, QN => n113944);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n7137, CK => CLK, Q => 
                           n119438, QN => n113945);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n7136, CK => CLK, Q => 
                           n119437, QN => n113946);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n7135, CK => CLK, Q => 
                           n119436, QN => n113947);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7134, CK => CLK, Q => 
                           n119435, QN => n113948);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7133, CK => CLK, Q => 
                           n119434, QN => n113949);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7132, CK => CLK, Q => 
                           n119433, QN => n113950);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7131, CK => CLK, Q => 
                           n119432, QN => n113951);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7130, CK => CLK, Q => 
                           n119431, QN => n113952);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7129, CK => CLK, Q => 
                           n119430, QN => n113953);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7128, CK => CLK, Q => 
                           n119429, QN => n113954);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7127, CK => CLK, Q => 
                           n119428, QN => n113955);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7126, CK => CLK, Q => 
                           n119427, QN => n113956);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7125, CK => CLK, Q => 
                           n119426, QN => n113957);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7124, CK => CLK, Q => 
                           n119425, QN => n113958);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7123, CK => CLK, Q => 
                           n119424, QN => n113959);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7122, CK => CLK, Q => 
                           n119423, QN => n113960);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7121, CK => CLK, Q => 
                           n119422, QN => n113961);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7120, CK => CLK, Q => 
                           n119421, QN => n113962);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7119, CK => CLK, Q => 
                           n119420, QN => n113963);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           n119419, QN => n113964);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7117, CK => CLK, Q => 
                           n119418, QN => n113965);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7116, CK => CLK, Q => 
                           n119417, QN => n113966);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7115, CK => CLK, Q => 
                           n119416, QN => n113967);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7114, CK => CLK, Q => 
                           n119415, QN => n113968);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7113, CK => CLK, Q => 
                           n119414, QN => n113969);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7112, CK => CLK, Q => 
                           n119413, QN => n113970);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7111, CK => CLK, Q => 
                           n119412, QN => n113971);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7110, CK => CLK, Q => 
                           n119411, QN => n113972);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7109, CK => CLK, Q => 
                           n119410, QN => n113973);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7108, CK => CLK, Q => 
                           n119409, QN => n113974);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => 
                           n119408, QN => n113975);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => 
                           n119407, QN => n113976);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => 
                           n119406, QN => n113977);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => 
                           n119405, QN => n113978);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => 
                           n119404, QN => n113979);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => 
                           n118264, QN => n114061);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => 
                           n118263, QN => n114062);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => 
                           n118262, QN => n114063);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => 
                           n118261, QN => n114064);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => 
                           n118260, QN => n114065);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => 
                           n118259, QN => n114066);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => 
                           n118258, QN => n114067);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => 
                           n118257, QN => n114068);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => 
                           n118256, QN => n114069);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => 
                           n118255, QN => n114070);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => 
                           n118254, QN => n114071);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => 
                           n118253, QN => n114072);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => 
                           n118252, QN => n114073);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => 
                           n118251, QN => n114074);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => 
                           n118250, QN => n114075);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => 
                           n118249, QN => n114076);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => 
                           n118248, QN => n114077);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => 
                           n118247, QN => n114078);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => 
                           n118246, QN => n114079);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => 
                           n118245, QN => n114080);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => 
                           n118244, QN => n114081);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => 
                           n118243, QN => n114082);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => 
                           n118242, QN => n114083);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => 
                           n118241, QN => n114084);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => 
                           n118240, QN => n114085);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => 
                           n118239, QN => n114086);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => 
                           n118238, QN => n114087);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => 
                           n118237, QN => n114088);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => 
                           n118236, QN => n114089);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => 
                           n118235, QN => n114090);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => 
                           n118234, QN => n114091);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => 
                           n118233, QN => n114092);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => 
                           n118232, QN => n114093);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => 
                           n118231, QN => n114094);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => 
                           n118230, QN => n114095);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => 
                           n118229, QN => n114096);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => 
                           n118228, QN => n114097);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => 
                           n118227, QN => n114098);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => 
                           n118226, QN => n114099);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => 
                           n118225, QN => n114100);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => 
                           n118224, QN => n114101);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => 
                           n118223, QN => n114102);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => 
                           n118222, QN => n114103);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => 
                           n118221, QN => n114104);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => 
                           n118220, QN => n114105);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => 
                           n118219, QN => n114106);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => 
                           n118218, QN => n114107);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => 
                           n118217, QN => n114108);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => 
                           n118216, QN => n114109);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => 
                           n118215, QN => n114110);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => 
                           n118214, QN => n114111);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => 
                           n118213, QN => n114112);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => 
                           n118212, QN => n114113);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => 
                           n118211, QN => n114114);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => 
                           n118210, QN => n114115);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => 
                           n118209, QN => n114116);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => 
                           n118208, QN => n114117);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => 
                           n118207, QN => n114118);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => 
                           n118206, QN => n114119);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => 
                           n118205, QN => n114120);
   OUT1_reg_63_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => OUT1_63_port
                           , QN => n119403);
   OUT1_reg_62_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => OUT1_62_port
                           , QN => n119402);
   OUT1_reg_61_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => OUT1_61_port
                           , QN => n119401);
   OUT1_reg_60_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => OUT1_60_port
                           , QN => n119400);
   OUT2_reg_63_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => OUT2_63_port
                           , QN => n119399);
   OUT2_reg_62_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => OUT2_62_port
                           , QN => n119398);
   OUT2_reg_61_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => OUT2_61_port
                           , QN => n119397);
   OUT2_reg_60_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => OUT2_60_port
                           , QN => n119396);
   OUT2_reg_59_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => OUT2_59_port
                           , QN => n119395);
   OUT2_reg_58_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => OUT2_58_port
                           , QN => n119394);
   OUT2_reg_57_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => OUT2_57_port
                           , QN => n119393);
   OUT2_reg_56_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => OUT2_56_port
                           , QN => n119392);
   OUT2_reg_55_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => OUT2_55_port
                           , QN => n119391);
   OUT2_reg_54_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => OUT2_54_port
                           , QN => n119390);
   OUT2_reg_53_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => OUT2_53_port
                           , QN => n119389);
   OUT2_reg_52_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => OUT2_52_port
                           , QN => n119388);
   OUT2_reg_51_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => OUT2_51_port
                           , QN => n119387);
   OUT2_reg_50_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => OUT2_50_port
                           , QN => n119386);
   OUT2_reg_49_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => OUT2_49_port
                           , QN => n119385);
   OUT2_reg_48_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => OUT2_48_port
                           , QN => n119384);
   OUT2_reg_47_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => OUT2_47_port
                           , QN => n119383);
   OUT2_reg_46_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => OUT2_46_port
                           , QN => n119382);
   OUT2_reg_45_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => OUT2_45_port
                           , QN => n119381);
   OUT2_reg_44_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => OUT2_44_port
                           , QN => n119380);
   OUT2_reg_43_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => OUT2_43_port
                           , QN => n119379);
   OUT2_reg_42_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => OUT2_42_port
                           , QN => n119378);
   OUT2_reg_41_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => OUT2_41_port
                           , QN => n119377);
   OUT2_reg_40_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => OUT2_40_port
                           , QN => n119376);
   OUT2_reg_39_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => OUT2_39_port
                           , QN => n119375);
   OUT2_reg_38_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => OUT2_38_port
                           , QN => n119374);
   OUT2_reg_37_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => OUT2_37_port
                           , QN => n119373);
   OUT2_reg_36_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => OUT2_36_port
                           , QN => n119372);
   OUT2_reg_35_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => OUT2_35_port
                           , QN => n119371);
   OUT2_reg_34_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => OUT2_34_port
                           , QN => n119370);
   OUT2_reg_33_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => OUT2_33_port
                           , QN => n119369);
   OUT2_reg_32_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => OUT2_32_port
                           , QN => n119368);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => OUT2_31_port
                           , QN => n119367);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5341, CK => CLK, Q => OUT2_30_port
                           , QN => n119366);
   U83326 : NOR3_X1 port map( A1 => n120018, A2 => ADD_RD2(2), A3 => n117973, 
                           ZN => n117945);
   U83327 : NOR3_X1 port map( A1 => n120018, A2 => ADD_RD2(1), A3 => n117971, 
                           ZN => n117953);
   U83328 : NOR3_X1 port map( A1 => n117971, A2 => n120018, A3 => n117973, ZN 
                           => n117948);
   U83329 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n120018
                           , ZN => n117954);
   U83330 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n120216
                           , ZN => n116445);
   U83331 : BUF_X1 port map( A => n120827, Z => n120829);
   U83332 : BUF_X1 port map( A => n120828, Z => n120833);
   U83333 : BUF_X1 port map( A => n120828, Z => n120832);
   U83334 : BUF_X1 port map( A => n120827, Z => n120831);
   U83335 : BUF_X1 port map( A => n120827, Z => n120830);
   U83336 : BUF_X1 port map( A => n116528, Z => n119863);
   U83337 : BUF_X1 port map( A => n116528, Z => n119864);
   U83338 : BUF_X1 port map( A => n116528, Z => n119865);
   U83339 : BUF_X1 port map( A => n116528, Z => n119866);
   U83340 : BUF_X1 port map( A => n116528, Z => n119862);
   U83341 : BUF_X1 port map( A => n113767, Z => n120822);
   U83342 : BUF_X1 port map( A => n113767, Z => n120823);
   U83343 : BUF_X1 port map( A => n113767, Z => n120824);
   U83344 : BUF_X1 port map( A => n113767, Z => n120825);
   U83345 : BUF_X1 port map( A => n120543, Z => n120545);
   U83346 : BUF_X1 port map( A => n120246, Z => n120248);
   U83347 : BUF_X1 port map( A => n120259, Z => n120261);
   U83348 : BUF_X1 port map( A => n120518, Z => n120520);
   U83349 : BUF_X1 port map( A => n120568, Z => n120570);
   U83350 : BUF_X1 port map( A => n120372, Z => n120374);
   U83351 : BUF_X1 port map( A => n120335, Z => n120337);
   U83352 : BUF_X1 port map( A => n120284, Z => n120286);
   U83353 : BUF_X1 port map( A => n120409, Z => n120411);
   U83354 : BUF_X1 port map( A => n120310, Z => n120312);
   U83355 : BUF_X1 port map( A => n120297, Z => n120299);
   U83356 : BUF_X1 port map( A => n120544, Z => n120549);
   U83357 : BUF_X1 port map( A => n120544, Z => n120548);
   U83358 : BUF_X1 port map( A => n120543, Z => n120547);
   U83359 : BUF_X1 port map( A => n120543, Z => n120546);
   U83360 : BUF_X1 port map( A => n120246, Z => n120249);
   U83361 : BUF_X1 port map( A => n120246, Z => n120250);
   U83362 : BUF_X1 port map( A => n120247, Z => n120251);
   U83363 : BUF_X1 port map( A => n120259, Z => n120262);
   U83364 : BUF_X1 port map( A => n120259, Z => n120263);
   U83365 : BUF_X1 port map( A => n120247, Z => n120252);
   U83366 : BUF_X1 port map( A => n120518, Z => n120521);
   U83367 : BUF_X1 port map( A => n120518, Z => n120522);
   U83368 : BUF_X1 port map( A => n120519, Z => n120523);
   U83369 : BUF_X1 port map( A => n120568, Z => n120571);
   U83370 : BUF_X1 port map( A => n120568, Z => n120572);
   U83371 : BUF_X1 port map( A => n120569, Z => n120573);
   U83372 : BUF_X1 port map( A => n120519, Z => n120524);
   U83373 : BUF_X1 port map( A => n120372, Z => n120375);
   U83374 : BUF_X1 port map( A => n120372, Z => n120376);
   U83375 : BUF_X1 port map( A => n120373, Z => n120377);
   U83376 : BUF_X1 port map( A => n120335, Z => n120338);
   U83377 : BUF_X1 port map( A => n120335, Z => n120339);
   U83378 : BUF_X1 port map( A => n120336, Z => n120340);
   U83379 : BUF_X1 port map( A => n120284, Z => n120287);
   U83380 : BUF_X1 port map( A => n120284, Z => n120288);
   U83381 : BUF_X1 port map( A => n120285, Z => n120289);
   U83382 : BUF_X1 port map( A => n120260, Z => n120264);
   U83383 : BUF_X1 port map( A => n120409, Z => n120412);
   U83384 : BUF_X1 port map( A => n120409, Z => n120413);
   U83385 : BUF_X1 port map( A => n120410, Z => n120414);
   U83386 : BUF_X1 port map( A => n120310, Z => n120313);
   U83387 : BUF_X1 port map( A => n120310, Z => n120314);
   U83388 : BUF_X1 port map( A => n120311, Z => n120315);
   U83389 : BUF_X1 port map( A => n120569, Z => n120574);
   U83390 : BUF_X1 port map( A => n120373, Z => n120378);
   U83391 : BUF_X1 port map( A => n120336, Z => n120341);
   U83392 : BUF_X1 port map( A => n120285, Z => n120290);
   U83393 : BUF_X1 port map( A => n120260, Z => n120265);
   U83394 : BUF_X1 port map( A => n120297, Z => n120300);
   U83395 : BUF_X1 port map( A => n120297, Z => n120301);
   U83396 : BUF_X1 port map( A => n120298, Z => n120302);
   U83397 : BUF_X1 port map( A => n120410, Z => n120415);
   U83398 : BUF_X1 port map( A => n120298, Z => n120303);
   U83399 : BUF_X1 port map( A => n120311, Z => n120316);
   U83400 : BUF_X1 port map( A => n114139, Z => n120434);
   U83401 : BUF_X1 port map( A => n114139, Z => n120435);
   U83402 : BUF_X1 port map( A => n114139, Z => n120436);
   U83403 : BUF_X1 port map( A => n114139, Z => n120437);
   U83404 : BUF_X1 port map( A => n114139, Z => n120438);
   U83405 : BUF_X1 port map( A => n114645, Z => n120240);
   U83406 : BUF_X1 port map( A => n114645, Z => n120241);
   U83407 : BUF_X1 port map( A => n114645, Z => n120242);
   U83408 : BUF_X1 port map( A => n114645, Z => n120243);
   U83409 : BUF_X1 port map( A => n114645, Z => n120244);
   U83410 : BUF_X1 port map( A => n113897, Z => n120611);
   U83411 : BUF_X1 port map( A => n113897, Z => n120612);
   U83412 : BUF_X1 port map( A => n113897, Z => n120613);
   U83413 : BUF_X1 port map( A => n113897, Z => n120614);
   U83414 : BUF_X1 port map( A => n113897, Z => n120615);
   U83415 : BUF_X1 port map( A => n113904, Z => n120599);
   U83416 : BUF_X1 port map( A => n113904, Z => n120600);
   U83417 : BUF_X1 port map( A => n113904, Z => n120601);
   U83418 : BUF_X1 port map( A => n113904, Z => n120602);
   U83419 : BUF_X1 port map( A => n113904, Z => n120603);
   U83420 : BUF_X1 port map( A => n113991, Z => n120537);
   U83421 : BUF_X1 port map( A => n113991, Z => n120538);
   U83422 : BUF_X1 port map( A => n113991, Z => n120539);
   U83423 : BUF_X1 port map( A => n113991, Z => n120540);
   U83424 : BUF_X1 port map( A => n113991, Z => n120541);
   U83425 : BUF_X1 port map( A => n114214, Z => n120379);
   U83426 : BUF_X1 port map( A => n114579, Z => n120253);
   U83427 : BUF_X1 port map( A => n114579, Z => n120254);
   U83428 : BUF_X1 port map( A => n114579, Z => n120255);
   U83429 : BUF_X1 port map( A => n114133, Z => n120464);
   U83430 : BUF_X1 port map( A => n114133, Z => n120465);
   U83431 : BUF_X1 port map( A => n114133, Z => n120466);
   U83432 : BUF_X1 port map( A => n114133, Z => n120467);
   U83433 : BUF_X1 port map( A => n114133, Z => n120468);
   U83434 : BUF_X1 port map( A => n114137, Z => n120440);
   U83435 : BUF_X1 port map( A => n114137, Z => n120441);
   U83436 : BUF_X1 port map( A => n114137, Z => n120442);
   U83437 : BUF_X1 port map( A => n114137, Z => n120443);
   U83438 : BUF_X1 port map( A => n114137, Z => n120444);
   U83439 : BUF_X1 port map( A => n114057, Z => n120512);
   U83440 : BUF_X1 port map( A => n114057, Z => n120513);
   U83441 : BUF_X1 port map( A => n114057, Z => n120514);
   U83442 : BUF_X1 port map( A => n114057, Z => n120515);
   U83443 : BUF_X1 port map( A => n114057, Z => n120516);
   U83444 : BUF_X1 port map( A => n114129, Z => n120488);
   U83445 : BUF_X1 port map( A => n114129, Z => n120489);
   U83446 : BUF_X1 port map( A => n114129, Z => n120490);
   U83447 : BUF_X1 port map( A => n114129, Z => n120491);
   U83448 : BUF_X1 port map( A => n114129, Z => n120492);
   U83449 : BUF_X1 port map( A => n114131, Z => n120476);
   U83450 : BUF_X1 port map( A => n114131, Z => n120477);
   U83451 : BUF_X1 port map( A => n114131, Z => n120478);
   U83452 : BUF_X1 port map( A => n114131, Z => n120479);
   U83453 : BUF_X1 port map( A => n114131, Z => n120480);
   U83454 : BUF_X1 port map( A => n114135, Z => n120452);
   U83455 : BUF_X1 port map( A => n114135, Z => n120453);
   U83456 : BUF_X1 port map( A => n114135, Z => n120454);
   U83457 : BUF_X1 port map( A => n114135, Z => n120455);
   U83458 : BUF_X1 port map( A => n114135, Z => n120456);
   U83459 : BUF_X1 port map( A => n113912, Z => n120575);
   U83460 : BUF_X1 port map( A => n113912, Z => n120576);
   U83461 : BUF_X1 port map( A => n113912, Z => n120577);
   U83462 : BUF_X1 port map( A => n113912, Z => n120578);
   U83463 : BUF_X1 port map( A => n113912, Z => n120579);
   U83464 : BUF_X1 port map( A => n114124, Z => n120500);
   U83465 : BUF_X1 port map( A => n114124, Z => n120501);
   U83466 : BUF_X1 port map( A => n114124, Z => n120502);
   U83467 : BUF_X1 port map( A => n114124, Z => n120503);
   U83468 : BUF_X1 port map( A => n114124, Z => n120504);
   U83469 : BUF_X1 port map( A => n113982, Z => n120550);
   U83470 : BUF_X1 port map( A => n113982, Z => n120551);
   U83471 : BUF_X1 port map( A => n113982, Z => n120552);
   U83472 : BUF_X1 port map( A => n113982, Z => n120553);
   U83473 : BUF_X1 port map( A => n113982, Z => n120554);
   U83474 : BUF_X1 port map( A => n113910, Z => n120587);
   U83475 : BUF_X1 port map( A => n113910, Z => n120588);
   U83476 : BUF_X1 port map( A => n113910, Z => n120589);
   U83477 : BUF_X1 port map( A => n113910, Z => n120590);
   U83478 : BUF_X1 port map( A => n113910, Z => n120591);
   U83479 : BUF_X1 port map( A => n113916, Z => n120562);
   U83480 : BUF_X1 port map( A => n113916, Z => n120563);
   U83481 : BUF_X1 port map( A => n113916, Z => n120564);
   U83482 : BUF_X1 port map( A => n113916, Z => n120565);
   U83483 : BUF_X1 port map( A => n113916, Z => n120566);
   U83484 : BUF_X1 port map( A => n114301, Z => n120354);
   U83485 : BUF_X1 port map( A => n114301, Z => n120355);
   U83486 : BUF_X1 port map( A => n114301, Z => n120356);
   U83487 : BUF_X1 port map( A => n114301, Z => n120357);
   U83488 : BUF_X1 port map( A => n114301, Z => n120358);
   U83489 : BUF_X1 port map( A => n114236, Z => n120366);
   U83490 : BUF_X1 port map( A => n114236, Z => n120367);
   U83491 : BUF_X1 port map( A => n114236, Z => n120368);
   U83492 : BUF_X1 port map( A => n114236, Z => n120369);
   U83493 : BUF_X1 port map( A => n114236, Z => n120370);
   U83494 : BUF_X1 port map( A => n114307, Z => n120329);
   U83495 : BUF_X1 port map( A => n114307, Z => n120330);
   U83496 : BUF_X1 port map( A => n114307, Z => n120331);
   U83497 : BUF_X1 port map( A => n114307, Z => n120332);
   U83498 : BUF_X1 port map( A => n114307, Z => n120333);
   U83499 : BUF_X1 port map( A => n114212, Z => n120391);
   U83500 : BUF_X1 port map( A => n114212, Z => n120392);
   U83501 : BUF_X1 port map( A => n114212, Z => n120393);
   U83502 : BUF_X1 port map( A => n114212, Z => n120394);
   U83503 : BUF_X1 port map( A => n114212, Z => n120395);
   U83504 : BUF_X1 port map( A => n114373, Z => n120317);
   U83505 : BUF_X1 port map( A => n114373, Z => n120318);
   U83506 : BUF_X1 port map( A => n114373, Z => n120319);
   U83507 : BUF_X1 port map( A => n114373, Z => n120320);
   U83508 : BUF_X1 port map( A => n114373, Z => n120321);
   U83509 : BUF_X1 port map( A => n114511, Z => n120278);
   U83510 : BUF_X1 port map( A => n114511, Z => n120279);
   U83511 : BUF_X1 port map( A => n114511, Z => n120280);
   U83512 : BUF_X1 port map( A => n114511, Z => n120281);
   U83513 : BUF_X1 port map( A => n114511, Z => n120282);
   U83514 : BUF_X1 port map( A => n114576, Z => n120266);
   U83515 : BUF_X1 port map( A => n114576, Z => n120267);
   U83516 : BUF_X1 port map( A => n114576, Z => n120268);
   U83517 : BUF_X1 port map( A => n114576, Z => n120269);
   U83518 : BUF_X1 port map( A => n114576, Z => n120270);
   U83519 : BUF_X1 port map( A => n114579, Z => n120256);
   U83520 : BUF_X1 port map( A => n114579, Z => n120257);
   U83521 : BUF_X1 port map( A => n114147, Z => n120403);
   U83522 : BUF_X1 port map( A => n114147, Z => n120404);
   U83523 : BUF_X1 port map( A => n114147, Z => n120405);
   U83524 : BUF_X1 port map( A => n114147, Z => n120406);
   U83525 : BUF_X1 port map( A => n114147, Z => n120407);
   U83526 : BUF_X1 port map( A => n114379, Z => n120304);
   U83527 : BUF_X1 port map( A => n114379, Z => n120305);
   U83528 : BUF_X1 port map( A => n114379, Z => n120306);
   U83529 : BUF_X1 port map( A => n114379, Z => n120307);
   U83530 : BUF_X1 port map( A => n114214, Z => n120380);
   U83531 : BUF_X1 port map( A => n114214, Z => n120381);
   U83532 : BUF_X1 port map( A => n114214, Z => n120382);
   U83533 : BUF_X1 port map( A => n114214, Z => n120383);
   U83534 : BUF_X1 port map( A => n114140, Z => n120428);
   U83535 : BUF_X1 port map( A => n114140, Z => n120429);
   U83536 : BUF_X1 port map( A => n114140, Z => n120430);
   U83537 : BUF_X1 port map( A => n114140, Z => n120431);
   U83538 : BUF_X1 port map( A => n114140, Z => n120432);
   U83539 : BUF_X1 port map( A => n114143, Z => n120416);
   U83540 : BUF_X1 port map( A => n114143, Z => n120417);
   U83541 : BUF_X1 port map( A => n114143, Z => n120418);
   U83542 : BUF_X1 port map( A => n114143, Z => n120419);
   U83543 : BUF_X1 port map( A => n114143, Z => n120420);
   U83544 : BUF_X1 port map( A => n114304, Z => n120342);
   U83545 : BUF_X1 port map( A => n114304, Z => n120343);
   U83546 : BUF_X1 port map( A => n114304, Z => n120344);
   U83547 : BUF_X1 port map( A => n114304, Z => n120345);
   U83548 : BUF_X1 port map( A => n114304, Z => n120346);
   U83549 : BUF_X1 port map( A => n114445, Z => n120291);
   U83550 : BUF_X1 port map( A => n114445, Z => n120292);
   U83551 : BUF_X1 port map( A => n114445, Z => n120293);
   U83552 : BUF_X1 port map( A => n114445, Z => n120294);
   U83553 : BUF_X1 port map( A => n114445, Z => n120295);
   U83554 : BUF_X1 port map( A => n114053, Z => n120525);
   U83555 : BUF_X1 port map( A => n114053, Z => n120526);
   U83556 : BUF_X1 port map( A => n114053, Z => n120527);
   U83557 : BUF_X1 port map( A => n114053, Z => n120528);
   U83558 : BUF_X1 port map( A => n114053, Z => n120529);
   U83559 : BUF_X1 port map( A => n114379, Z => n120308);
   U83560 : BUF_X1 port map( A => n114689, Z => n120100);
   U83561 : BUF_X1 port map( A => n114689, Z => n120096);
   U83562 : BUF_X1 port map( A => n114689, Z => n120097);
   U83563 : BUF_X1 port map( A => n114689, Z => n120098);
   U83564 : BUF_X1 port map( A => n114689, Z => n120099);
   U83565 : BUF_X1 port map( A => n113767, Z => n120821);
   U83566 : BUF_X1 port map( A => n113766, Z => n120827);
   U83567 : BUF_X1 port map( A => n113766, Z => n120828);
   U83568 : OAI21_X1 port map( B1 => n113894, B2 => n114141, A => n120624, ZN 
                           => n114139);
   U83569 : NAND2_X1 port map( A1 => n116447, A2 => n116463, ZN => n114689);
   U83570 : BUF_X1 port map( A => n116522, Z => n119887);
   U83571 : BUF_X1 port map( A => n116522, Z => n119888);
   U83572 : BUF_X1 port map( A => n116522, Z => n119889);
   U83573 : BUF_X1 port map( A => n116522, Z => n119890);
   U83574 : BUF_X1 port map( A => n114691, Z => n120088);
   U83575 : BUF_X1 port map( A => n114698, Z => n120064);
   U83576 : BUF_X1 port map( A => n116522, Z => n119886);
   U83577 : BUF_X1 port map( A => n114691, Z => n120084);
   U83578 : BUF_X1 port map( A => n114698, Z => n120060);
   U83579 : BUF_X1 port map( A => n114691, Z => n120085);
   U83580 : BUF_X1 port map( A => n114698, Z => n120061);
   U83581 : BUF_X1 port map( A => n114691, Z => n120086);
   U83582 : BUF_X1 port map( A => n114698, Z => n120062);
   U83583 : BUF_X1 port map( A => n114691, Z => n120087);
   U83584 : BUF_X1 port map( A => n114698, Z => n120063);
   U83585 : BUF_X1 port map( A => n116490, Z => n120025);
   U83586 : BUF_X1 port map( A => n116490, Z => n120026);
   U83587 : BUF_X1 port map( A => n116490, Z => n120027);
   U83588 : BUF_X1 port map( A => n116490, Z => n120028);
   U83589 : BUF_X1 port map( A => n114662, Z => n120202);
   U83590 : BUF_X1 port map( A => n116490, Z => n120024);
   U83591 : BUF_X1 port map( A => n114662, Z => n120198);
   U83592 : BUF_X1 port map( A => n114662, Z => n120199);
   U83593 : BUF_X1 port map( A => n114662, Z => n120200);
   U83594 : BUF_X1 port map( A => n114662, Z => n120201);
   U83595 : BUF_X1 port map( A => n114657, Z => n120226);
   U83596 : BUF_X1 port map( A => n114657, Z => n120222);
   U83597 : BUF_X1 port map( A => n114657, Z => n120223);
   U83598 : BUF_X1 port map( A => n114657, Z => n120224);
   U83599 : BUF_X1 port map( A => n114657, Z => n120225);
   U83600 : BUF_X1 port map( A => n116495, Z => n120001);
   U83601 : BUF_X1 port map( A => n116502, Z => n119977);
   U83602 : BUF_X1 port map( A => n116507, Z => n119953);
   U83603 : BUF_X1 port map( A => n116495, Z => n120002);
   U83604 : BUF_X1 port map( A => n116502, Z => n119978);
   U83605 : BUF_X1 port map( A => n116507, Z => n119954);
   U83606 : BUF_X1 port map( A => n116495, Z => n120003);
   U83607 : BUF_X1 port map( A => n116502, Z => n119979);
   U83608 : BUF_X1 port map( A => n116507, Z => n119955);
   U83609 : BUF_X1 port map( A => n116495, Z => n120004);
   U83610 : BUF_X1 port map( A => n116502, Z => n119980);
   U83611 : BUF_X1 port map( A => n116507, Z => n119956);
   U83612 : BUF_X1 port map( A => n114669, Z => n120178);
   U83613 : BUF_X1 port map( A => n114675, Z => n120154);
   U83614 : BUF_X1 port map( A => n116495, Z => n120000);
   U83615 : BUF_X1 port map( A => n116502, Z => n119976);
   U83616 : BUF_X1 port map( A => n116507, Z => n119952);
   U83617 : BUF_X1 port map( A => n114669, Z => n120174);
   U83618 : BUF_X1 port map( A => n114675, Z => n120150);
   U83619 : BUF_X1 port map( A => n114669, Z => n120175);
   U83620 : BUF_X1 port map( A => n114675, Z => n120151);
   U83621 : BUF_X1 port map( A => n114669, Z => n120176);
   U83622 : BUF_X1 port map( A => n114675, Z => n120152);
   U83623 : BUF_X1 port map( A => n114669, Z => n120177);
   U83624 : BUF_X1 port map( A => n114675, Z => n120153);
   U83625 : BUF_X1 port map( A => n116523, Z => n119881);
   U83626 : BUF_X1 port map( A => n116523, Z => n119882);
   U83627 : BUF_X1 port map( A => n116523, Z => n119883);
   U83628 : BUF_X1 port map( A => n116523, Z => n119884);
   U83629 : BUF_X1 port map( A => n116523, Z => n119880);
   U83630 : BUF_X1 port map( A => n116529, Z => n119857);
   U83631 : BUF_X1 port map( A => n116529, Z => n119858);
   U83632 : BUF_X1 port map( A => n116529, Z => n119859);
   U83633 : BUF_X1 port map( A => n116529, Z => n119860);
   U83634 : BUF_X1 port map( A => n114693, Z => n120082);
   U83635 : BUF_X1 port map( A => n114700, Z => n120058);
   U83636 : BUF_X1 port map( A => n116529, Z => n119856);
   U83637 : BUF_X1 port map( A => n114693, Z => n120078);
   U83638 : BUF_X1 port map( A => n114700, Z => n120054);
   U83639 : BUF_X1 port map( A => n114693, Z => n120079);
   U83640 : BUF_X1 port map( A => n114700, Z => n120055);
   U83641 : BUF_X1 port map( A => n114693, Z => n120080);
   U83642 : BUF_X1 port map( A => n114700, Z => n120056);
   U83643 : BUF_X1 port map( A => n114693, Z => n120081);
   U83644 : BUF_X1 port map( A => n114700, Z => n120057);
   U83645 : BUF_X1 port map( A => n116492, Z => n120013);
   U83646 : BUF_X1 port map( A => n116499, Z => n119989);
   U83647 : BUF_X1 port map( A => n116487, Z => n120037);
   U83648 : BUF_X1 port map( A => n116504, Z => n119965);
   U83649 : BUF_X1 port map( A => n116492, Z => n120014);
   U83650 : BUF_X1 port map( A => n116499, Z => n119990);
   U83651 : BUF_X1 port map( A => n116487, Z => n120038);
   U83652 : BUF_X1 port map( A => n116504, Z => n119966);
   U83653 : BUF_X1 port map( A => n116492, Z => n120015);
   U83654 : BUF_X1 port map( A => n116499, Z => n119991);
   U83655 : BUF_X1 port map( A => n116487, Z => n120039);
   U83656 : BUF_X1 port map( A => n116504, Z => n119967);
   U83657 : BUF_X1 port map( A => n116492, Z => n120016);
   U83658 : BUF_X1 port map( A => n116499, Z => n119992);
   U83659 : BUF_X1 port map( A => n116487, Z => n120040);
   U83660 : BUF_X1 port map( A => n116504, Z => n119968);
   U83661 : BUF_X1 port map( A => n114672, Z => n120166);
   U83662 : BUF_X1 port map( A => n114672, Z => n120163);
   U83663 : BUF_X1 port map( A => n114672, Z => n120164);
   U83664 : BUF_X1 port map( A => n114672, Z => n120165);
   U83665 : BUF_X1 port map( A => n114654, Z => n120238);
   U83666 : BUF_X1 port map( A => n114654, Z => n120235);
   U83667 : BUF_X1 port map( A => n114654, Z => n120236);
   U83668 : BUF_X1 port map( A => n114654, Z => n120237);
   U83669 : BUF_X1 port map( A => n114659, Z => n120214);
   U83670 : BUF_X1 port map( A => n114666, Z => n120190);
   U83671 : BUF_X1 port map( A => n114659, Z => n120211);
   U83672 : BUF_X1 port map( A => n114666, Z => n120187);
   U83673 : BUF_X1 port map( A => n114659, Z => n120212);
   U83674 : BUF_X1 port map( A => n114666, Z => n120188);
   U83675 : BUF_X1 port map( A => n114659, Z => n120213);
   U83676 : BUF_X1 port map( A => n114666, Z => n120189);
   U83677 : BUF_X1 port map( A => n114690, Z => n120094);
   U83678 : BUF_X1 port map( A => n114690, Z => n120090);
   U83679 : BUF_X1 port map( A => n114690, Z => n120091);
   U83680 : BUF_X1 port map( A => n114690, Z => n120092);
   U83681 : BUF_X1 port map( A => n114690, Z => n120093);
   U83682 : BUF_X1 port map( A => n116521, Z => n119893);
   U83683 : BUF_X1 port map( A => n116521, Z => n119894);
   U83684 : BUF_X1 port map( A => n116521, Z => n119895);
   U83685 : BUF_X1 port map( A => n116521, Z => n119896);
   U83686 : BUF_X1 port map( A => n116521, Z => n119892);
   U83687 : BUF_X1 port map( A => n114688, Z => n120106);
   U83688 : BUF_X1 port map( A => n114688, Z => n120102);
   U83689 : BUF_X1 port map( A => n114688, Z => n120103);
   U83690 : BUF_X1 port map( A => n114688, Z => n120104);
   U83691 : BUF_X1 port map( A => n114688, Z => n120105);
   U83692 : BUF_X1 port map( A => n116519, Z => n119905);
   U83693 : BUF_X1 port map( A => n116519, Z => n119906);
   U83694 : BUF_X1 port map( A => n116519, Z => n119907);
   U83695 : BUF_X1 port map( A => n116519, Z => n119908);
   U83696 : BUF_X1 port map( A => n116519, Z => n119904);
   U83697 : BUF_X1 port map( A => n116520, Z => n119899);
   U83698 : BUF_X1 port map( A => n116520, Z => n119900);
   U83699 : BUF_X1 port map( A => n116520, Z => n119901);
   U83700 : BUF_X1 port map( A => n116520, Z => n119902);
   U83701 : BUF_X1 port map( A => n116520, Z => n119898);
   U83702 : BUF_X1 port map( A => n114670, Z => n120172);
   U83703 : BUF_X1 port map( A => n114676, Z => n120148);
   U83704 : BUF_X1 port map( A => n114670, Z => n120168);
   U83705 : BUF_X1 port map( A => n114676, Z => n120144);
   U83706 : BUF_X1 port map( A => n114670, Z => n120169);
   U83707 : BUF_X1 port map( A => n114676, Z => n120145);
   U83708 : BUF_X1 port map( A => n114670, Z => n120170);
   U83709 : BUF_X1 port map( A => n114676, Z => n120146);
   U83710 : BUF_X1 port map( A => n114670, Z => n120171);
   U83711 : BUF_X1 port map( A => n114676, Z => n120147);
   U83712 : BUF_X1 port map( A => n116497, Z => n119995);
   U83713 : BUF_X1 port map( A => n116503, Z => n119971);
   U83714 : BUF_X1 port map( A => n116508, Z => n119947);
   U83715 : BUF_X1 port map( A => n116497, Z => n119996);
   U83716 : BUF_X1 port map( A => n116503, Z => n119972);
   U83717 : BUF_X1 port map( A => n116508, Z => n119948);
   U83718 : BUF_X1 port map( A => n116497, Z => n119997);
   U83719 : BUF_X1 port map( A => n116503, Z => n119973);
   U83720 : BUF_X1 port map( A => n116508, Z => n119949);
   U83721 : BUF_X1 port map( A => n116497, Z => n119998);
   U83722 : BUF_X1 port map( A => n116503, Z => n119974);
   U83723 : BUF_X1 port map( A => n116508, Z => n119950);
   U83724 : BUF_X1 port map( A => n114664, Z => n120196);
   U83725 : BUF_X1 port map( A => n116497, Z => n119994);
   U83726 : BUF_X1 port map( A => n116503, Z => n119970);
   U83727 : BUF_X1 port map( A => n116508, Z => n119946);
   U83728 : BUF_X1 port map( A => n114664, Z => n120192);
   U83729 : BUF_X1 port map( A => n114664, Z => n120193);
   U83730 : BUF_X1 port map( A => n114664, Z => n120194);
   U83731 : BUF_X1 port map( A => n114664, Z => n120195);
   U83732 : NAND2_X1 port map( A1 => n120628, A2 => n120248, ZN => n114645);
   U83733 : NAND2_X1 port map( A1 => n120628, A2 => n120617, ZN => n113897);
   U83734 : NAND2_X1 port map( A1 => n120628, A2 => n120605, ZN => n113904);
   U83735 : BUF_X1 port map( A => n114213, Z => n120389);
   U83736 : BUF_X1 port map( A => n114132, Z => n120470);
   U83737 : BUF_X1 port map( A => n114136, Z => n120446);
   U83738 : BUF_X1 port map( A => n114128, Z => n120494);
   U83739 : BUF_X1 port map( A => n114130, Z => n120482);
   U83740 : BUF_X1 port map( A => n114134, Z => n120458);
   U83741 : BUF_X1 port map( A => n113911, Z => n120581);
   U83742 : BUF_X1 port map( A => n114122, Z => n120506);
   U83743 : BUF_X1 port map( A => n113980, Z => n120556);
   U83744 : BUF_X1 port map( A => n113909, Z => n120593);
   U83745 : BUF_X1 port map( A => n114300, Z => n120360);
   U83746 : BUF_X1 port map( A => n114211, Z => n120397);
   U83747 : BUF_X1 port map( A => n114372, Z => n120323);
   U83748 : BUF_X1 port map( A => n114575, Z => n120272);
   U83749 : BUF_X1 port map( A => n114142, Z => n120422);
   U83750 : BUF_X1 port map( A => n114303, Z => n120348);
   U83751 : BUF_X1 port map( A => n114213, Z => n120385);
   U83752 : BUF_X1 port map( A => n114052, Z => n120531);
   U83753 : BUF_X1 port map( A => n113895, Z => n120617);
   U83754 : BUF_X1 port map( A => n113902, Z => n120605);
   U83755 : BUF_X1 port map( A => n114132, Z => n120471);
   U83756 : BUF_X1 port map( A => n114132, Z => n120472);
   U83757 : BUF_X1 port map( A => n114132, Z => n120473);
   U83758 : BUF_X1 port map( A => n114132, Z => n120474);
   U83759 : BUF_X1 port map( A => n114136, Z => n120447);
   U83760 : BUF_X1 port map( A => n114136, Z => n120448);
   U83761 : BUF_X1 port map( A => n114136, Z => n120449);
   U83762 : BUF_X1 port map( A => n114136, Z => n120450);
   U83763 : BUF_X1 port map( A => n114128, Z => n120495);
   U83764 : BUF_X1 port map( A => n114128, Z => n120496);
   U83765 : BUF_X1 port map( A => n114128, Z => n120497);
   U83766 : BUF_X1 port map( A => n114128, Z => n120498);
   U83767 : BUF_X1 port map( A => n114130, Z => n120483);
   U83768 : BUF_X1 port map( A => n114130, Z => n120484);
   U83769 : BUF_X1 port map( A => n114130, Z => n120485);
   U83770 : BUF_X1 port map( A => n114130, Z => n120486);
   U83771 : BUF_X1 port map( A => n114134, Z => n120459);
   U83772 : BUF_X1 port map( A => n114134, Z => n120460);
   U83773 : BUF_X1 port map( A => n114134, Z => n120461);
   U83774 : BUF_X1 port map( A => n114134, Z => n120462);
   U83775 : BUF_X1 port map( A => n113911, Z => n120582);
   U83776 : BUF_X1 port map( A => n113911, Z => n120583);
   U83777 : BUF_X1 port map( A => n113911, Z => n120584);
   U83778 : BUF_X1 port map( A => n113911, Z => n120585);
   U83779 : BUF_X1 port map( A => n114122, Z => n120507);
   U83780 : BUF_X1 port map( A => n114122, Z => n120508);
   U83781 : BUF_X1 port map( A => n114122, Z => n120509);
   U83782 : BUF_X1 port map( A => n114122, Z => n120510);
   U83783 : BUF_X1 port map( A => n113980, Z => n120557);
   U83784 : BUF_X1 port map( A => n113980, Z => n120558);
   U83785 : BUF_X1 port map( A => n113980, Z => n120559);
   U83786 : BUF_X1 port map( A => n113980, Z => n120560);
   U83787 : BUF_X1 port map( A => n113909, Z => n120594);
   U83788 : BUF_X1 port map( A => n113909, Z => n120595);
   U83789 : BUF_X1 port map( A => n113909, Z => n120596);
   U83790 : BUF_X1 port map( A => n113909, Z => n120597);
   U83791 : BUF_X1 port map( A => n114300, Z => n120361);
   U83792 : BUF_X1 port map( A => n114300, Z => n120362);
   U83793 : BUF_X1 port map( A => n114300, Z => n120363);
   U83794 : BUF_X1 port map( A => n114300, Z => n120364);
   U83795 : BUF_X1 port map( A => n114211, Z => n120398);
   U83796 : BUF_X1 port map( A => n114211, Z => n120399);
   U83797 : BUF_X1 port map( A => n114211, Z => n120400);
   U83798 : BUF_X1 port map( A => n114211, Z => n120401);
   U83799 : BUF_X1 port map( A => n114372, Z => n120324);
   U83800 : BUF_X1 port map( A => n114372, Z => n120325);
   U83801 : BUF_X1 port map( A => n114372, Z => n120326);
   U83802 : BUF_X1 port map( A => n114372, Z => n120327);
   U83803 : BUF_X1 port map( A => n114575, Z => n120273);
   U83804 : BUF_X1 port map( A => n114575, Z => n120274);
   U83805 : BUF_X1 port map( A => n114575, Z => n120275);
   U83806 : BUF_X1 port map( A => n114575, Z => n120276);
   U83807 : BUF_X1 port map( A => n114213, Z => n120386);
   U83808 : BUF_X1 port map( A => n114142, Z => n120423);
   U83809 : BUF_X1 port map( A => n114142, Z => n120424);
   U83810 : BUF_X1 port map( A => n114142, Z => n120425);
   U83811 : BUF_X1 port map( A => n114142, Z => n120426);
   U83812 : BUF_X1 port map( A => n114303, Z => n120349);
   U83813 : BUF_X1 port map( A => n114303, Z => n120350);
   U83814 : BUF_X1 port map( A => n114303, Z => n120351);
   U83815 : BUF_X1 port map( A => n114303, Z => n120352);
   U83816 : BUF_X1 port map( A => n114213, Z => n120387);
   U83817 : BUF_X1 port map( A => n114052, Z => n120532);
   U83818 : BUF_X1 port map( A => n114052, Z => n120533);
   U83819 : BUF_X1 port map( A => n114052, Z => n120534);
   U83820 : BUF_X1 port map( A => n114052, Z => n120535);
   U83821 : BUF_X1 port map( A => n113895, Z => n120618);
   U83822 : BUF_X1 port map( A => n113895, Z => n120619);
   U83823 : BUF_X1 port map( A => n113895, Z => n120620);
   U83824 : BUF_X1 port map( A => n113895, Z => n120621);
   U83825 : BUF_X1 port map( A => n113902, Z => n120606);
   U83826 : BUF_X1 port map( A => n113902, Z => n120607);
   U83827 : BUF_X1 port map( A => n113902, Z => n120608);
   U83828 : BUF_X1 port map( A => n113902, Z => n120609);
   U83829 : BUF_X1 port map( A => n116513, Z => n119941);
   U83830 : BUF_X1 port map( A => n116515, Z => n119929);
   U83831 : BUF_X1 port map( A => n116517, Z => n119917);
   U83832 : BUF_X1 port map( A => n116513, Z => n119942);
   U83833 : BUF_X1 port map( A => n116515, Z => n119930);
   U83834 : BUF_X1 port map( A => n116517, Z => n119918);
   U83835 : BUF_X1 port map( A => n116513, Z => n119943);
   U83836 : BUF_X1 port map( A => n116515, Z => n119931);
   U83837 : BUF_X1 port map( A => n116517, Z => n119919);
   U83838 : BUF_X1 port map( A => n116513, Z => n119944);
   U83839 : BUF_X1 port map( A => n116515, Z => n119932);
   U83840 : BUF_X1 port map( A => n116517, Z => n119920);
   U83841 : BUF_X1 port map( A => n114686, Z => n120118);
   U83842 : BUF_X1 port map( A => n114686, Z => n120114);
   U83843 : BUF_X1 port map( A => n114696, Z => n120072);
   U83844 : BUF_X1 port map( A => n114686, Z => n120115);
   U83845 : BUF_X1 port map( A => n114684, Z => n120130);
   U83846 : BUF_X1 port map( A => n114682, Z => n120142);
   U83847 : BUF_X1 port map( A => n114696, Z => n120076);
   U83848 : BUF_X1 port map( A => n116513, Z => n119940);
   U83849 : BUF_X1 port map( A => n116515, Z => n119928);
   U83850 : BUF_X1 port map( A => n116517, Z => n119916);
   U83851 : BUF_X1 port map( A => n114684, Z => n120126);
   U83852 : BUF_X1 port map( A => n114682, Z => n120138);
   U83853 : BUF_X1 port map( A => n114684, Z => n120127);
   U83854 : BUF_X1 port map( A => n114682, Z => n120139);
   U83855 : BUF_X1 port map( A => n114696, Z => n120073);
   U83856 : BUF_X1 port map( A => n114686, Z => n120116);
   U83857 : BUF_X1 port map( A => n114686, Z => n120117);
   U83858 : BUF_X1 port map( A => n114684, Z => n120128);
   U83859 : BUF_X1 port map( A => n114682, Z => n120140);
   U83860 : BUF_X1 port map( A => n114696, Z => n120074);
   U83861 : BUF_X1 port map( A => n114684, Z => n120129);
   U83862 : BUF_X1 port map( A => n114682, Z => n120141);
   U83863 : BUF_X1 port map( A => n114696, Z => n120075);
   U83864 : BUF_X1 port map( A => n116531, Z => n119851);
   U83865 : BUF_X1 port map( A => n116526, Z => n119875);
   U83866 : BUF_X1 port map( A => n116531, Z => n119852);
   U83867 : BUF_X1 port map( A => n116526, Z => n119876);
   U83868 : BUF_X1 port map( A => n116531, Z => n119853);
   U83869 : BUF_X1 port map( A => n116526, Z => n119877);
   U83870 : BUF_X1 port map( A => n116531, Z => n119854);
   U83871 : BUF_X1 port map( A => n116526, Z => n119878);
   U83872 : BUF_X1 port map( A => n114702, Z => n120052);
   U83873 : BUF_X1 port map( A => n116531, Z => n119850);
   U83874 : BUF_X1 port map( A => n116526, Z => n119874);
   U83875 : BUF_X1 port map( A => n114702, Z => n120048);
   U83876 : BUF_X1 port map( A => n114702, Z => n120049);
   U83877 : BUF_X1 port map( A => n114702, Z => n120050);
   U83878 : BUF_X1 port map( A => n114702, Z => n120051);
   U83879 : BUF_X1 port map( A => n114213, Z => n120388);
   U83880 : NAND2_X1 port map( A1 => n120625, A2 => n120360, ZN => n114301);
   U83881 : NAND2_X1 port map( A1 => n120625, A2 => n120374, ZN => n114236);
   U83882 : NAND2_X1 port map( A1 => n120625, A2 => n120411, ZN => n114147);
   U83883 : NAND2_X1 port map( A1 => n120625, A2 => n120385, ZN => n114214);
   U83884 : NAND2_X1 port map( A1 => n120626, A2 => n120506, ZN => n114124);
   U83885 : NAND2_X1 port map( A1 => n120627, A2 => n120556, ZN => n113982);
   U83886 : NAND2_X1 port map( A1 => n120626, A2 => n120470, ZN => n114133);
   U83887 : NAND2_X1 port map( A1 => n120626, A2 => n120446, ZN => n114137);
   U83888 : NAND2_X1 port map( A1 => n120627, A2 => n120520, ZN => n114057);
   U83889 : NAND2_X1 port map( A1 => n120626, A2 => n120494, ZN => n114129);
   U83890 : NAND2_X1 port map( A1 => n120626, A2 => n120482, ZN => n114131);
   U83891 : NAND2_X1 port map( A1 => n120626, A2 => n120458, ZN => n114135);
   U83892 : NAND2_X1 port map( A1 => n120627, A2 => n120581, ZN => n113912);
   U83893 : NAND2_X1 port map( A1 => n120627, A2 => n120593, ZN => n113910);
   U83894 : NAND2_X1 port map( A1 => n120627, A2 => n120570, ZN => n113916);
   U83895 : NAND2_X1 port map( A1 => n120626, A2 => n120337, ZN => n114307);
   U83896 : NAND2_X1 port map( A1 => n120626, A2 => n120397, ZN => n114212);
   U83897 : NAND2_X1 port map( A1 => n120627, A2 => n120323, ZN => n114373);
   U83898 : NAND2_X1 port map( A1 => n120627, A2 => n120286, ZN => n114511);
   U83899 : NAND2_X1 port map( A1 => n120627, A2 => n120272, ZN => n114576);
   U83900 : NAND2_X1 port map( A1 => n120627, A2 => n120261, ZN => n114579);
   U83901 : NAND2_X1 port map( A1 => n120627, A2 => n120545, ZN => n113991);
   U83902 : NAND2_X1 port map( A1 => n120626, A2 => n120434, ZN => n114140);
   U83903 : NAND2_X1 port map( A1 => n120626, A2 => n120422, ZN => n114143);
   U83904 : NAND2_X1 port map( A1 => n120626, A2 => n120348, ZN => n114304);
   U83905 : NAND2_X1 port map( A1 => n120627, A2 => n120299, ZN => n114445);
   U83906 : NAND2_X1 port map( A1 => n120627, A2 => n120531, ZN => n114053);
   U83907 : NAND2_X1 port map( A1 => n120626, A2 => n120312, ZN => n114379);
   U83908 : BUF_X1 port map( A => n116514, Z => n119935);
   U83909 : BUF_X1 port map( A => n116518, Z => n119911);
   U83910 : BUF_X1 port map( A => n116514, Z => n119936);
   U83911 : BUF_X1 port map( A => n116518, Z => n119912);
   U83912 : BUF_X1 port map( A => n116514, Z => n119937);
   U83913 : BUF_X1 port map( A => n116518, Z => n119913);
   U83914 : BUF_X1 port map( A => n116514, Z => n119938);
   U83915 : BUF_X1 port map( A => n116518, Z => n119914);
   U83916 : BUF_X1 port map( A => n114685, Z => n120124);
   U83917 : BUF_X1 port map( A => n114685, Z => n120120);
   U83918 : BUF_X1 port map( A => n114685, Z => n120121);
   U83919 : BUF_X1 port map( A => n114685, Z => n120122);
   U83920 : BUF_X1 port map( A => n114685, Z => n120123);
   U83921 : BUF_X1 port map( A => n114683, Z => n120136);
   U83922 : BUF_X1 port map( A => n114703, Z => n120046);
   U83923 : BUF_X1 port map( A => n116514, Z => n119934);
   U83924 : BUF_X1 port map( A => n116518, Z => n119910);
   U83925 : BUF_X1 port map( A => n114683, Z => n120132);
   U83926 : BUF_X1 port map( A => n114703, Z => n120042);
   U83927 : BUF_X1 port map( A => n114683, Z => n120133);
   U83928 : BUF_X1 port map( A => n114703, Z => n120043);
   U83929 : BUF_X1 port map( A => n114683, Z => n120134);
   U83930 : BUF_X1 port map( A => n114703, Z => n120044);
   U83931 : BUF_X1 port map( A => n114683, Z => n120135);
   U83932 : BUF_X1 port map( A => n114703, Z => n120045);
   U83933 : BUF_X1 port map( A => n116516, Z => n119923);
   U83934 : BUF_X1 port map( A => n116532, Z => n119845);
   U83935 : BUF_X1 port map( A => n116527, Z => n119869);
   U83936 : BUF_X1 port map( A => n116516, Z => n119924);
   U83937 : BUF_X1 port map( A => n116532, Z => n119846);
   U83938 : BUF_X1 port map( A => n116527, Z => n119870);
   U83939 : BUF_X1 port map( A => n116516, Z => n119925);
   U83940 : BUF_X1 port map( A => n116532, Z => n119847);
   U83941 : BUF_X1 port map( A => n116527, Z => n119871);
   U83942 : BUF_X1 port map( A => n116516, Z => n119926);
   U83943 : BUF_X1 port map( A => n116532, Z => n119848);
   U83944 : BUF_X1 port map( A => n116527, Z => n119872);
   U83945 : BUF_X1 port map( A => n114687, Z => n120112);
   U83946 : BUF_X1 port map( A => n114697, Z => n120070);
   U83947 : BUF_X1 port map( A => n116516, Z => n119922);
   U83948 : BUF_X1 port map( A => n116532, Z => n119844);
   U83949 : BUF_X1 port map( A => n116527, Z => n119868);
   U83950 : BUF_X1 port map( A => n114687, Z => n120108);
   U83951 : BUF_X1 port map( A => n114697, Z => n120066);
   U83952 : BUF_X1 port map( A => n114687, Z => n120109);
   U83953 : BUF_X1 port map( A => n114697, Z => n120067);
   U83954 : BUF_X1 port map( A => n114687, Z => n120110);
   U83955 : BUF_X1 port map( A => n114697, Z => n120068);
   U83956 : BUF_X1 port map( A => n114687, Z => n120111);
   U83957 : BUF_X1 port map( A => n114697, Z => n120069);
   U83958 : BUF_X1 port map( A => n116493, Z => n120007);
   U83959 : BUF_X1 port map( A => n116488, Z => n120031);
   U83960 : BUF_X1 port map( A => n116505, Z => n119959);
   U83961 : BUF_X1 port map( A => n116493, Z => n120008);
   U83962 : BUF_X1 port map( A => n116488, Z => n120032);
   U83963 : BUF_X1 port map( A => n116505, Z => n119960);
   U83964 : BUF_X1 port map( A => n116493, Z => n120009);
   U83965 : BUF_X1 port map( A => n116488, Z => n120033);
   U83966 : BUF_X1 port map( A => n116505, Z => n119961);
   U83967 : BUF_X1 port map( A => n116493, Z => n120010);
   U83968 : BUF_X1 port map( A => n116488, Z => n120034);
   U83969 : BUF_X1 port map( A => n116505, Z => n119962);
   U83970 : BUF_X1 port map( A => n114655, Z => n120232);
   U83971 : BUF_X1 port map( A => n114667, Z => n120184);
   U83972 : BUF_X1 port map( A => n116493, Z => n120006);
   U83973 : BUF_X1 port map( A => n116488, Z => n120030);
   U83974 : BUF_X1 port map( A => n116505, Z => n119958);
   U83975 : BUF_X1 port map( A => n114655, Z => n120228);
   U83976 : BUF_X1 port map( A => n114667, Z => n120180);
   U83977 : BUF_X1 port map( A => n114655, Z => n120229);
   U83978 : BUF_X1 port map( A => n114667, Z => n120181);
   U83979 : BUF_X1 port map( A => n114655, Z => n120230);
   U83980 : BUF_X1 port map( A => n114667, Z => n120182);
   U83981 : BUF_X1 port map( A => n114655, Z => n120231);
   U83982 : BUF_X1 port map( A => n114667, Z => n120183);
   U83983 : BUF_X1 port map( A => n116500, Z => n119983);
   U83984 : BUF_X1 port map( A => n116500, Z => n119984);
   U83985 : BUF_X1 port map( A => n116500, Z => n119985);
   U83986 : BUF_X1 port map( A => n116500, Z => n119986);
   U83987 : BUF_X1 port map( A => n114660, Z => n120208);
   U83988 : BUF_X1 port map( A => n114673, Z => n120160);
   U83989 : BUF_X1 port map( A => n116500, Z => n119982);
   U83990 : BUF_X1 port map( A => n114660, Z => n120204);
   U83991 : BUF_X1 port map( A => n114673, Z => n120156);
   U83992 : BUF_X1 port map( A => n114660, Z => n120205);
   U83993 : BUF_X1 port map( A => n114673, Z => n120157);
   U83994 : BUF_X1 port map( A => n114660, Z => n120206);
   U83995 : BUF_X1 port map( A => n114673, Z => n120158);
   U83996 : BUF_X1 port map( A => n114660, Z => n120207);
   U83997 : BUF_X1 port map( A => n114673, Z => n120159);
   U83998 : BUF_X1 port map( A => n114672, Z => n120162);
   U83999 : BUF_X1 port map( A => n116492, Z => n120012);
   U84000 : BUF_X1 port map( A => n116499, Z => n119988);
   U84001 : BUF_X1 port map( A => n116487, Z => n120036);
   U84002 : BUF_X1 port map( A => n116504, Z => n119964);
   U84003 : BUF_X1 port map( A => n114654, Z => n120234);
   U84004 : BUF_X1 port map( A => n114659, Z => n120210);
   U84005 : BUF_X1 port map( A => n114666, Z => n120186);
   U84006 : NAND2_X1 port map( A1 => n120628, A2 => n120829, ZN => n113767);
   U84007 : OAI21_X1 port map( B1 => n113893, B2 => n113894, A => n120623, ZN 
                           => n113766);
   U84008 : AND2_X1 port map( A1 => n117949, A2 => n117948, ZN => n116528);
   U84009 : BUF_X1 port map( A => n113914, Z => n120568);
   U84010 : BUF_X1 port map( A => n113990, Z => n120543);
   U84011 : BUF_X1 port map( A => n114643, Z => n120246);
   U84012 : BUF_X1 port map( A => n114577, Z => n120259);
   U84013 : BUF_X1 port map( A => n114055, Z => n120518);
   U84014 : BUF_X1 port map( A => n114234, Z => n120372);
   U84015 : BUF_X1 port map( A => n114305, Z => n120335);
   U84016 : BUF_X1 port map( A => n114509, Z => n120284);
   U84017 : BUF_X1 port map( A => n114145, Z => n120409);
   U84018 : BUF_X1 port map( A => n114377, Z => n120310);
   U84019 : BUF_X1 port map( A => n114443, Z => n120297);
   U84020 : BUF_X1 port map( A => n113990, Z => n120544);
   U84021 : BUF_X1 port map( A => n113914, Z => n120569);
   U84022 : BUF_X1 port map( A => n114643, Z => n120247);
   U84023 : BUF_X1 port map( A => n114055, Z => n120519);
   U84024 : BUF_X1 port map( A => n114234, Z => n120373);
   U84025 : BUF_X1 port map( A => n114305, Z => n120336);
   U84026 : BUF_X1 port map( A => n114509, Z => n120285);
   U84027 : BUF_X1 port map( A => n114577, Z => n120260);
   U84028 : BUF_X1 port map( A => n114145, Z => n120410);
   U84029 : BUF_X1 port map( A => n114443, Z => n120298);
   U84030 : BUF_X1 port map( A => n114377, Z => n120311);
   U84031 : NOR3_X1 port map( A1 => n116478, A2 => n120216, A3 => n116475, ZN 
                           => n116447);
   U84032 : NOR3_X1 port map( A1 => n116470, A2 => n116469, A3 => n116471, ZN 
                           => n116463);
   U84033 : NOR3_X1 port map( A1 => n117967, A2 => n117970, A3 => n117958, ZN 
                           => n117949);
   U84034 : OAI21_X1 port map( B1 => n113901, B2 => n113908, A => n120623, ZN 
                           => n113909);
   U84035 : OAI21_X1 port map( B1 => n113908, B2 => n114054, A => n120623, ZN 
                           => n114122);
   U84036 : OAI21_X1 port map( B1 => n113913, B2 => n114121, A => n120624, ZN 
                           => n114132);
   U84037 : OAI21_X1 port map( B1 => n113986, B2 => n114121, A => n120624, ZN 
                           => n114136);
   U84038 : OAI21_X1 port map( B1 => n113908, B2 => n114121, A => n120623, ZN 
                           => n114128);
   U84039 : OAI21_X1 port map( B1 => n113913, B2 => n114054, A => n120624, ZN 
                           => n114130);
   U84040 : OAI21_X1 port map( B1 => n113986, B2 => n114054, A => n120624, ZN 
                           => n114134);
   U84041 : OAI21_X1 port map( B1 => n113986, B2 => n114141, A => n120625, ZN 
                           => n114300);
   U84042 : OAI21_X1 port map( B1 => n113908, B2 => n114144, A => n120624, ZN 
                           => n114211);
   U84043 : OAI21_X1 port map( B1 => n113894, B2 => n114374, A => n120625, ZN 
                           => n114372);
   U84044 : OAI21_X1 port map( B1 => n113913, B2 => n114374, A => n120624, ZN 
                           => n114575);
   U84045 : OAI21_X1 port map( B1 => n113913, B2 => n114141, A => n120624, ZN 
                           => n114213);
   U84046 : OAI21_X1 port map( B1 => n113894, B2 => n114144, A => n120624, ZN 
                           => n114142);
   U84047 : OAI21_X1 port map( B1 => n113986, B2 => n114144, A => n120625, ZN 
                           => n114303);
   U84048 : OAI21_X1 port map( B1 => n113894, B2 => n114054, A => n120623, ZN 
                           => n114052);
   U84049 : OAI21_X1 port map( B1 => n113893, B2 => n113986, A => n120623, ZN 
                           => n113980);
   U84050 : OAI21_X1 port map( B1 => n113893, B2 => n113908, A => n120623, ZN 
                           => n113902);
   U84051 : OAI21_X1 port map( B1 => n113893, B2 => n113913, A => n120623, ZN 
                           => n113911);
   U84052 : OAI21_X1 port map( B1 => n113894, B2 => n113901, A => n120623, ZN 
                           => n113895);
   U84053 : BUF_X1 port map( A => n114658, Z => n120216);
   U84054 : BUF_X1 port map( A => n116491, Z => n120018);
   U84055 : BUF_X1 port map( A => n116491, Z => n120021);
   U84056 : BUF_X1 port map( A => n116491, Z => n120019);
   U84057 : BUF_X1 port map( A => n116491, Z => n120020);
   U84058 : BUF_X1 port map( A => n114658, Z => n120219);
   U84059 : BUF_X1 port map( A => n114658, Z => n120218);
   U84060 : BUF_X1 port map( A => n114658, Z => n120217);
   U84061 : NAND2_X1 port map( A1 => n116457, A2 => n116463, ZN => n114697);
   U84062 : NAND2_X1 port map( A1 => n116453, A2 => n116446, ZN => n114660);
   U84063 : NAND2_X1 port map( A1 => n116453, A2 => n116463, ZN => n114673);
   U84064 : NAND2_X1 port map( A1 => n116453, A2 => n116464, ZN => n114702);
   U84065 : NAND2_X1 port map( A1 => n117948, A2 => n117959, ZN => n116532);
   U84066 : NAND2_X1 port map( A1 => n117948, A2 => n117968, ZN => n116526);
   U84067 : NAND2_X1 port map( A1 => n117945, A2 => n117959, ZN => n116500);
   U84068 : NAND2_X1 port map( A1 => n117945, A2 => n117961, ZN => n116516);
   U84069 : NAND2_X1 port map( A1 => n117945, A2 => n117968, ZN => n116531);
   U84070 : NAND2_X1 port map( A1 => n117945, A2 => n117962, ZN => n116527);
   U84071 : NAND2_X1 port map( A1 => n114375, A2 => n114376, ZN => n113894);
   U84072 : NAND2_X1 port map( A1 => n116445, A2 => n116459, ZN => n114687);
   U84073 : BUF_X1 port map( A => n113892, Z => n120624);
   U84074 : BUF_X1 port map( A => n113892, Z => n120623);
   U84075 : BUF_X1 port map( A => n113892, Z => n120625);
   U84076 : BUF_X1 port map( A => n113892, Z => n120627);
   U84077 : BUF_X1 port map( A => n113892, Z => n120626);
   U84078 : NAND2_X1 port map( A1 => n116453, A2 => n116448, ZN => n114659);
   U84079 : NAND2_X1 port map( A1 => n116453, A2 => n116459, ZN => n114666);
   U84080 : NAND2_X1 port map( A1 => n116454, A2 => n116457, ZN => n114685);
   U84081 : NAND2_X1 port map( A1 => n116448, A2 => n116457, ZN => n114686);
   U84082 : NAND2_X1 port map( A1 => n116464, A2 => n116457, ZN => n114696);
   U84083 : NAND2_X1 port map( A1 => n116457, A2 => n116459, ZN => n114688);
   U84084 : NAND2_X1 port map( A1 => n116458, A2 => n116453, ZN => n114667);
   U84085 : NAND2_X1 port map( A1 => n116452, A2 => n116453, ZN => n114682);
   U84086 : NAND2_X1 port map( A1 => n117947, A2 => n117948, ZN => n116488);
   U84087 : NAND2_X1 port map( A1 => n117946, A2 => n117948, ZN => n116505);
   U84088 : NAND2_X1 port map( A1 => n117962, A2 => n117948, ZN => n116515);
   U84089 : NAND2_X1 port map( A1 => n117955, A2 => n117945, ZN => n116493);
   U84090 : NAND2_X1 port map( A1 => n117948, A2 => n117961, ZN => n116521);
   U84091 : NAND2_X1 port map( A1 => n117946, A2 => n117953, ZN => n116517);
   U84092 : NAND2_X1 port map( A1 => n117953, A2 => n117968, ZN => n116519);
   U84093 : OAI22_X1 port map( A1 => n113907, A2 => n120053, B1 => n114582, B2 
                           => n120047, ZN => n114781);
   U84094 : OAI22_X1 port map( A1 => n113906, A2 => n120053, B1 => n114581, B2 
                           => n120047, ZN => n114755);
   U84095 : OAI22_X1 port map( A1 => n113905, A2 => n120053, B1 => n114580, B2 
                           => n120047, ZN => n114729);
   U84096 : OAI22_X1 port map( A1 => n113903, A2 => n120053, B1 => n114578, B2 
                           => n120047, ZN => n114701);
   U84097 : NAND2_X1 port map( A1 => n116446, A2 => n116447, ZN => n114655);
   U84098 : NAND2_X1 port map( A1 => n116458, A2 => n116447, ZN => n114703);
   U84099 : NAND2_X1 port map( A1 => n117946, A2 => n117954, ZN => n116514);
   U84100 : NAND2_X1 port map( A1 => n117949, A2 => n117954, ZN => n116513);
   U84101 : NAND2_X1 port map( A1 => n117962, A2 => n117954, ZN => n116518);
   U84102 : NAND2_X1 port map( A1 => n116448, A2 => n116445, ZN => n114684);
   U84103 : NAND2_X1 port map( A1 => n117954, A2 => n117959, ZN => n116520);
   U84104 : NAND2_X1 port map( A1 => n116464, A2 => n116445, ZN => n114683);
   U84105 : BUF_X1 port map( A => n113891, Z => n120630);
   U84106 : BUF_X1 port map( A => n113889, Z => n120633);
   U84107 : BUF_X1 port map( A => n113887, Z => n120636);
   U84108 : BUF_X1 port map( A => n113885, Z => n120639);
   U84109 : BUF_X1 port map( A => n113883, Z => n120642);
   U84110 : BUF_X1 port map( A => n113881, Z => n120645);
   U84111 : BUF_X1 port map( A => n113879, Z => n120648);
   U84112 : BUF_X1 port map( A => n113877, Z => n120651);
   U84113 : BUF_X1 port map( A => n113875, Z => n120654);
   U84114 : BUF_X1 port map( A => n113873, Z => n120657);
   U84115 : BUF_X1 port map( A => n113871, Z => n120660);
   U84116 : BUF_X1 port map( A => n113869, Z => n120663);
   U84117 : BUF_X1 port map( A => n113867, Z => n120666);
   U84118 : BUF_X1 port map( A => n113865, Z => n120669);
   U84119 : BUF_X1 port map( A => n113863, Z => n120672);
   U84120 : BUF_X1 port map( A => n113861, Z => n120675);
   U84121 : BUF_X1 port map( A => n113859, Z => n120678);
   U84122 : BUF_X1 port map( A => n113857, Z => n120681);
   U84123 : BUF_X1 port map( A => n113855, Z => n120684);
   U84124 : BUF_X1 port map( A => n113853, Z => n120687);
   U84125 : BUF_X1 port map( A => n113851, Z => n120690);
   U84126 : BUF_X1 port map( A => n113849, Z => n120693);
   U84127 : BUF_X1 port map( A => n113847, Z => n120696);
   U84128 : BUF_X1 port map( A => n113845, Z => n120699);
   U84129 : BUF_X1 port map( A => n113843, Z => n120702);
   U84130 : BUF_X1 port map( A => n113841, Z => n120705);
   U84131 : BUF_X1 port map( A => n113839, Z => n120708);
   U84132 : BUF_X1 port map( A => n113837, Z => n120711);
   U84133 : BUF_X1 port map( A => n113835, Z => n120714);
   U84134 : BUF_X1 port map( A => n113833, Z => n120717);
   U84135 : BUF_X1 port map( A => n113831, Z => n120720);
   U84136 : BUF_X1 port map( A => n113829, Z => n120723);
   U84137 : BUF_X1 port map( A => n113827, Z => n120726);
   U84138 : BUF_X1 port map( A => n113825, Z => n120729);
   U84139 : BUF_X1 port map( A => n113823, Z => n120732);
   U84140 : BUF_X1 port map( A => n113821, Z => n120735);
   U84141 : BUF_X1 port map( A => n113819, Z => n120738);
   U84142 : BUF_X1 port map( A => n113817, Z => n120741);
   U84143 : BUF_X1 port map( A => n113815, Z => n120744);
   U84144 : BUF_X1 port map( A => n113813, Z => n120747);
   U84145 : BUF_X1 port map( A => n113811, Z => n120750);
   U84146 : BUF_X1 port map( A => n113809, Z => n120753);
   U84147 : BUF_X1 port map( A => n113807, Z => n120756);
   U84148 : BUF_X1 port map( A => n113805, Z => n120759);
   U84149 : BUF_X1 port map( A => n113803, Z => n120762);
   U84150 : BUF_X1 port map( A => n113801, Z => n120765);
   U84151 : BUF_X1 port map( A => n113799, Z => n120768);
   U84152 : BUF_X1 port map( A => n113797, Z => n120771);
   U84153 : BUF_X1 port map( A => n113795, Z => n120774);
   U84154 : BUF_X1 port map( A => n113793, Z => n120777);
   U84155 : BUF_X1 port map( A => n113791, Z => n120780);
   U84156 : BUF_X1 port map( A => n113789, Z => n120783);
   U84157 : BUF_X1 port map( A => n113787, Z => n120786);
   U84158 : BUF_X1 port map( A => n113785, Z => n120789);
   U84159 : BUF_X1 port map( A => n113783, Z => n120792);
   U84160 : BUF_X1 port map( A => n113781, Z => n120795);
   U84161 : BUF_X1 port map( A => n113779, Z => n120798);
   U84162 : BUF_X1 port map( A => n113777, Z => n120801);
   U84163 : BUF_X1 port map( A => n113775, Z => n120804);
   U84164 : BUF_X1 port map( A => n113773, Z => n120807);
   U84165 : BUF_X1 port map( A => n113771, Z => n120810);
   U84166 : BUF_X1 port map( A => n113770, Z => n120813);
   U84167 : BUF_X1 port map( A => n113769, Z => n120816);
   U84168 : BUF_X1 port map( A => n113768, Z => n120819);
   U84169 : BUF_X1 port map( A => n116491, Z => n120022);
   U84170 : BUF_X1 port map( A => n114658, Z => n120220);
   U84171 : BUF_X1 port map( A => n113771, Z => n120809);
   U84172 : BUF_X1 port map( A => n113770, Z => n120812);
   U84173 : BUF_X1 port map( A => n113769, Z => n120815);
   U84174 : BUF_X1 port map( A => n113768, Z => n120818);
   U84175 : BUF_X1 port map( A => n113891, Z => n120629);
   U84176 : BUF_X1 port map( A => n113889, Z => n120632);
   U84177 : BUF_X1 port map( A => n113887, Z => n120635);
   U84178 : BUF_X1 port map( A => n113885, Z => n120638);
   U84179 : BUF_X1 port map( A => n113883, Z => n120641);
   U84180 : BUF_X1 port map( A => n113881, Z => n120644);
   U84181 : BUF_X1 port map( A => n113879, Z => n120647);
   U84182 : BUF_X1 port map( A => n113877, Z => n120650);
   U84183 : BUF_X1 port map( A => n113875, Z => n120653);
   U84184 : BUF_X1 port map( A => n113873, Z => n120656);
   U84185 : BUF_X1 port map( A => n113871, Z => n120659);
   U84186 : BUF_X1 port map( A => n113869, Z => n120662);
   U84187 : BUF_X1 port map( A => n113867, Z => n120665);
   U84188 : BUF_X1 port map( A => n113865, Z => n120668);
   U84189 : BUF_X1 port map( A => n113863, Z => n120671);
   U84190 : BUF_X1 port map( A => n113861, Z => n120674);
   U84191 : BUF_X1 port map( A => n113859, Z => n120677);
   U84192 : BUF_X1 port map( A => n113857, Z => n120680);
   U84193 : BUF_X1 port map( A => n113855, Z => n120683);
   U84194 : BUF_X1 port map( A => n113853, Z => n120686);
   U84195 : BUF_X1 port map( A => n113851, Z => n120689);
   U84196 : BUF_X1 port map( A => n113849, Z => n120692);
   U84197 : BUF_X1 port map( A => n113847, Z => n120695);
   U84198 : BUF_X1 port map( A => n113845, Z => n120698);
   U84199 : BUF_X1 port map( A => n113843, Z => n120701);
   U84200 : BUF_X1 port map( A => n113841, Z => n120704);
   U84201 : BUF_X1 port map( A => n113839, Z => n120707);
   U84202 : BUF_X1 port map( A => n113837, Z => n120710);
   U84203 : BUF_X1 port map( A => n113835, Z => n120713);
   U84204 : BUF_X1 port map( A => n113833, Z => n120716);
   U84205 : BUF_X1 port map( A => n113831, Z => n120719);
   U84206 : BUF_X1 port map( A => n113829, Z => n120722);
   U84207 : BUF_X1 port map( A => n113827, Z => n120725);
   U84208 : BUF_X1 port map( A => n113825, Z => n120728);
   U84209 : BUF_X1 port map( A => n113823, Z => n120731);
   U84210 : BUF_X1 port map( A => n113821, Z => n120734);
   U84211 : BUF_X1 port map( A => n113819, Z => n120737);
   U84212 : BUF_X1 port map( A => n113817, Z => n120740);
   U84213 : BUF_X1 port map( A => n113815, Z => n120743);
   U84214 : BUF_X1 port map( A => n113813, Z => n120746);
   U84215 : BUF_X1 port map( A => n113811, Z => n120749);
   U84216 : BUF_X1 port map( A => n113809, Z => n120752);
   U84217 : BUF_X1 port map( A => n113807, Z => n120755);
   U84218 : BUF_X1 port map( A => n113805, Z => n120758);
   U84219 : BUF_X1 port map( A => n113803, Z => n120761);
   U84220 : BUF_X1 port map( A => n113801, Z => n120764);
   U84221 : BUF_X1 port map( A => n113799, Z => n120767);
   U84222 : BUF_X1 port map( A => n113797, Z => n120770);
   U84223 : BUF_X1 port map( A => n113795, Z => n120773);
   U84224 : BUF_X1 port map( A => n113793, Z => n120776);
   U84225 : BUF_X1 port map( A => n113791, Z => n120779);
   U84226 : BUF_X1 port map( A => n113789, Z => n120782);
   U84227 : BUF_X1 port map( A => n113787, Z => n120785);
   U84228 : BUF_X1 port map( A => n113785, Z => n120788);
   U84229 : BUF_X1 port map( A => n113783, Z => n120791);
   U84230 : BUF_X1 port map( A => n113781, Z => n120794);
   U84231 : BUF_X1 port map( A => n113779, Z => n120797);
   U84232 : BUF_X1 port map( A => n113777, Z => n120800);
   U84233 : BUF_X1 port map( A => n113775, Z => n120803);
   U84234 : BUF_X1 port map( A => n113773, Z => n120806);
   U84235 : NAND2_X1 port map( A1 => n116458, A2 => n116457, ZN => n114672);
   U84236 : OAI22_X1 port map( A1 => n120833, A2 => n113866, B1 => n120822, B2 
                           => n120665, ZN => n7435);
   U84237 : OAI22_X1 port map( A1 => n120833, A2 => n113864, B1 => n120822, B2 
                           => n120668, ZN => n7436);
   U84238 : OAI22_X1 port map( A1 => n120832, A2 => n113862, B1 => n120822, B2 
                           => n120671, ZN => n7437);
   U84239 : OAI22_X1 port map( A1 => n120832, A2 => n113860, B1 => n120822, B2 
                           => n120674, ZN => n7438);
   U84240 : OAI22_X1 port map( A1 => n120832, A2 => n113858, B1 => n120822, B2 
                           => n120677, ZN => n7439);
   U84241 : OAI22_X1 port map( A1 => n120832, A2 => n113856, B1 => n120822, B2 
                           => n120680, ZN => n7440);
   U84242 : OAI22_X1 port map( A1 => n120832, A2 => n113854, B1 => n120822, B2 
                           => n120683, ZN => n7441);
   U84243 : OAI22_X1 port map( A1 => n120832, A2 => n113852, B1 => n120822, B2 
                           => n120686, ZN => n7442);
   U84244 : OAI22_X1 port map( A1 => n120832, A2 => n113850, B1 => n120822, B2 
                           => n120689, ZN => n7443);
   U84245 : OAI22_X1 port map( A1 => n120832, A2 => n113848, B1 => n120822, B2 
                           => n120692, ZN => n7444);
   U84246 : OAI22_X1 port map( A1 => n120832, A2 => n113846, B1 => n120822, B2 
                           => n120695, ZN => n7445);
   U84247 : OAI22_X1 port map( A1 => n120832, A2 => n113844, B1 => n120822, B2 
                           => n120698, ZN => n7446);
   U84248 : OAI22_X1 port map( A1 => n120832, A2 => n113842, B1 => n120823, B2 
                           => n120701, ZN => n7447);
   U84249 : OAI22_X1 port map( A1 => n120832, A2 => n113840, B1 => n120823, B2 
                           => n120704, ZN => n7448);
   U84250 : OAI22_X1 port map( A1 => n120832, A2 => n113838, B1 => n120823, B2 
                           => n120707, ZN => n7449);
   U84251 : OAI22_X1 port map( A1 => n120831, A2 => n113836, B1 => n120823, B2 
                           => n120710, ZN => n7450);
   U84252 : OAI22_X1 port map( A1 => n120831, A2 => n113834, B1 => n120823, B2 
                           => n120713, ZN => n7451);
   U84253 : OAI22_X1 port map( A1 => n120831, A2 => n113832, B1 => n120823, B2 
                           => n120716, ZN => n7452);
   U84254 : OAI22_X1 port map( A1 => n120831, A2 => n113830, B1 => n120823, B2 
                           => n120719, ZN => n7453);
   U84255 : OAI22_X1 port map( A1 => n120831, A2 => n113828, B1 => n120823, B2 
                           => n120722, ZN => n7454);
   U84256 : OAI22_X1 port map( A1 => n120831, A2 => n113826, B1 => n120823, B2 
                           => n120725, ZN => n7455);
   U84257 : OAI22_X1 port map( A1 => n120831, A2 => n113824, B1 => n120823, B2 
                           => n120728, ZN => n7456);
   U84258 : OAI22_X1 port map( A1 => n120831, A2 => n113822, B1 => n120823, B2 
                           => n120731, ZN => n7457);
   U84259 : OAI22_X1 port map( A1 => n120831, A2 => n113820, B1 => n120823, B2 
                           => n120734, ZN => n7458);
   U84260 : OAI22_X1 port map( A1 => n120831, A2 => n113818, B1 => n120824, B2 
                           => n120737, ZN => n7459);
   U84261 : OAI22_X1 port map( A1 => n120831, A2 => n113816, B1 => n120824, B2 
                           => n120740, ZN => n7460);
   U84262 : OAI22_X1 port map( A1 => n120831, A2 => n113814, B1 => n120824, B2 
                           => n120743, ZN => n7461);
   U84263 : OAI22_X1 port map( A1 => n120830, A2 => n113812, B1 => n120824, B2 
                           => n120746, ZN => n7462);
   U84264 : OAI22_X1 port map( A1 => n120830, A2 => n113810, B1 => n120824, B2 
                           => n120749, ZN => n7463);
   U84265 : OAI22_X1 port map( A1 => n120830, A2 => n113808, B1 => n120824, B2 
                           => n120752, ZN => n7464);
   U84266 : OAI22_X1 port map( A1 => n120830, A2 => n113806, B1 => n120824, B2 
                           => n120755, ZN => n7465);
   U84267 : OAI22_X1 port map( A1 => n120830, A2 => n113804, B1 => n120824, B2 
                           => n120758, ZN => n7466);
   U84268 : OAI22_X1 port map( A1 => n120830, A2 => n113802, B1 => n120824, B2 
                           => n120761, ZN => n7467);
   U84269 : OAI22_X1 port map( A1 => n120830, A2 => n113800, B1 => n120824, B2 
                           => n120764, ZN => n7468);
   U84270 : OAI22_X1 port map( A1 => n120830, A2 => n113798, B1 => n120824, B2 
                           => n120767, ZN => n7469);
   U84271 : OAI22_X1 port map( A1 => n120831, A2 => n113796, B1 => n120824, B2 
                           => n120770, ZN => n7470);
   U84272 : OAI22_X1 port map( A1 => n120830, A2 => n113794, B1 => n120825, B2 
                           => n120773, ZN => n7471);
   U84273 : OAI22_X1 port map( A1 => n120830, A2 => n113792, B1 => n120825, B2 
                           => n120776, ZN => n7472);
   U84274 : OAI22_X1 port map( A1 => n120830, A2 => n113790, B1 => n120825, B2 
                           => n120779, ZN => n7473);
   U84275 : OAI22_X1 port map( A1 => n120830, A2 => n113788, B1 => n120825, B2 
                           => n120782, ZN => n7474);
   U84276 : OAI22_X1 port map( A1 => n120830, A2 => n113786, B1 => n120825, B2 
                           => n120785, ZN => n7475);
   U84277 : OAI22_X1 port map( A1 => n120829, A2 => n113784, B1 => n120825, B2 
                           => n120788, ZN => n7476);
   U84278 : OAI22_X1 port map( A1 => n120829, A2 => n113782, B1 => n120825, B2 
                           => n120791, ZN => n7477);
   U84279 : OAI22_X1 port map( A1 => n120829, A2 => n113780, B1 => n120825, B2 
                           => n120794, ZN => n7478);
   U84280 : OAI22_X1 port map( A1 => n120829, A2 => n113778, B1 => n120825, B2 
                           => n120797, ZN => n7479);
   U84281 : OAI22_X1 port map( A1 => n120829, A2 => n113776, B1 => n120825, B2 
                           => n120800, ZN => n7480);
   U84282 : OAI22_X1 port map( A1 => n120829, A2 => n113774, B1 => n120825, B2 
                           => n120803, ZN => n7481);
   U84283 : OAI22_X1 port map( A1 => n120829, A2 => n113772, B1 => n120825, B2 
                           => n120806, ZN => n7482);
   U84284 : NAND2_X1 port map( A1 => n117949, A2 => n117945, ZN => n116487);
   U84285 : NAND2_X1 port map( A1 => n117949, A2 => n117953, ZN => n116492);
   U84286 : NAND2_X1 port map( A1 => n117955, A2 => n117953, ZN => n116499);
   U84287 : NAND2_X1 port map( A1 => n117961, A2 => n117953, ZN => n116504);
   U84288 : OAI22_X1 port map( A1 => n120511, A2 => n114127, B1 => n120809, B2 
                           => n120505, ZN => n6843);
   U84289 : OAI22_X1 port map( A1 => n120511, A2 => n114126, B1 => n120812, B2 
                           => n120505, ZN => n6844);
   U84290 : OAI22_X1 port map( A1 => n120511, A2 => n114125, B1 => n120815, B2 
                           => n120505, ZN => n6845);
   U84291 : OAI22_X1 port map( A1 => n120511, A2 => n114123, B1 => n120818, B2 
                           => n120505, ZN => n6846);
   U84292 : OAI22_X1 port map( A1 => n120561, A2 => n113985, B1 => n120809, B2 
                           => n120555, ZN => n7099);
   U84293 : OAI22_X1 port map( A1 => n120561, A2 => n113984, B1 => n120812, B2 
                           => n120555, ZN => n7100);
   U84294 : OAI22_X1 port map( A1 => n120561, A2 => n113983, B1 => n120815, B2 
                           => n120555, ZN => n7101);
   U84295 : OAI22_X1 port map( A1 => n120561, A2 => n113981, B1 => n120818, B2 
                           => n120555, ZN => n7102);
   U84296 : OAI22_X1 port map( A1 => n120610, A2 => n113907, B1 => n120809, B2 
                           => n120604, ZN => n7355);
   U84297 : OAI22_X1 port map( A1 => n120610, A2 => n113906, B1 => n120812, B2 
                           => n120604, ZN => n7356);
   U84298 : OAI22_X1 port map( A1 => n120610, A2 => n113905, B1 => n120815, B2 
                           => n120604, ZN => n7357);
   U84299 : OAI22_X1 port map( A1 => n120610, A2 => n113903, B1 => n120818, B2 
                           => n120604, ZN => n7358);
   U84300 : NAND2_X1 port map( A1 => n116446, A2 => n116457, ZN => n114690);
   U84301 : OAI22_X1 port map( A1 => n120252, A2 => n114756, B1 => n120811, B2 
                           => n120245, ZN => n5496);
   U84302 : OAI22_X1 port map( A1 => n120252, A2 => n114730, B1 => n120814, B2 
                           => n120245, ZN => n5498);
   U84303 : OAI22_X1 port map( A1 => n120252, A2 => n114704, B1 => n120817, B2 
                           => n120245, ZN => n5500);
   U84304 : OAI22_X1 port map( A1 => n120252, A2 => n114644, B1 => n120820, B2 
                           => n120245, ZN => n5502);
   U84305 : OAI22_X1 port map( A1 => n120574, A2 => n113919, B1 => n120809, B2 
                           => n120567, ZN => n7163);
   U84306 : OAI22_X1 port map( A1 => n120574, A2 => n113918, B1 => n120812, B2 
                           => n120567, ZN => n7164);
   U84307 : OAI22_X1 port map( A1 => n120574, A2 => n113917, B1 => n120815, B2 
                           => n120567, ZN => n7165);
   U84308 : OAI22_X1 port map( A1 => n120574, A2 => n113915, B1 => n120818, B2 
                           => n120567, ZN => n7166);
   U84309 : OAI22_X1 port map( A1 => n120378, A2 => n114239, B1 => n120810, B2 
                           => n120371, ZN => n6139);
   U84310 : OAI22_X1 port map( A1 => n120378, A2 => n114238, B1 => n120813, B2 
                           => n120371, ZN => n6140);
   U84311 : OAI22_X1 port map( A1 => n120378, A2 => n114237, B1 => n120816, B2 
                           => n120371, ZN => n6141);
   U84312 : OAI22_X1 port map( A1 => n120378, A2 => n114235, B1 => n120819, B2 
                           => n120371, ZN => n6142);
   U84313 : OAI22_X1 port map( A1 => n120290, A2 => n114514, B1 => n120811, B2 
                           => n120283, ZN => n5691);
   U84314 : OAI22_X1 port map( A1 => n120290, A2 => n114513, B1 => n120814, B2 
                           => n120283, ZN => n5692);
   U84315 : OAI22_X1 port map( A1 => n120290, A2 => n114512, B1 => n120817, B2 
                           => n120283, ZN => n5693);
   U84316 : OAI22_X1 port map( A1 => n120290, A2 => n114510, B1 => n120820, B2 
                           => n120283, ZN => n5694);
   U84317 : OAI22_X1 port map( A1 => n120265, A2 => n114582, B1 => n120811, B2 
                           => n120258, ZN => n5563);
   U84318 : OAI22_X1 port map( A1 => n120265, A2 => n114581, B1 => n120814, B2 
                           => n120258, ZN => n5564);
   U84319 : OAI22_X1 port map( A1 => n120265, A2 => n114580, B1 => n120817, B2 
                           => n120258, ZN => n5565);
   U84320 : OAI22_X1 port map( A1 => n120265, A2 => n114578, B1 => n120820, B2 
                           => n120258, ZN => n5566);
   U84321 : OAI22_X1 port map( A1 => n120415, A2 => n114150, B1 => n120810, B2 
                           => n120408, ZN => n6331);
   U84322 : OAI22_X1 port map( A1 => n120415, A2 => n114149, B1 => n120813, B2 
                           => n120408, ZN => n6332);
   U84323 : OAI22_X1 port map( A1 => n120415, A2 => n114148, B1 => n120816, B2 
                           => n120408, ZN => n6333);
   U84324 : OAI22_X1 port map( A1 => n120415, A2 => n114146, B1 => n120819, B2 
                           => n120408, ZN => n6334);
   U84325 : OAI22_X1 port map( A1 => n120316, A2 => n114382, B1 => n120811, B2 
                           => n120309, ZN => n5819);
   U84326 : OAI22_X1 port map( A1 => n120316, A2 => n114381, B1 => n120814, B2 
                           => n120309, ZN => n5820);
   U84327 : OAI22_X1 port map( A1 => n120316, A2 => n114380, B1 => n120817, B2 
                           => n120309, ZN => n5821);
   U84328 : OAI22_X1 port map( A1 => n120316, A2 => n114378, B1 => n120820, B2 
                           => n120309, ZN => n5822);
   U84329 : OAI22_X1 port map( A1 => n120303, A2 => n114448, B1 => n120811, B2 
                           => n120296, ZN => n5755);
   U84330 : OAI22_X1 port map( A1 => n120303, A2 => n114447, B1 => n120814, B2 
                           => n120296, ZN => n5756);
   U84331 : OAI22_X1 port map( A1 => n120303, A2 => n114446, B1 => n120817, B2 
                           => n120296, ZN => n5757);
   U84332 : OAI22_X1 port map( A1 => n120303, A2 => n114444, B1 => n120820, B2 
                           => n120296, ZN => n5758);
   U84333 : NAND2_X1 port map( A1 => n116448, A2 => n116447, ZN => n114654);
   U84334 : OAI22_X1 port map( A1 => n120248, A2 => n116434, B1 => n120631, B2 
                           => n120240, ZN => n5376);
   U84335 : OAI22_X1 port map( A1 => n120248, A2 => n116406, B1 => n120634, B2 
                           => n120240, ZN => n5378);
   U84336 : OAI22_X1 port map( A1 => n120248, A2 => n116378, B1 => n120637, B2 
                           => n120240, ZN => n5380);
   U84337 : OAI22_X1 port map( A1 => n120248, A2 => n116350, B1 => n120640, B2 
                           => n120240, ZN => n5382);
   U84338 : OAI22_X1 port map( A1 => n120248, A2 => n116322, B1 => n120643, B2 
                           => n120240, ZN => n5384);
   U84339 : OAI22_X1 port map( A1 => n120248, A2 => n116294, B1 => n120646, B2 
                           => n120240, ZN => n5386);
   U84340 : OAI22_X1 port map( A1 => n120248, A2 => n116266, B1 => n120649, B2 
                           => n120240, ZN => n5388);
   U84341 : OAI22_X1 port map( A1 => n120248, A2 => n116238, B1 => n120652, B2 
                           => n120240, ZN => n5390);
   U84342 : OAI22_X1 port map( A1 => n120248, A2 => n116210, B1 => n120655, B2 
                           => n120240, ZN => n5392);
   U84343 : OAI22_X1 port map( A1 => n120248, A2 => n116182, B1 => n120658, B2 
                           => n120240, ZN => n5394);
   U84344 : OAI22_X1 port map( A1 => n120248, A2 => n116154, B1 => n120661, B2 
                           => n120240, ZN => n5396);
   U84345 : OAI22_X1 port map( A1 => n120248, A2 => n116126, B1 => n120664, B2 
                           => n120240, ZN => n5398);
   U84346 : OAI22_X1 port map( A1 => n120249, A2 => n116098, B1 => n120667, B2 
                           => n120241, ZN => n5400);
   U84347 : OAI22_X1 port map( A1 => n120249, A2 => n116070, B1 => n120670, B2 
                           => n120241, ZN => n5402);
   U84348 : OAI22_X1 port map( A1 => n120249, A2 => n116042, B1 => n120673, B2 
                           => n120241, ZN => n5404);
   U84349 : OAI22_X1 port map( A1 => n120249, A2 => n116014, B1 => n120676, B2 
                           => n120241, ZN => n5406);
   U84350 : OAI22_X1 port map( A1 => n120249, A2 => n115986, B1 => n120679, B2 
                           => n120241, ZN => n5408);
   U84351 : OAI22_X1 port map( A1 => n120249, A2 => n115958, B1 => n120682, B2 
                           => n120241, ZN => n5410);
   U84352 : OAI22_X1 port map( A1 => n120249, A2 => n115930, B1 => n120685, B2 
                           => n120241, ZN => n5412);
   U84353 : OAI22_X1 port map( A1 => n120249, A2 => n115902, B1 => n120688, B2 
                           => n120241, ZN => n5414);
   U84354 : OAI22_X1 port map( A1 => n120249, A2 => n115874, B1 => n120691, B2 
                           => n120241, ZN => n5416);
   U84355 : OAI22_X1 port map( A1 => n120249, A2 => n115846, B1 => n120694, B2 
                           => n120241, ZN => n5418);
   U84356 : OAI22_X1 port map( A1 => n120249, A2 => n115818, B1 => n120697, B2 
                           => n120241, ZN => n5420);
   U84357 : OAI22_X1 port map( A1 => n120249, A2 => n115790, B1 => n120700, B2 
                           => n120241, ZN => n5422);
   U84358 : OAI22_X1 port map( A1 => n120249, A2 => n115762, B1 => n120703, B2 
                           => n120242, ZN => n5424);
   U84359 : OAI22_X1 port map( A1 => n120250, A2 => n115734, B1 => n120706, B2 
                           => n120242, ZN => n5426);
   U84360 : OAI22_X1 port map( A1 => n120250, A2 => n115706, B1 => n120709, B2 
                           => n120242, ZN => n5428);
   U84361 : OAI22_X1 port map( A1 => n120250, A2 => n115678, B1 => n120712, B2 
                           => n120242, ZN => n5430);
   U84362 : OAI22_X1 port map( A1 => n120250, A2 => n115650, B1 => n120715, B2 
                           => n120242, ZN => n5432);
   U84363 : OAI22_X1 port map( A1 => n120250, A2 => n115622, B1 => n120718, B2 
                           => n120242, ZN => n5434);
   U84364 : OAI22_X1 port map( A1 => n120250, A2 => n115594, B1 => n120721, B2 
                           => n120242, ZN => n5436);
   U84365 : OAI22_X1 port map( A1 => n120250, A2 => n115566, B1 => n120724, B2 
                           => n120242, ZN => n5438);
   U84366 : OAI22_X1 port map( A1 => n120250, A2 => n115538, B1 => n120727, B2 
                           => n120242, ZN => n5440);
   U84367 : OAI22_X1 port map( A1 => n120250, A2 => n115510, B1 => n120730, B2 
                           => n120242, ZN => n5442);
   U84368 : OAI22_X1 port map( A1 => n120250, A2 => n115482, B1 => n120733, B2 
                           => n120242, ZN => n5444);
   U84369 : OAI22_X1 port map( A1 => n120250, A2 => n115454, B1 => n120736, B2 
                           => n120242, ZN => n5446);
   U84370 : OAI22_X1 port map( A1 => n120250, A2 => n115426, B1 => n120739, B2 
                           => n120243, ZN => n5448);
   U84371 : OAI22_X1 port map( A1 => n120250, A2 => n115398, B1 => n120742, B2 
                           => n120243, ZN => n5450);
   U84372 : OAI22_X1 port map( A1 => n120251, A2 => n115370, B1 => n120745, B2 
                           => n120243, ZN => n5452);
   U84373 : OAI22_X1 port map( A1 => n120251, A2 => n115342, B1 => n120748, B2 
                           => n120243, ZN => n5454);
   U84374 : OAI22_X1 port map( A1 => n120251, A2 => n115314, B1 => n120751, B2 
                           => n120243, ZN => n5456);
   U84375 : OAI22_X1 port map( A1 => n120251, A2 => n115286, B1 => n120754, B2 
                           => n120243, ZN => n5458);
   U84376 : OAI22_X1 port map( A1 => n120251, A2 => n115258, B1 => n120757, B2 
                           => n120243, ZN => n5460);
   U84377 : OAI22_X1 port map( A1 => n120251, A2 => n115230, B1 => n120760, B2 
                           => n120243, ZN => n5462);
   U84378 : OAI22_X1 port map( A1 => n120251, A2 => n115202, B1 => n120763, B2 
                           => n120243, ZN => n5464);
   U84379 : OAI22_X1 port map( A1 => n120251, A2 => n115174, B1 => n120766, B2 
                           => n120243, ZN => n5466);
   U84380 : OAI22_X1 port map( A1 => n120251, A2 => n115146, B1 => n120769, B2 
                           => n120243, ZN => n5468);
   U84381 : OAI22_X1 port map( A1 => n120251, A2 => n115118, B1 => n120772, B2 
                           => n120243, ZN => n5470);
   U84382 : OAI22_X1 port map( A1 => n120251, A2 => n115090, B1 => n120775, B2 
                           => n120244, ZN => n5472);
   U84383 : OAI22_X1 port map( A1 => n120251, A2 => n115062, B1 => n120778, B2 
                           => n120244, ZN => n5474);
   U84384 : OAI22_X1 port map( A1 => n120251, A2 => n115034, B1 => n120781, B2 
                           => n120244, ZN => n5476);
   U84385 : OAI22_X1 port map( A1 => n120252, A2 => n115006, B1 => n120784, B2 
                           => n120244, ZN => n5478);
   U84386 : OAI22_X1 port map( A1 => n120252, A2 => n114978, B1 => n120787, B2 
                           => n120244, ZN => n5480);
   U84387 : OAI22_X1 port map( A1 => n120252, A2 => n114950, B1 => n120790, B2 
                           => n120244, ZN => n5482);
   U84388 : OAI22_X1 port map( A1 => n120252, A2 => n114922, B1 => n120793, B2 
                           => n120244, ZN => n5484);
   U84389 : OAI22_X1 port map( A1 => n120252, A2 => n114894, B1 => n120796, B2 
                           => n120244, ZN => n5486);
   U84390 : OAI22_X1 port map( A1 => n120252, A2 => n114866, B1 => n120799, B2 
                           => n120244, ZN => n5488);
   U84391 : OAI22_X1 port map( A1 => n120252, A2 => n114838, B1 => n120802, B2 
                           => n120244, ZN => n5490);
   U84392 : OAI22_X1 port map( A1 => n120252, A2 => n114810, B1 => n120805, B2 
                           => n120244, ZN => n5492);
   U84393 : OAI22_X1 port map( A1 => n120252, A2 => n114782, B1 => n120808, B2 
                           => n120244, ZN => n5494);
   U84394 : OAI22_X1 port map( A1 => n120261, A2 => n114642, B1 => n120631, B2 
                           => n120253, ZN => n5503);
   U84395 : OAI22_X1 port map( A1 => n120261, A2 => n114641, B1 => n120634, B2 
                           => n120253, ZN => n5504);
   U84396 : OAI22_X1 port map( A1 => n120261, A2 => n114640, B1 => n120637, B2 
                           => n120253, ZN => n5505);
   U84397 : OAI22_X1 port map( A1 => n120261, A2 => n114639, B1 => n120640, B2 
                           => n120253, ZN => n5506);
   U84398 : OAI22_X1 port map( A1 => n120261, A2 => n114638, B1 => n120643, B2 
                           => n120253, ZN => n5507);
   U84399 : OAI22_X1 port map( A1 => n120261, A2 => n114637, B1 => n120646, B2 
                           => n120253, ZN => n5508);
   U84400 : OAI22_X1 port map( A1 => n120261, A2 => n114636, B1 => n120649, B2 
                           => n120253, ZN => n5509);
   U84401 : OAI22_X1 port map( A1 => n120261, A2 => n114635, B1 => n120652, B2 
                           => n120253, ZN => n5510);
   U84402 : OAI22_X1 port map( A1 => n120261, A2 => n114634, B1 => n120655, B2 
                           => n120253, ZN => n5511);
   U84403 : OAI22_X1 port map( A1 => n120261, A2 => n114633, B1 => n120658, B2 
                           => n120253, ZN => n5512);
   U84404 : OAI22_X1 port map( A1 => n120261, A2 => n114632, B1 => n120661, B2 
                           => n120253, ZN => n5513);
   U84405 : OAI22_X1 port map( A1 => n120261, A2 => n114631, B1 => n120664, B2 
                           => n120253, ZN => n5514);
   U84406 : OAI22_X1 port map( A1 => n120262, A2 => n114630, B1 => n120667, B2 
                           => n120254, ZN => n5515);
   U84407 : OAI22_X1 port map( A1 => n120262, A2 => n114629, B1 => n120670, B2 
                           => n120254, ZN => n5516);
   U84408 : OAI22_X1 port map( A1 => n120262, A2 => n114628, B1 => n120673, B2 
                           => n120254, ZN => n5517);
   U84409 : OAI22_X1 port map( A1 => n120262, A2 => n114627, B1 => n120676, B2 
                           => n120254, ZN => n5518);
   U84410 : OAI22_X1 port map( A1 => n120262, A2 => n114626, B1 => n120679, B2 
                           => n120254, ZN => n5519);
   U84411 : OAI22_X1 port map( A1 => n120262, A2 => n114625, B1 => n120682, B2 
                           => n120254, ZN => n5520);
   U84412 : OAI22_X1 port map( A1 => n120262, A2 => n114624, B1 => n120685, B2 
                           => n120254, ZN => n5521);
   U84413 : OAI22_X1 port map( A1 => n120262, A2 => n114623, B1 => n120688, B2 
                           => n120254, ZN => n5522);
   U84414 : OAI22_X1 port map( A1 => n120262, A2 => n114622, B1 => n120691, B2 
                           => n120254, ZN => n5523);
   U84415 : OAI22_X1 port map( A1 => n120262, A2 => n114621, B1 => n120694, B2 
                           => n120254, ZN => n5524);
   U84416 : OAI22_X1 port map( A1 => n120262, A2 => n114620, B1 => n120697, B2 
                           => n120254, ZN => n5525);
   U84417 : OAI22_X1 port map( A1 => n120262, A2 => n114619, B1 => n120700, B2 
                           => n120254, ZN => n5526);
   U84418 : OAI22_X1 port map( A1 => n120262, A2 => n114618, B1 => n120703, B2 
                           => n120255, ZN => n5527);
   U84419 : OAI22_X1 port map( A1 => n120263, A2 => n114617, B1 => n120706, B2 
                           => n120255, ZN => n5528);
   U84420 : OAI22_X1 port map( A1 => n120263, A2 => n114616, B1 => n120709, B2 
                           => n120255, ZN => n5529);
   U84421 : OAI22_X1 port map( A1 => n120263, A2 => n114615, B1 => n120712, B2 
                           => n120255, ZN => n5530);
   U84422 : OAI22_X1 port map( A1 => n120263, A2 => n114614, B1 => n120715, B2 
                           => n120255, ZN => n5531);
   U84423 : OAI22_X1 port map( A1 => n120263, A2 => n114613, B1 => n120718, B2 
                           => n120255, ZN => n5532);
   U84424 : OAI22_X1 port map( A1 => n120263, A2 => n114612, B1 => n120721, B2 
                           => n120255, ZN => n5533);
   U84425 : OAI22_X1 port map( A1 => n120263, A2 => n114611, B1 => n120724, B2 
                           => n120255, ZN => n5534);
   U84426 : OAI22_X1 port map( A1 => n120263, A2 => n114610, B1 => n120727, B2 
                           => n120255, ZN => n5535);
   U84427 : OAI22_X1 port map( A1 => n120263, A2 => n114609, B1 => n120730, B2 
                           => n120255, ZN => n5536);
   U84428 : OAI22_X1 port map( A1 => n120263, A2 => n114608, B1 => n120733, B2 
                           => n120255, ZN => n5537);
   U84429 : OAI22_X1 port map( A1 => n120263, A2 => n114607, B1 => n120736, B2 
                           => n120255, ZN => n5538);
   U84430 : OAI22_X1 port map( A1 => n120263, A2 => n114606, B1 => n120739, B2 
                           => n120256, ZN => n5539);
   U84431 : OAI22_X1 port map( A1 => n120263, A2 => n114605, B1 => n120742, B2 
                           => n120256, ZN => n5540);
   U84432 : OAI22_X1 port map( A1 => n120264, A2 => n114604, B1 => n120745, B2 
                           => n120256, ZN => n5541);
   U84433 : OAI22_X1 port map( A1 => n120264, A2 => n114603, B1 => n120748, B2 
                           => n120256, ZN => n5542);
   U84434 : OAI22_X1 port map( A1 => n120264, A2 => n114602, B1 => n120751, B2 
                           => n120256, ZN => n5543);
   U84435 : OAI22_X1 port map( A1 => n120264, A2 => n114601, B1 => n120754, B2 
                           => n120256, ZN => n5544);
   U84436 : OAI22_X1 port map( A1 => n120264, A2 => n114600, B1 => n120757, B2 
                           => n120256, ZN => n5545);
   U84437 : OAI22_X1 port map( A1 => n120264, A2 => n114599, B1 => n120760, B2 
                           => n120256, ZN => n5546);
   U84438 : OAI22_X1 port map( A1 => n120264, A2 => n114598, B1 => n120763, B2 
                           => n120256, ZN => n5547);
   U84439 : OAI22_X1 port map( A1 => n120286, A2 => n114574, B1 => n120631, B2 
                           => n120278, ZN => n5631);
   U84440 : OAI22_X1 port map( A1 => n120286, A2 => n114573, B1 => n120634, B2 
                           => n120278, ZN => n5632);
   U84441 : OAI22_X1 port map( A1 => n120286, A2 => n114572, B1 => n120637, B2 
                           => n120278, ZN => n5633);
   U84442 : OAI22_X1 port map( A1 => n120286, A2 => n114571, B1 => n120640, B2 
                           => n120278, ZN => n5634);
   U84443 : OAI22_X1 port map( A1 => n120286, A2 => n114570, B1 => n120643, B2 
                           => n120278, ZN => n5635);
   U84444 : OAI22_X1 port map( A1 => n120286, A2 => n114569, B1 => n120646, B2 
                           => n120278, ZN => n5636);
   U84445 : OAI22_X1 port map( A1 => n120286, A2 => n114568, B1 => n120649, B2 
                           => n120278, ZN => n5637);
   U84446 : OAI22_X1 port map( A1 => n120286, A2 => n114567, B1 => n120652, B2 
                           => n120278, ZN => n5638);
   U84447 : OAI22_X1 port map( A1 => n120286, A2 => n114566, B1 => n120655, B2 
                           => n120278, ZN => n5639);
   U84448 : OAI22_X1 port map( A1 => n120286, A2 => n114565, B1 => n120658, B2 
                           => n120278, ZN => n5640);
   U84449 : OAI22_X1 port map( A1 => n120286, A2 => n114564, B1 => n120661, B2 
                           => n120278, ZN => n5641);
   U84450 : OAI22_X1 port map( A1 => n120286, A2 => n114563, B1 => n120664, B2 
                           => n120278, ZN => n5642);
   U84451 : OAI22_X1 port map( A1 => n120287, A2 => n114562, B1 => n120667, B2 
                           => n120279, ZN => n5643);
   U84452 : OAI22_X1 port map( A1 => n120287, A2 => n114561, B1 => n120670, B2 
                           => n120279, ZN => n5644);
   U84453 : OAI22_X1 port map( A1 => n120287, A2 => n114560, B1 => n120673, B2 
                           => n120279, ZN => n5645);
   U84454 : OAI22_X1 port map( A1 => n120287, A2 => n114559, B1 => n120676, B2 
                           => n120279, ZN => n5646);
   U84455 : OAI22_X1 port map( A1 => n120287, A2 => n114558, B1 => n120679, B2 
                           => n120279, ZN => n5647);
   U84456 : OAI22_X1 port map( A1 => n120287, A2 => n114557, B1 => n120682, B2 
                           => n120279, ZN => n5648);
   U84457 : OAI22_X1 port map( A1 => n120287, A2 => n114556, B1 => n120685, B2 
                           => n120279, ZN => n5649);
   U84458 : OAI22_X1 port map( A1 => n120287, A2 => n114555, B1 => n120688, B2 
                           => n120279, ZN => n5650);
   U84459 : OAI22_X1 port map( A1 => n120287, A2 => n114554, B1 => n120691, B2 
                           => n120279, ZN => n5651);
   U84460 : OAI22_X1 port map( A1 => n120287, A2 => n114553, B1 => n120694, B2 
                           => n120279, ZN => n5652);
   U84461 : OAI22_X1 port map( A1 => n120287, A2 => n114552, B1 => n120697, B2 
                           => n120279, ZN => n5653);
   U84462 : OAI22_X1 port map( A1 => n120287, A2 => n114551, B1 => n120700, B2 
                           => n120279, ZN => n5654);
   U84463 : OAI22_X1 port map( A1 => n120287, A2 => n114550, B1 => n120703, B2 
                           => n120280, ZN => n5655);
   U84464 : OAI22_X1 port map( A1 => n120288, A2 => n114549, B1 => n120706, B2 
                           => n120280, ZN => n5656);
   U84465 : OAI22_X1 port map( A1 => n120288, A2 => n114548, B1 => n120709, B2 
                           => n120280, ZN => n5657);
   U84466 : OAI22_X1 port map( A1 => n120288, A2 => n114547, B1 => n120712, B2 
                           => n120280, ZN => n5658);
   U84467 : OAI22_X1 port map( A1 => n120288, A2 => n114546, B1 => n120715, B2 
                           => n120280, ZN => n5659);
   U84468 : OAI22_X1 port map( A1 => n120288, A2 => n114545, B1 => n120718, B2 
                           => n120280, ZN => n5660);
   U84469 : OAI22_X1 port map( A1 => n120288, A2 => n114544, B1 => n120721, B2 
                           => n120280, ZN => n5661);
   U84470 : OAI22_X1 port map( A1 => n120288, A2 => n114543, B1 => n120724, B2 
                           => n120280, ZN => n5662);
   U84471 : OAI22_X1 port map( A1 => n120288, A2 => n114542, B1 => n120727, B2 
                           => n120280, ZN => n5663);
   U84472 : OAI22_X1 port map( A1 => n120288, A2 => n114541, B1 => n120730, B2 
                           => n120280, ZN => n5664);
   U84473 : OAI22_X1 port map( A1 => n120288, A2 => n114540, B1 => n120733, B2 
                           => n120280, ZN => n5665);
   U84474 : OAI22_X1 port map( A1 => n120288, A2 => n114539, B1 => n120736, B2 
                           => n120280, ZN => n5666);
   U84475 : OAI22_X1 port map( A1 => n120288, A2 => n114538, B1 => n120739, B2 
                           => n120281, ZN => n5667);
   U84476 : OAI22_X1 port map( A1 => n120288, A2 => n114537, B1 => n120742, B2 
                           => n120281, ZN => n5668);
   U84477 : OAI22_X1 port map( A1 => n120289, A2 => n114536, B1 => n120745, B2 
                           => n120281, ZN => n5669);
   U84478 : OAI22_X1 port map( A1 => n120289, A2 => n114535, B1 => n120748, B2 
                           => n120281, ZN => n5670);
   U84479 : OAI22_X1 port map( A1 => n120289, A2 => n114534, B1 => n120751, B2 
                           => n120281, ZN => n5671);
   U84480 : OAI22_X1 port map( A1 => n120289, A2 => n114533, B1 => n120754, B2 
                           => n120281, ZN => n5672);
   U84481 : OAI22_X1 port map( A1 => n120289, A2 => n114532, B1 => n120757, B2 
                           => n120281, ZN => n5673);
   U84482 : OAI22_X1 port map( A1 => n120289, A2 => n114531, B1 => n120760, B2 
                           => n120281, ZN => n5674);
   U84483 : OAI22_X1 port map( A1 => n120289, A2 => n114530, B1 => n120763, B2 
                           => n120281, ZN => n5675);
   U84484 : OAI22_X1 port map( A1 => n120289, A2 => n114529, B1 => n120766, B2 
                           => n120281, ZN => n5676);
   U84485 : OAI22_X1 port map( A1 => n120289, A2 => n114528, B1 => n120769, B2 
                           => n120281, ZN => n5677);
   U84486 : OAI22_X1 port map( A1 => n120289, A2 => n114527, B1 => n120772, B2 
                           => n120281, ZN => n5678);
   U84487 : OAI22_X1 port map( A1 => n120289, A2 => n114526, B1 => n120775, B2 
                           => n120282, ZN => n5679);
   U84488 : OAI22_X1 port map( A1 => n120289, A2 => n114525, B1 => n120778, B2 
                           => n120282, ZN => n5680);
   U84489 : OAI22_X1 port map( A1 => n120289, A2 => n114524, B1 => n120781, B2 
                           => n120282, ZN => n5681);
   U84490 : OAI22_X1 port map( A1 => n120290, A2 => n114523, B1 => n120784, B2 
                           => n120282, ZN => n5682);
   U84491 : OAI22_X1 port map( A1 => n120290, A2 => n114522, B1 => n120787, B2 
                           => n120282, ZN => n5683);
   U84492 : OAI22_X1 port map( A1 => n120290, A2 => n114521, B1 => n120790, B2 
                           => n120282, ZN => n5684);
   U84493 : OAI22_X1 port map( A1 => n120290, A2 => n114520, B1 => n120793, B2 
                           => n120282, ZN => n5685);
   U84494 : OAI22_X1 port map( A1 => n120290, A2 => n114519, B1 => n120796, B2 
                           => n120282, ZN => n5686);
   U84495 : OAI22_X1 port map( A1 => n120290, A2 => n114518, B1 => n120799, B2 
                           => n120282, ZN => n5687);
   U84496 : OAI22_X1 port map( A1 => n120290, A2 => n114517, B1 => n120802, B2 
                           => n120282, ZN => n5688);
   U84497 : OAI22_X1 port map( A1 => n120290, A2 => n114516, B1 => n120805, B2 
                           => n120282, ZN => n5689);
   U84498 : OAI22_X1 port map( A1 => n120290, A2 => n114515, B1 => n120808, B2 
                           => n120282, ZN => n5690);
   U84499 : OAI22_X1 port map( A1 => n120264, A2 => n114597, B1 => n120766, B2 
                           => n120256, ZN => n5548);
   U84500 : OAI22_X1 port map( A1 => n120264, A2 => n114596, B1 => n120769, B2 
                           => n120256, ZN => n5549);
   U84501 : OAI22_X1 port map( A1 => n120264, A2 => n114595, B1 => n120772, B2 
                           => n120256, ZN => n5550);
   U84502 : OAI22_X1 port map( A1 => n120264, A2 => n114594, B1 => n120775, B2 
                           => n120257, ZN => n5551);
   U84503 : OAI22_X1 port map( A1 => n120264, A2 => n114593, B1 => n120778, B2 
                           => n120257, ZN => n5552);
   U84504 : OAI22_X1 port map( A1 => n120264, A2 => n114592, B1 => n120781, B2 
                           => n120257, ZN => n5553);
   U84505 : OAI22_X1 port map( A1 => n120265, A2 => n114591, B1 => n120784, B2 
                           => n120257, ZN => n5554);
   U84506 : OAI22_X1 port map( A1 => n120265, A2 => n114590, B1 => n120787, B2 
                           => n120257, ZN => n5555);
   U84507 : OAI22_X1 port map( A1 => n120265, A2 => n114589, B1 => n120790, B2 
                           => n120257, ZN => n5556);
   U84508 : OAI22_X1 port map( A1 => n120265, A2 => n114588, B1 => n120793, B2 
                           => n120257, ZN => n5557);
   U84509 : OAI22_X1 port map( A1 => n120265, A2 => n114587, B1 => n120796, B2 
                           => n120257, ZN => n5558);
   U84510 : OAI22_X1 port map( A1 => n120265, A2 => n114586, B1 => n120799, B2 
                           => n120257, ZN => n5559);
   U84511 : OAI22_X1 port map( A1 => n120265, A2 => n114585, B1 => n120802, B2 
                           => n120257, ZN => n5560);
   U84512 : OAI22_X1 port map( A1 => n120265, A2 => n114584, B1 => n120805, B2 
                           => n120257, ZN => n5561);
   U84513 : OAI22_X1 port map( A1 => n120265, A2 => n114583, B1 => n120808, B2 
                           => n120257, ZN => n5562);
   U84514 : OAI22_X1 port map( A1 => n120312, A2 => n114442, B1 => n120631, B2 
                           => n120304, ZN => n5759);
   U84515 : OAI22_X1 port map( A1 => n120312, A2 => n114441, B1 => n120634, B2 
                           => n120304, ZN => n5760);
   U84516 : OAI22_X1 port map( A1 => n120312, A2 => n114440, B1 => n120637, B2 
                           => n120304, ZN => n5761);
   U84517 : OAI22_X1 port map( A1 => n120312, A2 => n114439, B1 => n120640, B2 
                           => n120304, ZN => n5762);
   U84518 : OAI22_X1 port map( A1 => n120312, A2 => n114438, B1 => n120643, B2 
                           => n120304, ZN => n5763);
   U84519 : OAI22_X1 port map( A1 => n120312, A2 => n114437, B1 => n120646, B2 
                           => n120304, ZN => n5764);
   U84520 : OAI22_X1 port map( A1 => n120312, A2 => n114436, B1 => n120649, B2 
                           => n120304, ZN => n5765);
   U84521 : OAI22_X1 port map( A1 => n120312, A2 => n114435, B1 => n120652, B2 
                           => n120304, ZN => n5766);
   U84522 : OAI22_X1 port map( A1 => n120312, A2 => n114434, B1 => n120655, B2 
                           => n120304, ZN => n5767);
   U84523 : OAI22_X1 port map( A1 => n120312, A2 => n114433, B1 => n120658, B2 
                           => n120304, ZN => n5768);
   U84524 : OAI22_X1 port map( A1 => n120312, A2 => n114432, B1 => n120661, B2 
                           => n120304, ZN => n5769);
   U84525 : OAI22_X1 port map( A1 => n120312, A2 => n114431, B1 => n120664, B2 
                           => n120304, ZN => n5770);
   U84526 : OAI22_X1 port map( A1 => n120313, A2 => n114430, B1 => n120667, B2 
                           => n120305, ZN => n5771);
   U84527 : OAI22_X1 port map( A1 => n120313, A2 => n114429, B1 => n120670, B2 
                           => n120305, ZN => n5772);
   U84528 : OAI22_X1 port map( A1 => n120313, A2 => n114428, B1 => n120673, B2 
                           => n120305, ZN => n5773);
   U84529 : OAI22_X1 port map( A1 => n120313, A2 => n114427, B1 => n120676, B2 
                           => n120305, ZN => n5774);
   U84530 : OAI22_X1 port map( A1 => n120313, A2 => n114426, B1 => n120679, B2 
                           => n120305, ZN => n5775);
   U84531 : OAI22_X1 port map( A1 => n120313, A2 => n114425, B1 => n120682, B2 
                           => n120305, ZN => n5776);
   U84532 : OAI22_X1 port map( A1 => n120313, A2 => n114424, B1 => n120685, B2 
                           => n120305, ZN => n5777);
   U84533 : OAI22_X1 port map( A1 => n120313, A2 => n114423, B1 => n120688, B2 
                           => n120305, ZN => n5778);
   U84534 : OAI22_X1 port map( A1 => n120313, A2 => n114422, B1 => n120691, B2 
                           => n120305, ZN => n5779);
   U84535 : OAI22_X1 port map( A1 => n120313, A2 => n114421, B1 => n120694, B2 
                           => n120305, ZN => n5780);
   U84536 : OAI22_X1 port map( A1 => n120313, A2 => n114420, B1 => n120697, B2 
                           => n120305, ZN => n5781);
   U84537 : OAI22_X1 port map( A1 => n120313, A2 => n114419, B1 => n120700, B2 
                           => n120305, ZN => n5782);
   U84538 : OAI22_X1 port map( A1 => n120313, A2 => n114418, B1 => n120703, B2 
                           => n120306, ZN => n5783);
   U84539 : OAI22_X1 port map( A1 => n120314, A2 => n114417, B1 => n120706, B2 
                           => n120306, ZN => n5784);
   U84540 : OAI22_X1 port map( A1 => n120314, A2 => n114416, B1 => n120709, B2 
                           => n120306, ZN => n5785);
   U84541 : OAI22_X1 port map( A1 => n120314, A2 => n114415, B1 => n120712, B2 
                           => n120306, ZN => n5786);
   U84542 : OAI22_X1 port map( A1 => n120314, A2 => n114414, B1 => n120715, B2 
                           => n120306, ZN => n5787);
   U84543 : OAI22_X1 port map( A1 => n120314, A2 => n114413, B1 => n120718, B2 
                           => n120306, ZN => n5788);
   U84544 : OAI22_X1 port map( A1 => n120314, A2 => n114412, B1 => n120721, B2 
                           => n120306, ZN => n5789);
   U84545 : OAI22_X1 port map( A1 => n120314, A2 => n114411, B1 => n120724, B2 
                           => n120306, ZN => n5790);
   U84546 : OAI22_X1 port map( A1 => n120314, A2 => n114410, B1 => n120727, B2 
                           => n120306, ZN => n5791);
   U84547 : OAI22_X1 port map( A1 => n120314, A2 => n114409, B1 => n120730, B2 
                           => n120306, ZN => n5792);
   U84548 : OAI22_X1 port map( A1 => n120314, A2 => n114408, B1 => n120733, B2 
                           => n120306, ZN => n5793);
   U84549 : OAI22_X1 port map( A1 => n120314, A2 => n114407, B1 => n120736, B2 
                           => n120306, ZN => n5794);
   U84550 : OAI22_X1 port map( A1 => n120314, A2 => n114406, B1 => n120739, B2 
                           => n120307, ZN => n5795);
   U84551 : OAI22_X1 port map( A1 => n120314, A2 => n114405, B1 => n120742, B2 
                           => n120307, ZN => n5796);
   U84552 : OAI22_X1 port map( A1 => n120315, A2 => n114404, B1 => n120745, B2 
                           => n120307, ZN => n5797);
   U84553 : OAI22_X1 port map( A1 => n120315, A2 => n114403, B1 => n120748, B2 
                           => n120307, ZN => n5798);
   U84554 : OAI22_X1 port map( A1 => n120315, A2 => n114402, B1 => n120751, B2 
                           => n120307, ZN => n5799);
   U84555 : OAI22_X1 port map( A1 => n120315, A2 => n114401, B1 => n120754, B2 
                           => n120307, ZN => n5800);
   U84556 : OAI22_X1 port map( A1 => n120315, A2 => n114400, B1 => n120757, B2 
                           => n120307, ZN => n5801);
   U84557 : OAI22_X1 port map( A1 => n120315, A2 => n114399, B1 => n120760, B2 
                           => n120307, ZN => n5802);
   U84558 : OAI22_X1 port map( A1 => n120315, A2 => n114398, B1 => n120763, B2 
                           => n120307, ZN => n5803);
   U84559 : OAI22_X1 port map( A1 => n120315, A2 => n114397, B1 => n120766, B2 
                           => n120307, ZN => n5804);
   U84560 : OAI22_X1 port map( A1 => n120315, A2 => n114396, B1 => n120769, B2 
                           => n120307, ZN => n5805);
   U84561 : OAI22_X1 port map( A1 => n120315, A2 => n114395, B1 => n120772, B2 
                           => n120307, ZN => n5806);
   U84562 : OAI22_X1 port map( A1 => n120315, A2 => n114394, B1 => n120775, B2 
                           => n120308, ZN => n5807);
   U84563 : OAI22_X1 port map( A1 => n120315, A2 => n114393, B1 => n120778, B2 
                           => n120308, ZN => n5808);
   U84564 : OAI22_X1 port map( A1 => n120315, A2 => n114392, B1 => n120781, B2 
                           => n120308, ZN => n5809);
   U84565 : OAI22_X1 port map( A1 => n120316, A2 => n114391, B1 => n120784, B2 
                           => n120308, ZN => n5810);
   U84566 : OAI22_X1 port map( A1 => n120316, A2 => n114390, B1 => n120787, B2 
                           => n120308, ZN => n5811);
   U84567 : OAI22_X1 port map( A1 => n120316, A2 => n114389, B1 => n120790, B2 
                           => n120308, ZN => n5812);
   U84568 : OAI22_X1 port map( A1 => n120316, A2 => n114388, B1 => n120793, B2 
                           => n120308, ZN => n5813);
   U84569 : OAI22_X1 port map( A1 => n120316, A2 => n114387, B1 => n120796, B2 
                           => n120308, ZN => n5814);
   U84570 : OAI22_X1 port map( A1 => n120316, A2 => n114386, B1 => n120799, B2 
                           => n120308, ZN => n5815);
   U84571 : OAI22_X1 port map( A1 => n120316, A2 => n114385, B1 => n120802, B2 
                           => n120308, ZN => n5816);
   U84572 : OAI22_X1 port map( A1 => n120316, A2 => n114384, B1 => n120805, B2 
                           => n120308, ZN => n5817);
   U84573 : OAI22_X1 port map( A1 => n120299, A2 => n114508, B1 => n120631, B2 
                           => n120291, ZN => n5695);
   U84574 : OAI22_X1 port map( A1 => n120299, A2 => n114507, B1 => n120634, B2 
                           => n120291, ZN => n5696);
   U84575 : OAI22_X1 port map( A1 => n120299, A2 => n114506, B1 => n120637, B2 
                           => n120291, ZN => n5697);
   U84576 : OAI22_X1 port map( A1 => n120299, A2 => n114505, B1 => n120640, B2 
                           => n120291, ZN => n5698);
   U84577 : OAI22_X1 port map( A1 => n120299, A2 => n114504, B1 => n120643, B2 
                           => n120291, ZN => n5699);
   U84578 : OAI22_X1 port map( A1 => n120299, A2 => n114503, B1 => n120646, B2 
                           => n120291, ZN => n5700);
   U84579 : OAI22_X1 port map( A1 => n120299, A2 => n114502, B1 => n120649, B2 
                           => n120291, ZN => n5701);
   U84580 : OAI22_X1 port map( A1 => n120299, A2 => n114501, B1 => n120652, B2 
                           => n120291, ZN => n5702);
   U84581 : OAI22_X1 port map( A1 => n120299, A2 => n114500, B1 => n120655, B2 
                           => n120291, ZN => n5703);
   U84582 : OAI22_X1 port map( A1 => n120299, A2 => n114499, B1 => n120658, B2 
                           => n120291, ZN => n5704);
   U84583 : OAI22_X1 port map( A1 => n120299, A2 => n114498, B1 => n120661, B2 
                           => n120291, ZN => n5705);
   U84584 : OAI22_X1 port map( A1 => n120299, A2 => n114497, B1 => n120664, B2 
                           => n120291, ZN => n5706);
   U84585 : OAI22_X1 port map( A1 => n120300, A2 => n114496, B1 => n120667, B2 
                           => n120292, ZN => n5707);
   U84586 : OAI22_X1 port map( A1 => n120300, A2 => n114495, B1 => n120670, B2 
                           => n120292, ZN => n5708);
   U84587 : OAI22_X1 port map( A1 => n120300, A2 => n114494, B1 => n120673, B2 
                           => n120292, ZN => n5709);
   U84588 : OAI22_X1 port map( A1 => n120300, A2 => n114493, B1 => n120676, B2 
                           => n120292, ZN => n5710);
   U84589 : OAI22_X1 port map( A1 => n120300, A2 => n114492, B1 => n120679, B2 
                           => n120292, ZN => n5711);
   U84590 : OAI22_X1 port map( A1 => n120300, A2 => n114491, B1 => n120682, B2 
                           => n120292, ZN => n5712);
   U84591 : OAI22_X1 port map( A1 => n120300, A2 => n114490, B1 => n120685, B2 
                           => n120292, ZN => n5713);
   U84592 : OAI22_X1 port map( A1 => n120300, A2 => n114489, B1 => n120688, B2 
                           => n120292, ZN => n5714);
   U84593 : OAI22_X1 port map( A1 => n120300, A2 => n114488, B1 => n120691, B2 
                           => n120292, ZN => n5715);
   U84594 : OAI22_X1 port map( A1 => n120300, A2 => n114487, B1 => n120694, B2 
                           => n120292, ZN => n5716);
   U84595 : OAI22_X1 port map( A1 => n120300, A2 => n114486, B1 => n120697, B2 
                           => n120292, ZN => n5717);
   U84596 : OAI22_X1 port map( A1 => n120300, A2 => n114485, B1 => n120700, B2 
                           => n120292, ZN => n5718);
   U84597 : OAI22_X1 port map( A1 => n120300, A2 => n114484, B1 => n120703, B2 
                           => n120293, ZN => n5719);
   U84598 : OAI22_X1 port map( A1 => n120301, A2 => n114483, B1 => n120706, B2 
                           => n120293, ZN => n5720);
   U84599 : OAI22_X1 port map( A1 => n120301, A2 => n114482, B1 => n120709, B2 
                           => n120293, ZN => n5721);
   U84600 : OAI22_X1 port map( A1 => n120301, A2 => n114481, B1 => n120712, B2 
                           => n120293, ZN => n5722);
   U84601 : OAI22_X1 port map( A1 => n120301, A2 => n114480, B1 => n120715, B2 
                           => n120293, ZN => n5723);
   U84602 : OAI22_X1 port map( A1 => n120301, A2 => n114479, B1 => n120718, B2 
                           => n120293, ZN => n5724);
   U84603 : OAI22_X1 port map( A1 => n120301, A2 => n114478, B1 => n120721, B2 
                           => n120293, ZN => n5725);
   U84604 : OAI22_X1 port map( A1 => n120301, A2 => n114477, B1 => n120724, B2 
                           => n120293, ZN => n5726);
   U84605 : OAI22_X1 port map( A1 => n120301, A2 => n114476, B1 => n120727, B2 
                           => n120293, ZN => n5727);
   U84606 : OAI22_X1 port map( A1 => n120301, A2 => n114475, B1 => n120730, B2 
                           => n120293, ZN => n5728);
   U84607 : OAI22_X1 port map( A1 => n120301, A2 => n114474, B1 => n120733, B2 
                           => n120293, ZN => n5729);
   U84608 : OAI22_X1 port map( A1 => n120301, A2 => n114473, B1 => n120736, B2 
                           => n120293, ZN => n5730);
   U84609 : OAI22_X1 port map( A1 => n120301, A2 => n114472, B1 => n120739, B2 
                           => n120294, ZN => n5731);
   U84610 : OAI22_X1 port map( A1 => n120301, A2 => n114471, B1 => n120742, B2 
                           => n120294, ZN => n5732);
   U84611 : OAI22_X1 port map( A1 => n120302, A2 => n114470, B1 => n120745, B2 
                           => n120294, ZN => n5733);
   U84612 : OAI22_X1 port map( A1 => n120302, A2 => n114469, B1 => n120748, B2 
                           => n120294, ZN => n5734);
   U84613 : OAI22_X1 port map( A1 => n120302, A2 => n114468, B1 => n120751, B2 
                           => n120294, ZN => n5735);
   U84614 : OAI22_X1 port map( A1 => n120302, A2 => n114467, B1 => n120754, B2 
                           => n120294, ZN => n5736);
   U84615 : OAI22_X1 port map( A1 => n120302, A2 => n114466, B1 => n120757, B2 
                           => n120294, ZN => n5737);
   U84616 : OAI22_X1 port map( A1 => n120302, A2 => n114465, B1 => n120760, B2 
                           => n120294, ZN => n5738);
   U84617 : OAI22_X1 port map( A1 => n120302, A2 => n114464, B1 => n120763, B2 
                           => n120294, ZN => n5739);
   U84618 : OAI22_X1 port map( A1 => n120302, A2 => n114463, B1 => n120766, B2 
                           => n120294, ZN => n5740);
   U84619 : OAI22_X1 port map( A1 => n120302, A2 => n114462, B1 => n120769, B2 
                           => n120294, ZN => n5741);
   U84620 : OAI22_X1 port map( A1 => n120302, A2 => n114461, B1 => n120772, B2 
                           => n120294, ZN => n5742);
   U84621 : OAI22_X1 port map( A1 => n120302, A2 => n114460, B1 => n120775, B2 
                           => n120295, ZN => n5743);
   U84622 : OAI22_X1 port map( A1 => n120302, A2 => n114459, B1 => n120778, B2 
                           => n120295, ZN => n5744);
   U84623 : OAI22_X1 port map( A1 => n120302, A2 => n114458, B1 => n120781, B2 
                           => n120295, ZN => n5745);
   U84624 : OAI22_X1 port map( A1 => n120303, A2 => n114457, B1 => n120784, B2 
                           => n120295, ZN => n5746);
   U84625 : OAI22_X1 port map( A1 => n120303, A2 => n114456, B1 => n120787, B2 
                           => n120295, ZN => n5747);
   U84626 : OAI22_X1 port map( A1 => n120303, A2 => n114455, B1 => n120790, B2 
                           => n120295, ZN => n5748);
   U84627 : OAI22_X1 port map( A1 => n120303, A2 => n114454, B1 => n120793, B2 
                           => n120295, ZN => n5749);
   U84628 : OAI22_X1 port map( A1 => n120303, A2 => n114453, B1 => n120796, B2 
                           => n120295, ZN => n5750);
   U84629 : OAI22_X1 port map( A1 => n120303, A2 => n114452, B1 => n120799, B2 
                           => n120295, ZN => n5751);
   U84630 : OAI22_X1 port map( A1 => n120303, A2 => n114451, B1 => n120802, B2 
                           => n120295, ZN => n5752);
   U84631 : OAI22_X1 port map( A1 => n120303, A2 => n114450, B1 => n120805, B2 
                           => n120295, ZN => n5753);
   U84632 : OAI22_X1 port map( A1 => n120303, A2 => n114449, B1 => n120808, B2 
                           => n120295, ZN => n5754);
   U84633 : OAI22_X1 port map( A1 => n120316, A2 => n114383, B1 => n120808, B2 
                           => n120308, ZN => n5818);
   U84634 : OAI22_X1 port map( A1 => n120545, A2 => n114051, B1 => n120629, B2 
                           => n120537, ZN => n6975);
   U84635 : OAI22_X1 port map( A1 => n120549, A2 => n114050, B1 => n120632, B2 
                           => n120537, ZN => n6976);
   U84636 : OAI22_X1 port map( A1 => n120549, A2 => n114049, B1 => n120635, B2 
                           => n120537, ZN => n6977);
   U84637 : OAI22_X1 port map( A1 => n120549, A2 => n114048, B1 => n120638, B2 
                           => n120537, ZN => n6978);
   U84638 : OAI22_X1 port map( A1 => n120549, A2 => n114047, B1 => n120641, B2 
                           => n120537, ZN => n6979);
   U84639 : OAI22_X1 port map( A1 => n120549, A2 => n114046, B1 => n120644, B2 
                           => n120537, ZN => n6980);
   U84640 : OAI22_X1 port map( A1 => n120549, A2 => n114045, B1 => n120647, B2 
                           => n120537, ZN => n6981);
   U84641 : OAI22_X1 port map( A1 => n120549, A2 => n114044, B1 => n120650, B2 
                           => n120537, ZN => n6982);
   U84642 : OAI22_X1 port map( A1 => n120549, A2 => n114043, B1 => n120653, B2 
                           => n120537, ZN => n6983);
   U84643 : OAI22_X1 port map( A1 => n120549, A2 => n114042, B1 => n120656, B2 
                           => n120537, ZN => n6984);
   U84644 : OAI22_X1 port map( A1 => n120549, A2 => n114041, B1 => n120659, B2 
                           => n120537, ZN => n6985);
   U84645 : OAI22_X1 port map( A1 => n120549, A2 => n114040, B1 => n120662, B2 
                           => n120537, ZN => n6986);
   U84646 : OAI22_X1 port map( A1 => n120549, A2 => n114039, B1 => n120665, B2 
                           => n120538, ZN => n6987);
   U84647 : OAI22_X1 port map( A1 => n120549, A2 => n114038, B1 => n120668, B2 
                           => n120538, ZN => n6988);
   U84648 : OAI22_X1 port map( A1 => n120548, A2 => n114037, B1 => n120671, B2 
                           => n120538, ZN => n6989);
   U84649 : OAI22_X1 port map( A1 => n120548, A2 => n114036, B1 => n120674, B2 
                           => n120538, ZN => n6990);
   U84650 : OAI22_X1 port map( A1 => n120548, A2 => n114035, B1 => n120677, B2 
                           => n120538, ZN => n6991);
   U84651 : OAI22_X1 port map( A1 => n120548, A2 => n114034, B1 => n120680, B2 
                           => n120538, ZN => n6992);
   U84652 : OAI22_X1 port map( A1 => n120548, A2 => n114033, B1 => n120683, B2 
                           => n120538, ZN => n6993);
   U84653 : OAI22_X1 port map( A1 => n120548, A2 => n114032, B1 => n120686, B2 
                           => n120538, ZN => n6994);
   U84654 : OAI22_X1 port map( A1 => n120548, A2 => n114031, B1 => n120689, B2 
                           => n120538, ZN => n6995);
   U84655 : OAI22_X1 port map( A1 => n120548, A2 => n114030, B1 => n120692, B2 
                           => n120538, ZN => n6996);
   U84656 : OAI22_X1 port map( A1 => n120548, A2 => n114029, B1 => n120695, B2 
                           => n120538, ZN => n6997);
   U84657 : OAI22_X1 port map( A1 => n120548, A2 => n114028, B1 => n120698, B2 
                           => n120538, ZN => n6998);
   U84658 : OAI22_X1 port map( A1 => n120548, A2 => n114027, B1 => n120701, B2 
                           => n120539, ZN => n6999);
   U84659 : OAI22_X1 port map( A1 => n120548, A2 => n114026, B1 => n120704, B2 
                           => n120539, ZN => n7000);
   U84660 : OAI22_X1 port map( A1 => n120548, A2 => n114025, B1 => n120707, B2 
                           => n120539, ZN => n7001);
   U84661 : OAI22_X1 port map( A1 => n120547, A2 => n114024, B1 => n120710, B2 
                           => n120539, ZN => n7002);
   U84662 : OAI22_X1 port map( A1 => n120547, A2 => n114023, B1 => n120713, B2 
                           => n120539, ZN => n7003);
   U84663 : OAI22_X1 port map( A1 => n120547, A2 => n114022, B1 => n120716, B2 
                           => n120539, ZN => n7004);
   U84664 : OAI22_X1 port map( A1 => n120547, A2 => n114021, B1 => n120719, B2 
                           => n120539, ZN => n7005);
   U84665 : OAI22_X1 port map( A1 => n120547, A2 => n114020, B1 => n120722, B2 
                           => n120539, ZN => n7006);
   U84666 : OAI22_X1 port map( A1 => n120547, A2 => n114019, B1 => n120725, B2 
                           => n120539, ZN => n7007);
   U84667 : OAI22_X1 port map( A1 => n120547, A2 => n114018, B1 => n120728, B2 
                           => n120539, ZN => n7008);
   U84668 : OAI22_X1 port map( A1 => n120547, A2 => n114017, B1 => n120731, B2 
                           => n120539, ZN => n7009);
   U84669 : OAI22_X1 port map( A1 => n120547, A2 => n114016, B1 => n120734, B2 
                           => n120539, ZN => n7010);
   U84670 : OAI22_X1 port map( A1 => n120547, A2 => n114015, B1 => n120737, B2 
                           => n120540, ZN => n7011);
   U84671 : OAI22_X1 port map( A1 => n120547, A2 => n114014, B1 => n120740, B2 
                           => n120540, ZN => n7012);
   U84672 : OAI22_X1 port map( A1 => n120547, A2 => n114013, B1 => n120743, B2 
                           => n120540, ZN => n7013);
   U84673 : OAI22_X1 port map( A1 => n120546, A2 => n114012, B1 => n120746, B2 
                           => n120540, ZN => n7014);
   U84674 : OAI22_X1 port map( A1 => n120546, A2 => n114011, B1 => n120749, B2 
                           => n120540, ZN => n7015);
   U84675 : OAI22_X1 port map( A1 => n120546, A2 => n114010, B1 => n120752, B2 
                           => n120540, ZN => n7016);
   U84676 : OAI22_X1 port map( A1 => n120546, A2 => n114009, B1 => n120755, B2 
                           => n120540, ZN => n7017);
   U84677 : OAI22_X1 port map( A1 => n120546, A2 => n114008, B1 => n120758, B2 
                           => n120540, ZN => n7018);
   U84678 : OAI22_X1 port map( A1 => n120546, A2 => n114007, B1 => n120761, B2 
                           => n120540, ZN => n7019);
   U84679 : OAI22_X1 port map( A1 => n120546, A2 => n114006, B1 => n120764, B2 
                           => n120540, ZN => n7020);
   U84680 : OAI22_X1 port map( A1 => n120546, A2 => n114005, B1 => n120767, B2 
                           => n120540, ZN => n7021);
   U84681 : OAI22_X1 port map( A1 => n120547, A2 => n114004, B1 => n120770, B2 
                           => n120540, ZN => n7022);
   U84682 : OAI22_X1 port map( A1 => n120546, A2 => n114003, B1 => n120773, B2 
                           => n120541, ZN => n7023);
   U84683 : OAI22_X1 port map( A1 => n120546, A2 => n114002, B1 => n120776, B2 
                           => n120541, ZN => n7024);
   U84684 : OAI22_X1 port map( A1 => n120546, A2 => n114001, B1 => n120779, B2 
                           => n120541, ZN => n7025);
   U84685 : OAI22_X1 port map( A1 => n120546, A2 => n114000, B1 => n120782, B2 
                           => n120541, ZN => n7026);
   U84686 : OAI22_X1 port map( A1 => n120546, A2 => n113999, B1 => n120785, B2 
                           => n120541, ZN => n7027);
   U84687 : OAI22_X1 port map( A1 => n120545, A2 => n113998, B1 => n120788, B2 
                           => n120541, ZN => n7028);
   U84688 : OAI22_X1 port map( A1 => n120545, A2 => n113997, B1 => n120791, B2 
                           => n120541, ZN => n7029);
   U84689 : OAI22_X1 port map( A1 => n120545, A2 => n113996, B1 => n120794, B2 
                           => n120541, ZN => n7030);
   U84690 : OAI22_X1 port map( A1 => n120545, A2 => n113995, B1 => n120797, B2 
                           => n120541, ZN => n7031);
   U84691 : OAI22_X1 port map( A1 => n120545, A2 => n113994, B1 => n120800, B2 
                           => n120541, ZN => n7032);
   U84692 : OAI22_X1 port map( A1 => n120545, A2 => n113993, B1 => n120803, B2 
                           => n120541, ZN => n7033);
   U84693 : OAI22_X1 port map( A1 => n120545, A2 => n113992, B1 => n120806, B2 
                           => n120541, ZN => n7034);
   U84694 : OAI22_X1 port map( A1 => n120829, A2 => n113890, B1 => n120821, B2 
                           => n120629, ZN => n7423);
   U84695 : OAI22_X1 port map( A1 => n120833, A2 => n113888, B1 => n120821, B2 
                           => n120632, ZN => n7424);
   U84696 : OAI22_X1 port map( A1 => n120833, A2 => n113886, B1 => n120821, B2 
                           => n120635, ZN => n7425);
   U84697 : OAI22_X1 port map( A1 => n120833, A2 => n113884, B1 => n120821, B2 
                           => n120638, ZN => n7426);
   U84698 : OAI22_X1 port map( A1 => n120833, A2 => n113882, B1 => n120821, B2 
                           => n120641, ZN => n7427);
   U84699 : OAI22_X1 port map( A1 => n120833, A2 => n113880, B1 => n120821, B2 
                           => n120644, ZN => n7428);
   U84700 : OAI22_X1 port map( A1 => n120833, A2 => n113878, B1 => n120821, B2 
                           => n120647, ZN => n7429);
   U84701 : OAI22_X1 port map( A1 => n120833, A2 => n113876, B1 => n120821, B2 
                           => n120650, ZN => n7430);
   U84702 : OAI22_X1 port map( A1 => n120833, A2 => n113874, B1 => n120821, B2 
                           => n120653, ZN => n7431);
   U84703 : OAI22_X1 port map( A1 => n120833, A2 => n113872, B1 => n120821, B2 
                           => n120656, ZN => n7432);
   U84704 : OAI22_X1 port map( A1 => n120833, A2 => n113870, B1 => n120821, B2 
                           => n120659, ZN => n7433);
   U84705 : OAI22_X1 port map( A1 => n120833, A2 => n113868, B1 => n120821, B2 
                           => n120662, ZN => n7434);
   U84706 : OAI22_X1 port map( A1 => n120390, A2 => n114233, B1 => n120630, B2 
                           => n120379, ZN => n6143);
   U84707 : OAI22_X1 port map( A1 => n120390, A2 => n114232, B1 => n120633, B2 
                           => n120379, ZN => n6144);
   U84708 : OAI22_X1 port map( A1 => n120390, A2 => n114231, B1 => n120636, B2 
                           => n120379, ZN => n6145);
   U84709 : OAI22_X1 port map( A1 => n120390, A2 => n114230, B1 => n120639, B2 
                           => n120379, ZN => n6146);
   U84710 : OAI22_X1 port map( A1 => n120389, A2 => n114229, B1 => n120642, B2 
                           => n120379, ZN => n6147);
   U84711 : OAI22_X1 port map( A1 => n120389, A2 => n114228, B1 => n120645, B2 
                           => n120379, ZN => n6148);
   U84712 : OAI22_X1 port map( A1 => n120389, A2 => n114227, B1 => n120648, B2 
                           => n120379, ZN => n6149);
   U84713 : OAI22_X1 port map( A1 => n120389, A2 => n114226, B1 => n120651, B2 
                           => n120379, ZN => n6150);
   U84714 : OAI22_X1 port map( A1 => n120389, A2 => n114225, B1 => n120654, B2 
                           => n120379, ZN => n6151);
   U84715 : OAI22_X1 port map( A1 => n120389, A2 => n114224, B1 => n120657, B2 
                           => n120379, ZN => n6152);
   U84716 : OAI22_X1 port map( A1 => n120389, A2 => n114223, B1 => n120660, B2 
                           => n120379, ZN => n6153);
   U84717 : OAI22_X1 port map( A1 => n120389, A2 => n114222, B1 => n120663, B2 
                           => n120379, ZN => n6154);
   U84718 : OAI22_X1 port map( A1 => n120389, A2 => n114221, B1 => n120666, B2 
                           => n120380, ZN => n6155);
   U84719 : OAI22_X1 port map( A1 => n120389, A2 => n114220, B1 => n120669, B2 
                           => n120380, ZN => n6156);
   U84720 : OAI22_X1 port map( A1 => n120389, A2 => n114219, B1 => n120672, B2 
                           => n120380, ZN => n6157);
   U84721 : OAI22_X1 port map( A1 => n120389, A2 => n114218, B1 => n120675, B2 
                           => n120380, ZN => n6158);
   U84722 : OAI22_X1 port map( A1 => n120389, A2 => n114217, B1 => n120678, B2 
                           => n120380, ZN => n6159);
   U84723 : OAI22_X1 port map( A1 => n120388, A2 => n114216, B1 => n120681, B2 
                           => n120380, ZN => n6160);
   U84724 : OAI22_X1 port map( A1 => n120388, A2 => n114215, B1 => n120684, B2 
                           => n120380, ZN => n6161);
   U84725 : OAI22_X1 port map( A1 => n120570, A2 => n113979, B1 => n120629, B2 
                           => n120562, ZN => n7103);
   U84726 : OAI22_X1 port map( A1 => n120570, A2 => n113978, B1 => n120632, B2 
                           => n120562, ZN => n7104);
   U84727 : OAI22_X1 port map( A1 => n120570, A2 => n113977, B1 => n120635, B2 
                           => n120562, ZN => n7105);
   U84728 : OAI22_X1 port map( A1 => n120570, A2 => n113976, B1 => n120638, B2 
                           => n120562, ZN => n7106);
   U84729 : OAI22_X1 port map( A1 => n120570, A2 => n113975, B1 => n120641, B2 
                           => n120562, ZN => n7107);
   U84730 : OAI22_X1 port map( A1 => n120570, A2 => n113974, B1 => n120644, B2 
                           => n120562, ZN => n7108);
   U84731 : OAI22_X1 port map( A1 => n120570, A2 => n113973, B1 => n120647, B2 
                           => n120562, ZN => n7109);
   U84732 : OAI22_X1 port map( A1 => n120570, A2 => n113972, B1 => n120650, B2 
                           => n120562, ZN => n7110);
   U84733 : OAI22_X1 port map( A1 => n120570, A2 => n113971, B1 => n120653, B2 
                           => n120562, ZN => n7111);
   U84734 : OAI22_X1 port map( A1 => n120570, A2 => n113970, B1 => n120656, B2 
                           => n120562, ZN => n7112);
   U84735 : OAI22_X1 port map( A1 => n120570, A2 => n113969, B1 => n120659, B2 
                           => n120562, ZN => n7113);
   U84736 : OAI22_X1 port map( A1 => n120570, A2 => n113968, B1 => n120662, B2 
                           => n120562, ZN => n7114);
   U84737 : OAI22_X1 port map( A1 => n120571, A2 => n113967, B1 => n120665, B2 
                           => n120563, ZN => n7115);
   U84738 : OAI22_X1 port map( A1 => n120571, A2 => n113966, B1 => n120668, B2 
                           => n120563, ZN => n7116);
   U84739 : OAI22_X1 port map( A1 => n120571, A2 => n113965, B1 => n120671, B2 
                           => n120563, ZN => n7117);
   U84740 : OAI22_X1 port map( A1 => n120571, A2 => n113964, B1 => n120674, B2 
                           => n120563, ZN => n7118);
   U84741 : OAI22_X1 port map( A1 => n120571, A2 => n113963, B1 => n120677, B2 
                           => n120563, ZN => n7119);
   U84742 : OAI22_X1 port map( A1 => n120571, A2 => n113962, B1 => n120680, B2 
                           => n120563, ZN => n7120);
   U84743 : OAI22_X1 port map( A1 => n120571, A2 => n113961, B1 => n120683, B2 
                           => n120563, ZN => n7121);
   U84744 : OAI22_X1 port map( A1 => n120571, A2 => n113960, B1 => n120686, B2 
                           => n120563, ZN => n7122);
   U84745 : OAI22_X1 port map( A1 => n120571, A2 => n113959, B1 => n120689, B2 
                           => n120563, ZN => n7123);
   U84746 : OAI22_X1 port map( A1 => n120571, A2 => n113958, B1 => n120692, B2 
                           => n120563, ZN => n7124);
   U84747 : OAI22_X1 port map( A1 => n120571, A2 => n113957, B1 => n120695, B2 
                           => n120563, ZN => n7125);
   U84748 : OAI22_X1 port map( A1 => n120571, A2 => n113956, B1 => n120698, B2 
                           => n120563, ZN => n7126);
   U84749 : OAI22_X1 port map( A1 => n120571, A2 => n113955, B1 => n120701, B2 
                           => n120564, ZN => n7127);
   U84750 : OAI22_X1 port map( A1 => n120572, A2 => n113954, B1 => n120704, B2 
                           => n120564, ZN => n7128);
   U84751 : OAI22_X1 port map( A1 => n120572, A2 => n113953, B1 => n120707, B2 
                           => n120564, ZN => n7129);
   U84752 : OAI22_X1 port map( A1 => n120572, A2 => n113952, B1 => n120710, B2 
                           => n120564, ZN => n7130);
   U84753 : OAI22_X1 port map( A1 => n120572, A2 => n113951, B1 => n120713, B2 
                           => n120564, ZN => n7131);
   U84754 : OAI22_X1 port map( A1 => n120572, A2 => n113950, B1 => n120716, B2 
                           => n120564, ZN => n7132);
   U84755 : OAI22_X1 port map( A1 => n120572, A2 => n113949, B1 => n120719, B2 
                           => n120564, ZN => n7133);
   U84756 : OAI22_X1 port map( A1 => n120572, A2 => n113948, B1 => n120722, B2 
                           => n120564, ZN => n7134);
   U84757 : OAI22_X1 port map( A1 => n120572, A2 => n113947, B1 => n120725, B2 
                           => n120564, ZN => n7135);
   U84758 : OAI22_X1 port map( A1 => n120572, A2 => n113946, B1 => n120728, B2 
                           => n120564, ZN => n7136);
   U84759 : OAI22_X1 port map( A1 => n120572, A2 => n113945, B1 => n120731, B2 
                           => n120564, ZN => n7137);
   U84760 : OAI22_X1 port map( A1 => n120572, A2 => n113944, B1 => n120734, B2 
                           => n120564, ZN => n7138);
   U84761 : OAI22_X1 port map( A1 => n120572, A2 => n113943, B1 => n120737, B2 
                           => n120565, ZN => n7139);
   U84762 : OAI22_X1 port map( A1 => n120572, A2 => n113942, B1 => n120740, B2 
                           => n120565, ZN => n7140);
   U84763 : OAI22_X1 port map( A1 => n120573, A2 => n113941, B1 => n120743, B2 
                           => n120565, ZN => n7141);
   U84764 : OAI22_X1 port map( A1 => n120573, A2 => n113940, B1 => n120746, B2 
                           => n120565, ZN => n7142);
   U84765 : OAI22_X1 port map( A1 => n120573, A2 => n113939, B1 => n120749, B2 
                           => n120565, ZN => n7143);
   U84766 : OAI22_X1 port map( A1 => n120573, A2 => n113938, B1 => n120752, B2 
                           => n120565, ZN => n7144);
   U84767 : OAI22_X1 port map( A1 => n120573, A2 => n113937, B1 => n120755, B2 
                           => n120565, ZN => n7145);
   U84768 : OAI22_X1 port map( A1 => n120573, A2 => n113936, B1 => n120758, B2 
                           => n120565, ZN => n7146);
   U84769 : OAI22_X1 port map( A1 => n120573, A2 => n113935, B1 => n120761, B2 
                           => n120565, ZN => n7147);
   U84770 : OAI22_X1 port map( A1 => n120573, A2 => n113934, B1 => n120764, B2 
                           => n120565, ZN => n7148);
   U84771 : OAI22_X1 port map( A1 => n120573, A2 => n113933, B1 => n120767, B2 
                           => n120565, ZN => n7149);
   U84772 : OAI22_X1 port map( A1 => n120573, A2 => n113932, B1 => n120770, B2 
                           => n120565, ZN => n7150);
   U84773 : OAI22_X1 port map( A1 => n120573, A2 => n113931, B1 => n120773, B2 
                           => n120566, ZN => n7151);
   U84774 : OAI22_X1 port map( A1 => n120573, A2 => n113930, B1 => n120776, B2 
                           => n120566, ZN => n7152);
   U84775 : OAI22_X1 port map( A1 => n120573, A2 => n113929, B1 => n120779, B2 
                           => n120566, ZN => n7153);
   U84776 : OAI22_X1 port map( A1 => n120574, A2 => n113928, B1 => n120782, B2 
                           => n120566, ZN => n7154);
   U84777 : OAI22_X1 port map( A1 => n120574, A2 => n113927, B1 => n120785, B2 
                           => n120566, ZN => n7155);
   U84778 : OAI22_X1 port map( A1 => n120574, A2 => n113926, B1 => n120788, B2 
                           => n120566, ZN => n7156);
   U84779 : OAI22_X1 port map( A1 => n120574, A2 => n113925, B1 => n120791, B2 
                           => n120566, ZN => n7157);
   U84780 : OAI22_X1 port map( A1 => n120574, A2 => n113924, B1 => n120794, B2 
                           => n120566, ZN => n7158);
   U84781 : OAI22_X1 port map( A1 => n120574, A2 => n113923, B1 => n120797, B2 
                           => n120566, ZN => n7159);
   U84782 : OAI22_X1 port map( A1 => n120574, A2 => n113922, B1 => n120800, B2 
                           => n120566, ZN => n7160);
   U84783 : OAI22_X1 port map( A1 => n120574, A2 => n113921, B1 => n120803, B2 
                           => n120566, ZN => n7161);
   U84784 : OAI22_X1 port map( A1 => n120574, A2 => n113920, B1 => n120806, B2 
                           => n120566, ZN => n7162);
   U84785 : OAI22_X1 port map( A1 => n120374, A2 => n114299, B1 => n120630, B2 
                           => n120366, ZN => n6079);
   U84786 : OAI22_X1 port map( A1 => n120374, A2 => n114298, B1 => n120633, B2 
                           => n120366, ZN => n6080);
   U84787 : OAI22_X1 port map( A1 => n120374, A2 => n114297, B1 => n120636, B2 
                           => n120366, ZN => n6081);
   U84788 : OAI22_X1 port map( A1 => n120374, A2 => n114296, B1 => n120639, B2 
                           => n120366, ZN => n6082);
   U84789 : OAI22_X1 port map( A1 => n120374, A2 => n114295, B1 => n120642, B2 
                           => n120366, ZN => n6083);
   U84790 : OAI22_X1 port map( A1 => n120374, A2 => n114294, B1 => n120645, B2 
                           => n120366, ZN => n6084);
   U84791 : OAI22_X1 port map( A1 => n120374, A2 => n114293, B1 => n120648, B2 
                           => n120366, ZN => n6085);
   U84792 : OAI22_X1 port map( A1 => n120374, A2 => n114292, B1 => n120651, B2 
                           => n120366, ZN => n6086);
   U84793 : OAI22_X1 port map( A1 => n120374, A2 => n114291, B1 => n120654, B2 
                           => n120366, ZN => n6087);
   U84794 : OAI22_X1 port map( A1 => n120374, A2 => n114290, B1 => n120657, B2 
                           => n120366, ZN => n6088);
   U84795 : OAI22_X1 port map( A1 => n120374, A2 => n114289, B1 => n120660, B2 
                           => n120366, ZN => n6089);
   U84796 : OAI22_X1 port map( A1 => n120374, A2 => n114288, B1 => n120663, B2 
                           => n120366, ZN => n6090);
   U84797 : OAI22_X1 port map( A1 => n120375, A2 => n114287, B1 => n120666, B2 
                           => n120367, ZN => n6091);
   U84798 : OAI22_X1 port map( A1 => n120375, A2 => n114286, B1 => n120669, B2 
                           => n120367, ZN => n6092);
   U84799 : OAI22_X1 port map( A1 => n120375, A2 => n114285, B1 => n120672, B2 
                           => n120367, ZN => n6093);
   U84800 : OAI22_X1 port map( A1 => n120375, A2 => n114284, B1 => n120675, B2 
                           => n120367, ZN => n6094);
   U84801 : OAI22_X1 port map( A1 => n120375, A2 => n114283, B1 => n120678, B2 
                           => n120367, ZN => n6095);
   U84802 : OAI22_X1 port map( A1 => n120375, A2 => n114282, B1 => n120681, B2 
                           => n120367, ZN => n6096);
   U84803 : OAI22_X1 port map( A1 => n120375, A2 => n114281, B1 => n120684, B2 
                           => n120367, ZN => n6097);
   U84804 : OAI22_X1 port map( A1 => n120375, A2 => n114280, B1 => n120687, B2 
                           => n120367, ZN => n6098);
   U84805 : OAI22_X1 port map( A1 => n120375, A2 => n114279, B1 => n120690, B2 
                           => n120367, ZN => n6099);
   U84806 : OAI22_X1 port map( A1 => n120375, A2 => n114278, B1 => n120693, B2 
                           => n120367, ZN => n6100);
   U84807 : OAI22_X1 port map( A1 => n120375, A2 => n114277, B1 => n120696, B2 
                           => n120367, ZN => n6101);
   U84808 : OAI22_X1 port map( A1 => n120375, A2 => n114276, B1 => n120699, B2 
                           => n120367, ZN => n6102);
   U84809 : OAI22_X1 port map( A1 => n120375, A2 => n114275, B1 => n120702, B2 
                           => n120368, ZN => n6103);
   U84810 : OAI22_X1 port map( A1 => n120376, A2 => n114274, B1 => n120705, B2 
                           => n120368, ZN => n6104);
   U84811 : OAI22_X1 port map( A1 => n120376, A2 => n114273, B1 => n120708, B2 
                           => n120368, ZN => n6105);
   U84812 : OAI22_X1 port map( A1 => n120376, A2 => n114272, B1 => n120711, B2 
                           => n120368, ZN => n6106);
   U84813 : OAI22_X1 port map( A1 => n120376, A2 => n114271, B1 => n120714, B2 
                           => n120368, ZN => n6107);
   U84814 : OAI22_X1 port map( A1 => n120376, A2 => n114270, B1 => n120717, B2 
                           => n120368, ZN => n6108);
   U84815 : OAI22_X1 port map( A1 => n120376, A2 => n114269, B1 => n120720, B2 
                           => n120368, ZN => n6109);
   U84816 : OAI22_X1 port map( A1 => n120376, A2 => n114268, B1 => n120723, B2 
                           => n120368, ZN => n6110);
   U84817 : OAI22_X1 port map( A1 => n120376, A2 => n114267, B1 => n120726, B2 
                           => n120368, ZN => n6111);
   U84818 : OAI22_X1 port map( A1 => n120376, A2 => n114266, B1 => n120729, B2 
                           => n120368, ZN => n6112);
   U84819 : OAI22_X1 port map( A1 => n120376, A2 => n114265, B1 => n120732, B2 
                           => n120368, ZN => n6113);
   U84820 : OAI22_X1 port map( A1 => n120376, A2 => n114264, B1 => n120735, B2 
                           => n120368, ZN => n6114);
   U84821 : OAI22_X1 port map( A1 => n120376, A2 => n114263, B1 => n120738, B2 
                           => n120369, ZN => n6115);
   U84822 : OAI22_X1 port map( A1 => n120376, A2 => n114262, B1 => n120741, B2 
                           => n120369, ZN => n6116);
   U84823 : OAI22_X1 port map( A1 => n120377, A2 => n114261, B1 => n120744, B2 
                           => n120369, ZN => n6117);
   U84824 : OAI22_X1 port map( A1 => n120377, A2 => n114260, B1 => n120747, B2 
                           => n120369, ZN => n6118);
   U84825 : OAI22_X1 port map( A1 => n120377, A2 => n114259, B1 => n120750, B2 
                           => n120369, ZN => n6119);
   U84826 : OAI22_X1 port map( A1 => n120377, A2 => n114258, B1 => n120753, B2 
                           => n120369, ZN => n6120);
   U84827 : OAI22_X1 port map( A1 => n120377, A2 => n114257, B1 => n120756, B2 
                           => n120369, ZN => n6121);
   U84828 : OAI22_X1 port map( A1 => n120377, A2 => n114256, B1 => n120759, B2 
                           => n120369, ZN => n6122);
   U84829 : OAI22_X1 port map( A1 => n120377, A2 => n114255, B1 => n120762, B2 
                           => n120369, ZN => n6123);
   U84830 : OAI22_X1 port map( A1 => n120377, A2 => n114254, B1 => n120765, B2 
                           => n120369, ZN => n6124);
   U84831 : OAI22_X1 port map( A1 => n120377, A2 => n114253, B1 => n120768, B2 
                           => n120369, ZN => n6125);
   U84832 : OAI22_X1 port map( A1 => n120377, A2 => n114252, B1 => n120771, B2 
                           => n120369, ZN => n6126);
   U84833 : OAI22_X1 port map( A1 => n120377, A2 => n114251, B1 => n120774, B2 
                           => n120370, ZN => n6127);
   U84834 : OAI22_X1 port map( A1 => n120377, A2 => n114250, B1 => n120777, B2 
                           => n120370, ZN => n6128);
   U84835 : OAI22_X1 port map( A1 => n120377, A2 => n114249, B1 => n120780, B2 
                           => n120370, ZN => n6129);
   U84836 : OAI22_X1 port map( A1 => n120378, A2 => n114248, B1 => n120783, B2 
                           => n120370, ZN => n6130);
   U84837 : OAI22_X1 port map( A1 => n120378, A2 => n114247, B1 => n120786, B2 
                           => n120370, ZN => n6131);
   U84838 : OAI22_X1 port map( A1 => n120378, A2 => n114246, B1 => n120789, B2 
                           => n120370, ZN => n6132);
   U84839 : OAI22_X1 port map( A1 => n120378, A2 => n114245, B1 => n120792, B2 
                           => n120370, ZN => n6133);
   U84840 : OAI22_X1 port map( A1 => n120378, A2 => n114244, B1 => n120795, B2 
                           => n120370, ZN => n6134);
   U84841 : OAI22_X1 port map( A1 => n120378, A2 => n114243, B1 => n120798, B2 
                           => n120370, ZN => n6135);
   U84842 : OAI22_X1 port map( A1 => n120378, A2 => n114242, B1 => n120801, B2 
                           => n120370, ZN => n6136);
   U84843 : OAI22_X1 port map( A1 => n120378, A2 => n114241, B1 => n120804, B2 
                           => n120370, ZN => n6137);
   U84844 : OAI22_X1 port map( A1 => n120378, A2 => n114240, B1 => n120807, B2 
                           => n120370, ZN => n6138);
   U84845 : OAI22_X1 port map( A1 => n120411, A2 => n114210, B1 => n120630, B2 
                           => n120403, ZN => n6271);
   U84846 : OAI22_X1 port map( A1 => n120411, A2 => n114209, B1 => n120633, B2 
                           => n120403, ZN => n6272);
   U84847 : OAI22_X1 port map( A1 => n120411, A2 => n114208, B1 => n120636, B2 
                           => n120403, ZN => n6273);
   U84848 : OAI22_X1 port map( A1 => n120411, A2 => n114207, B1 => n120639, B2 
                           => n120403, ZN => n6274);
   U84849 : OAI22_X1 port map( A1 => n120411, A2 => n114206, B1 => n120642, B2 
                           => n120403, ZN => n6275);
   U84850 : OAI22_X1 port map( A1 => n120411, A2 => n114205, B1 => n120645, B2 
                           => n120403, ZN => n6276);
   U84851 : OAI22_X1 port map( A1 => n120411, A2 => n114204, B1 => n120648, B2 
                           => n120403, ZN => n6277);
   U84852 : OAI22_X1 port map( A1 => n120411, A2 => n114203, B1 => n120651, B2 
                           => n120403, ZN => n6278);
   U84853 : OAI22_X1 port map( A1 => n120411, A2 => n114202, B1 => n120654, B2 
                           => n120403, ZN => n6279);
   U84854 : OAI22_X1 port map( A1 => n120411, A2 => n114201, B1 => n120657, B2 
                           => n120403, ZN => n6280);
   U84855 : OAI22_X1 port map( A1 => n120411, A2 => n114200, B1 => n120660, B2 
                           => n120403, ZN => n6281);
   U84856 : OAI22_X1 port map( A1 => n120411, A2 => n114199, B1 => n120663, B2 
                           => n120403, ZN => n6282);
   U84857 : OAI22_X1 port map( A1 => n120412, A2 => n114198, B1 => n120666, B2 
                           => n120404, ZN => n6283);
   U84858 : OAI22_X1 port map( A1 => n120412, A2 => n114197, B1 => n120669, B2 
                           => n120404, ZN => n6284);
   U84859 : OAI22_X1 port map( A1 => n120412, A2 => n114196, B1 => n120672, B2 
                           => n120404, ZN => n6285);
   U84860 : OAI22_X1 port map( A1 => n120412, A2 => n114195, B1 => n120675, B2 
                           => n120404, ZN => n6286);
   U84861 : OAI22_X1 port map( A1 => n120412, A2 => n114194, B1 => n120678, B2 
                           => n120404, ZN => n6287);
   U84862 : OAI22_X1 port map( A1 => n120412, A2 => n114193, B1 => n120681, B2 
                           => n120404, ZN => n6288);
   U84863 : OAI22_X1 port map( A1 => n120412, A2 => n114192, B1 => n120684, B2 
                           => n120404, ZN => n6289);
   U84864 : OAI22_X1 port map( A1 => n120412, A2 => n114191, B1 => n120687, B2 
                           => n120404, ZN => n6290);
   U84865 : OAI22_X1 port map( A1 => n120412, A2 => n114190, B1 => n120690, B2 
                           => n120404, ZN => n6291);
   U84866 : OAI22_X1 port map( A1 => n120412, A2 => n114189, B1 => n120693, B2 
                           => n120404, ZN => n6292);
   U84867 : OAI22_X1 port map( A1 => n120412, A2 => n114188, B1 => n120696, B2 
                           => n120404, ZN => n6293);
   U84868 : OAI22_X1 port map( A1 => n120412, A2 => n114187, B1 => n120699, B2 
                           => n120404, ZN => n6294);
   U84869 : OAI22_X1 port map( A1 => n120412, A2 => n114186, B1 => n120702, B2 
                           => n120405, ZN => n6295);
   U84870 : OAI22_X1 port map( A1 => n120413, A2 => n114185, B1 => n120705, B2 
                           => n120405, ZN => n6296);
   U84871 : OAI22_X1 port map( A1 => n120413, A2 => n114184, B1 => n120708, B2 
                           => n120405, ZN => n6297);
   U84872 : OAI22_X1 port map( A1 => n120413, A2 => n114183, B1 => n120711, B2 
                           => n120405, ZN => n6298);
   U84873 : OAI22_X1 port map( A1 => n120413, A2 => n114182, B1 => n120714, B2 
                           => n120405, ZN => n6299);
   U84874 : OAI22_X1 port map( A1 => n120413, A2 => n114181, B1 => n120717, B2 
                           => n120405, ZN => n6300);
   U84875 : OAI22_X1 port map( A1 => n120413, A2 => n114180, B1 => n120720, B2 
                           => n120405, ZN => n6301);
   U84876 : OAI22_X1 port map( A1 => n120413, A2 => n114179, B1 => n120723, B2 
                           => n120405, ZN => n6302);
   U84877 : OAI22_X1 port map( A1 => n120413, A2 => n114178, B1 => n120726, B2 
                           => n120405, ZN => n6303);
   U84878 : OAI22_X1 port map( A1 => n120413, A2 => n114177, B1 => n120729, B2 
                           => n120405, ZN => n6304);
   U84879 : OAI22_X1 port map( A1 => n120413, A2 => n114176, B1 => n120732, B2 
                           => n120405, ZN => n6305);
   U84880 : OAI22_X1 port map( A1 => n120413, A2 => n114175, B1 => n120735, B2 
                           => n120405, ZN => n6306);
   U84881 : OAI22_X1 port map( A1 => n120413, A2 => n114174, B1 => n120738, B2 
                           => n120406, ZN => n6307);
   U84882 : OAI22_X1 port map( A1 => n120413, A2 => n114173, B1 => n120741, B2 
                           => n120406, ZN => n6308);
   U84883 : OAI22_X1 port map( A1 => n120414, A2 => n114172, B1 => n120744, B2 
                           => n120406, ZN => n6309);
   U84884 : OAI22_X1 port map( A1 => n120414, A2 => n114171, B1 => n120747, B2 
                           => n120406, ZN => n6310);
   U84885 : OAI22_X1 port map( A1 => n120414, A2 => n114170, B1 => n120750, B2 
                           => n120406, ZN => n6311);
   U84886 : OAI22_X1 port map( A1 => n120414, A2 => n114169, B1 => n120753, B2 
                           => n120406, ZN => n6312);
   U84887 : OAI22_X1 port map( A1 => n120414, A2 => n114168, B1 => n120756, B2 
                           => n120406, ZN => n6313);
   U84888 : OAI22_X1 port map( A1 => n120414, A2 => n114167, B1 => n120759, B2 
                           => n120406, ZN => n6314);
   U84889 : OAI22_X1 port map( A1 => n120414, A2 => n114166, B1 => n120762, B2 
                           => n120406, ZN => n6315);
   U84890 : OAI22_X1 port map( A1 => n120414, A2 => n114165, B1 => n120765, B2 
                           => n120406, ZN => n6316);
   U84891 : OAI22_X1 port map( A1 => n120414, A2 => n114164, B1 => n120768, B2 
                           => n120406, ZN => n6317);
   U84892 : OAI22_X1 port map( A1 => n120414, A2 => n114163, B1 => n120771, B2 
                           => n120406, ZN => n6318);
   U84893 : OAI22_X1 port map( A1 => n120414, A2 => n114162, B1 => n120774, B2 
                           => n120407, ZN => n6319);
   U84894 : OAI22_X1 port map( A1 => n120414, A2 => n114161, B1 => n120777, B2 
                           => n120407, ZN => n6320);
   U84895 : OAI22_X1 port map( A1 => n120414, A2 => n114160, B1 => n120780, B2 
                           => n120407, ZN => n6321);
   U84896 : OAI22_X1 port map( A1 => n120415, A2 => n114159, B1 => n120783, B2 
                           => n120407, ZN => n6322);
   U84897 : OAI22_X1 port map( A1 => n120415, A2 => n114158, B1 => n120786, B2 
                           => n120407, ZN => n6323);
   U84898 : OAI22_X1 port map( A1 => n120415, A2 => n114157, B1 => n120789, B2 
                           => n120407, ZN => n6324);
   U84899 : OAI22_X1 port map( A1 => n120415, A2 => n114156, B1 => n120792, B2 
                           => n120407, ZN => n6325);
   U84900 : OAI22_X1 port map( A1 => n120415, A2 => n114155, B1 => n120795, B2 
                           => n120407, ZN => n6326);
   U84901 : OAI22_X1 port map( A1 => n120415, A2 => n114154, B1 => n120798, B2 
                           => n120407, ZN => n6327);
   U84902 : OAI22_X1 port map( A1 => n120415, A2 => n114153, B1 => n120801, B2 
                           => n120407, ZN => n6328);
   U84903 : OAI22_X1 port map( A1 => n120415, A2 => n114152, B1 => n120804, B2 
                           => n120407, ZN => n6329);
   U84904 : OAI22_X1 port map( A1 => n120415, A2 => n114151, B1 => n120807, B2 
                           => n120407, ZN => n6330);
   U84905 : OAI21_X1 port map( B1 => n113901, B2 => n113913, A => n120623, ZN 
                           => n113914);
   U84906 : OAI21_X1 port map( B1 => n113901, B2 => n113986, A => n120623, ZN 
                           => n113990);
   U84907 : BUF_X1 port map( A => n113891, Z => n120631);
   U84908 : BUF_X1 port map( A => n113889, Z => n120634);
   U84909 : BUF_X1 port map( A => n113887, Z => n120637);
   U84910 : BUF_X1 port map( A => n113885, Z => n120640);
   U84911 : BUF_X1 port map( A => n113883, Z => n120643);
   U84912 : BUF_X1 port map( A => n113881, Z => n120646);
   U84913 : BUF_X1 port map( A => n113879, Z => n120649);
   U84914 : BUF_X1 port map( A => n113877, Z => n120652);
   U84915 : BUF_X1 port map( A => n113875, Z => n120655);
   U84916 : BUF_X1 port map( A => n113873, Z => n120658);
   U84917 : BUF_X1 port map( A => n113871, Z => n120661);
   U84918 : BUF_X1 port map( A => n113869, Z => n120664);
   U84919 : BUF_X1 port map( A => n113867, Z => n120667);
   U84920 : BUF_X1 port map( A => n113865, Z => n120670);
   U84921 : BUF_X1 port map( A => n113863, Z => n120673);
   U84922 : BUF_X1 port map( A => n113861, Z => n120676);
   U84923 : BUF_X1 port map( A => n113859, Z => n120679);
   U84924 : BUF_X1 port map( A => n113857, Z => n120682);
   U84925 : BUF_X1 port map( A => n113855, Z => n120685);
   U84926 : BUF_X1 port map( A => n113853, Z => n120688);
   U84927 : BUF_X1 port map( A => n113851, Z => n120691);
   U84928 : BUF_X1 port map( A => n113849, Z => n120694);
   U84929 : BUF_X1 port map( A => n113847, Z => n120697);
   U84930 : BUF_X1 port map( A => n113845, Z => n120700);
   U84931 : BUF_X1 port map( A => n113843, Z => n120703);
   U84932 : BUF_X1 port map( A => n113841, Z => n120706);
   U84933 : BUF_X1 port map( A => n113839, Z => n120709);
   U84934 : BUF_X1 port map( A => n113837, Z => n120712);
   U84935 : BUF_X1 port map( A => n113835, Z => n120715);
   U84936 : BUF_X1 port map( A => n113833, Z => n120718);
   U84937 : BUF_X1 port map( A => n113831, Z => n120721);
   U84938 : BUF_X1 port map( A => n113829, Z => n120724);
   U84939 : BUF_X1 port map( A => n113827, Z => n120727);
   U84940 : BUF_X1 port map( A => n113825, Z => n120730);
   U84941 : BUF_X1 port map( A => n113823, Z => n120733);
   U84942 : BUF_X1 port map( A => n113821, Z => n120736);
   U84943 : BUF_X1 port map( A => n113819, Z => n120739);
   U84944 : BUF_X1 port map( A => n113817, Z => n120742);
   U84945 : BUF_X1 port map( A => n113815, Z => n120745);
   U84946 : BUF_X1 port map( A => n113813, Z => n120748);
   U84947 : BUF_X1 port map( A => n113811, Z => n120751);
   U84948 : BUF_X1 port map( A => n113809, Z => n120754);
   U84949 : BUF_X1 port map( A => n113807, Z => n120757);
   U84950 : BUF_X1 port map( A => n113805, Z => n120760);
   U84951 : BUF_X1 port map( A => n113803, Z => n120763);
   U84952 : BUF_X1 port map( A => n113801, Z => n120766);
   U84953 : BUF_X1 port map( A => n113799, Z => n120769);
   U84954 : BUF_X1 port map( A => n113797, Z => n120772);
   U84955 : BUF_X1 port map( A => n113795, Z => n120775);
   U84956 : BUF_X1 port map( A => n113793, Z => n120778);
   U84957 : BUF_X1 port map( A => n113791, Z => n120781);
   U84958 : BUF_X1 port map( A => n113789, Z => n120784);
   U84959 : BUF_X1 port map( A => n113787, Z => n120787);
   U84960 : BUF_X1 port map( A => n113785, Z => n120790);
   U84961 : BUF_X1 port map( A => n113783, Z => n120793);
   U84962 : BUF_X1 port map( A => n113781, Z => n120796);
   U84963 : BUF_X1 port map( A => n113779, Z => n120799);
   U84964 : BUF_X1 port map( A => n113777, Z => n120802);
   U84965 : BUF_X1 port map( A => n113775, Z => n120805);
   U84966 : BUF_X1 port map( A => n113771, Z => n120811);
   U84967 : BUF_X1 port map( A => n113770, Z => n120814);
   U84968 : BUF_X1 port map( A => n113769, Z => n120817);
   U84969 : BUF_X1 port map( A => n113768, Z => n120820);
   U84970 : BUF_X1 port map( A => n113773, Z => n120808);
   U84971 : OAI21_X1 port map( B1 => n113986, B2 => n114374, A => n120624, ZN 
                           => n114643);
   U84972 : OAI21_X1 port map( B1 => n113908, B2 => n114141, A => n120624, ZN 
                           => n114145);
   U84973 : OAI21_X1 port map( B1 => n113908, B2 => n114374, A => n120625, ZN 
                           => n114443);
   U84974 : OAI21_X1 port map( B1 => n113894, B2 => n114121, A => n120623, ZN 
                           => n114055);
   U84975 : OAI21_X1 port map( B1 => n113913, B2 => n114144, A => n120624, ZN 
                           => n114234);
   U84976 : OAI21_X1 port map( B1 => n113894, B2 => n114371, A => n120625, ZN 
                           => n114305);
   U84977 : OAI21_X1 port map( B1 => n113913, B2 => n114371, A => n120625, ZN 
                           => n114509);
   U84978 : OAI21_X1 port map( B1 => n113986, B2 => n114371, A => n120625, ZN 
                           => n114577);
   U84979 : OAI21_X1 port map( B1 => n113908, B2 => n114371, A => n120625, ZN 
                           => n114377);
   U84980 : AND2_X1 port map( A1 => n116453, A2 => n116454, ZN => n114662);
   U84981 : AND2_X1 port map( A1 => n117945, A2 => n117946, ZN => n116490);
   U84982 : AND2_X1 port map( A1 => n117953, A2 => n117959, ZN => n116523);
   U84983 : AND2_X1 port map( A1 => n116445, A2 => n116446, ZN => n114657);
   U84984 : AND2_X1 port map( A1 => n116445, A2 => n116463, ZN => n114676);
   U84985 : AND2_X1 port map( A1 => n116452, A2 => n116457, ZN => n114670);
   U84986 : AND2_X1 port map( A1 => n117955, A2 => n117948, ZN => n116503);
   U84987 : AND2_X1 port map( A1 => n117947, A2 => n117945, ZN => n116502);
   U84988 : AND2_X1 port map( A1 => n117947, A2 => n117953, ZN => n116497);
   U84989 : AND2_X1 port map( A1 => n117962, A2 => n117953, ZN => n116507);
   U84990 : AND2_X1 port map( A1 => n117947, A2 => n117954, ZN => n116495);
   U84991 : AND2_X1 port map( A1 => n117961, A2 => n117954, ZN => n116508);
   U84992 : AND2_X1 port map( A1 => n116452, A2 => n116447, ZN => n114664);
   U84993 : AND2_X1 port map( A1 => n116464, A2 => n116447, ZN => n114675);
   U84994 : AND2_X1 port map( A1 => n117955, A2 => n117954, ZN => n116529);
   U84995 : AND2_X1 port map( A1 => n117968, A2 => n117954, ZN => n116522);
   U84996 : AND2_X1 port map( A1 => n116454, A2 => n116447, ZN => n114691);
   U84997 : AND2_X1 port map( A1 => n116459, A2 => n116447, ZN => n114698);
   U84998 : AND2_X1 port map( A1 => n116452, A2 => n116445, ZN => n114669);
   U84999 : AND2_X1 port map( A1 => n116454, A2 => n116445, ZN => n114693);
   U85000 : AND2_X1 port map( A1 => n116458, A2 => n116445, ZN => n114700);
   U85001 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n116471
                           , ZN => n116448);
   U85002 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n117970
                           , ZN => n117959);
   U85003 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n117967
                           , ZN => n117968);
   U85004 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n116470
                           , ZN => n116459);
   U85005 : NOR3_X1 port map( A1 => n117967, A2 => ADD_RD2(4), A3 => n117958, 
                           ZN => n117961);
   U85006 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n116469
                           , ZN => n116446);
   U85007 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n116464);
   U85008 : NOR3_X1 port map( A1 => n117970, A2 => ADD_RD2(3), A3 => n117967, 
                           ZN => n117962);
   U85009 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n117946);
   U85010 : NOR3_X1 port map( A1 => n116470, A2 => ADD_RD1(0), A3 => n116471, 
                           ZN => n116458);
   U85011 : NOR3_X1 port map( A1 => n117970, A2 => ADD_RD2(0), A3 => n117958, 
                           ZN => n117955);
   U85012 : NOR3_X1 port map( A1 => n116469, A2 => ADD_RD1(3), A3 => n116471, 
                           ZN => n116454);
   U85013 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n117958
                           , ZN => n117947);
   U85014 : NOR3_X1 port map( A1 => n116469, A2 => ADD_RD1(4), A3 => n116470, 
                           ZN => n116452);
   U85015 : OAI222_X1 port map( A1 => n113968, A2 => n119904, B1 => n90359, B2 
                           => n119898, C1 => n99364, C2 => n119892, ZN => 
                           n117709);
   U85016 : OAI222_X1 port map( A1 => n113967, A2 => n119905, B1 => n90358, B2 
                           => n119899, C1 => n99363, C2 => n119893, ZN => 
                           n117687);
   U85017 : OAI222_X1 port map( A1 => n113966, A2 => n119905, B1 => n90357, B2 
                           => n119899, C1 => n99362, C2 => n119893, ZN => 
                           n117665);
   U85018 : OAI222_X1 port map( A1 => n113965, A2 => n119905, B1 => n90356, B2 
                           => n119899, C1 => n99361, C2 => n119893, ZN => 
                           n117643);
   U85019 : OAI222_X1 port map( A1 => n113964, A2 => n119905, B1 => n90355, B2 
                           => n119899, C1 => n99360, C2 => n119893, ZN => 
                           n117621);
   U85020 : OAI222_X1 port map( A1 => n113963, A2 => n119905, B1 => n90354, B2 
                           => n119899, C1 => n99359, C2 => n119893, ZN => 
                           n117599);
   U85021 : OAI222_X1 port map( A1 => n113962, A2 => n119905, B1 => n90353, B2 
                           => n119899, C1 => n99358, C2 => n119893, ZN => 
                           n117577);
   U85022 : OAI222_X1 port map( A1 => n113961, A2 => n119905, B1 => n90352, B2 
                           => n119899, C1 => n99357, C2 => n119893, ZN => 
                           n117555);
   U85023 : OAI222_X1 port map( A1 => n113960, A2 => n119905, B1 => n90351, B2 
                           => n119899, C1 => n99356, C2 => n119893, ZN => 
                           n117532);
   U85024 : OAI222_X1 port map( A1 => n113959, A2 => n119905, B1 => n90350, B2 
                           => n119899, C1 => n99355, C2 => n119893, ZN => 
                           n117509);
   U85025 : OAI222_X1 port map( A1 => n113958, A2 => n119905, B1 => n90349, B2 
                           => n119899, C1 => n99354, C2 => n119893, ZN => 
                           n117486);
   U85026 : OAI222_X1 port map( A1 => n113957, A2 => n119905, B1 => n90348, B2 
                           => n119899, C1 => n99353, C2 => n119893, ZN => 
                           n117463);
   U85027 : OAI222_X1 port map( A1 => n113956, A2 => n119905, B1 => n90347, B2 
                           => n119899, C1 => n99352, C2 => n119893, ZN => 
                           n117440);
   U85028 : OAI222_X1 port map( A1 => n113955, A2 => n119906, B1 => n90346, B2 
                           => n119900, C1 => n99351, C2 => n119894, ZN => 
                           n117417);
   U85029 : OAI222_X1 port map( A1 => n113954, A2 => n119906, B1 => n90345, B2 
                           => n119900, C1 => n99350, C2 => n119894, ZN => 
                           n117394);
   U85030 : OAI222_X1 port map( A1 => n113953, A2 => n119906, B1 => n90344, B2 
                           => n119900, C1 => n99349, C2 => n119894, ZN => 
                           n117371);
   U85031 : OAI222_X1 port map( A1 => n113952, A2 => n119906, B1 => n90343, B2 
                           => n119900, C1 => n99348, C2 => n119894, ZN => 
                           n117348);
   U85032 : OAI222_X1 port map( A1 => n113951, A2 => n119906, B1 => n90342, B2 
                           => n119900, C1 => n99347, C2 => n119894, ZN => 
                           n117325);
   U85033 : OAI222_X1 port map( A1 => n113950, A2 => n119906, B1 => n90341, B2 
                           => n119900, C1 => n99346, C2 => n119894, ZN => 
                           n117302);
   U85034 : OAI222_X1 port map( A1 => n113949, A2 => n119906, B1 => n90340, B2 
                           => n119900, C1 => n99345, C2 => n119894, ZN => 
                           n117279);
   U85035 : OAI222_X1 port map( A1 => n113948, A2 => n119906, B1 => n90339, B2 
                           => n119900, C1 => n99344, C2 => n119894, ZN => 
                           n117256);
   U85036 : OAI222_X1 port map( A1 => n113947, A2 => n119906, B1 => n90338, B2 
                           => n119900, C1 => n99343, C2 => n119894, ZN => 
                           n117233);
   U85037 : OAI222_X1 port map( A1 => n113946, A2 => n119906, B1 => n90337, B2 
                           => n119900, C1 => n99342, C2 => n119894, ZN => 
                           n117210);
   U85038 : OAI222_X1 port map( A1 => n113945, A2 => n119906, B1 => n90336, B2 
                           => n119900, C1 => n99341, C2 => n119894, ZN => 
                           n117187);
   U85039 : OAI222_X1 port map( A1 => n113944, A2 => n119906, B1 => n90335, B2 
                           => n119900, C1 => n99340, C2 => n119894, ZN => 
                           n117164);
   U85040 : OAI222_X1 port map( A1 => n113943, A2 => n119907, B1 => n90334, B2 
                           => n119901, C1 => n99339, C2 => n119895, ZN => 
                           n117141);
   U85041 : OAI222_X1 port map( A1 => n113942, A2 => n119907, B1 => n90333, B2 
                           => n119901, C1 => n99338, C2 => n119895, ZN => 
                           n117118);
   U85042 : OAI222_X1 port map( A1 => n113941, A2 => n119907, B1 => n90332, B2 
                           => n119901, C1 => n99337, C2 => n119895, ZN => 
                           n117095);
   U85043 : OAI222_X1 port map( A1 => n113940, A2 => n119907, B1 => n90331, B2 
                           => n119901, C1 => n99336, C2 => n119895, ZN => 
                           n117072);
   U85044 : OAI222_X1 port map( A1 => n113939, A2 => n119907, B1 => n90330, B2 
                           => n119901, C1 => n99335, C2 => n119895, ZN => 
                           n117049);
   U85045 : OAI222_X1 port map( A1 => n113938, A2 => n119907, B1 => n90329, B2 
                           => n119901, C1 => n99334, C2 => n119895, ZN => 
                           n117026);
   U85046 : OAI222_X1 port map( A1 => n113937, A2 => n119907, B1 => n90328, B2 
                           => n119901, C1 => n99333, C2 => n119895, ZN => 
                           n117003);
   U85047 : OAI222_X1 port map( A1 => n113936, A2 => n119907, B1 => n90327, B2 
                           => n119901, C1 => n99332, C2 => n119895, ZN => 
                           n116980);
   U85048 : OAI222_X1 port map( A1 => n113935, A2 => n119907, B1 => n90326, B2 
                           => n119901, C1 => n99331, C2 => n119895, ZN => 
                           n116957);
   U85049 : OAI222_X1 port map( A1 => n113934, A2 => n119907, B1 => n90325, B2 
                           => n119901, C1 => n99330, C2 => n119895, ZN => 
                           n116934);
   U85050 : OAI222_X1 port map( A1 => n113933, A2 => n119907, B1 => n90324, B2 
                           => n119901, C1 => n99329, C2 => n119895, ZN => 
                           n116911);
   U85051 : OAI222_X1 port map( A1 => n113932, A2 => n119907, B1 => n90323, B2 
                           => n119901, C1 => n99328, C2 => n119895, ZN => 
                           n116888);
   U85052 : OAI222_X1 port map( A1 => n113931, A2 => n119908, B1 => n90322, B2 
                           => n119902, C1 => n99327, C2 => n119896, ZN => 
                           n116865);
   U85053 : OAI222_X1 port map( A1 => n113930, A2 => n119908, B1 => n90321, B2 
                           => n119902, C1 => n99326, C2 => n119896, ZN => 
                           n116842);
   U85054 : OAI222_X1 port map( A1 => n113929, A2 => n119908, B1 => n90320, B2 
                           => n119902, C1 => n99325, C2 => n119896, ZN => 
                           n116819);
   U85055 : OAI222_X1 port map( A1 => n113928, A2 => n119908, B1 => n90319, B2 
                           => n119902, C1 => n99324, C2 => n119896, ZN => 
                           n116796);
   U85056 : OAI222_X1 port map( A1 => n113927, A2 => n119908, B1 => n90318, B2 
                           => n119902, C1 => n99323, C2 => n119896, ZN => 
                           n116773);
   U85057 : OAI222_X1 port map( A1 => n113926, A2 => n119908, B1 => n90317, B2 
                           => n119902, C1 => n99322, C2 => n119896, ZN => 
                           n116750);
   U85058 : OAI222_X1 port map( A1 => n113925, A2 => n119908, B1 => n90316, B2 
                           => n119902, C1 => n99321, C2 => n119896, ZN => 
                           n116727);
   U85059 : OAI222_X1 port map( A1 => n113924, A2 => n119908, B1 => n90315, B2 
                           => n119902, C1 => n99320, C2 => n119896, ZN => 
                           n116704);
   U85060 : OAI222_X1 port map( A1 => n113923, A2 => n119908, B1 => n90314, B2 
                           => n119902, C1 => n99319, C2 => n119896, ZN => 
                           n116681);
   U85061 : OAI222_X1 port map( A1 => n113922, A2 => n119908, B1 => n90313, B2 
                           => n119902, C1 => n99318, C2 => n119896, ZN => 
                           n116658);
   U85062 : OAI222_X1 port map( A1 => n113921, A2 => n119908, B1 => n90312, B2 
                           => n119902, C1 => n99317, C2 => n119896, ZN => 
                           n116635);
   U85063 : OAI222_X1 port map( A1 => n113920, A2 => n119908, B1 => n90311, B2 
                           => n119902, C1 => n99316, C2 => n119896, ZN => 
                           n116612);
   U85064 : OAI222_X1 port map( A1 => n99131, A2 => n120105, B1 => n120099, B2 
                           => n115146, C1 => n113933, C2 => n120093, ZN => 
                           n115165);
   U85065 : OAI222_X1 port map( A1 => n99130, A2 => n120105, B1 => n120099, B2 
                           => n115118, C1 => n113932, C2 => n120093, ZN => 
                           n115137);
   U85066 : OAI222_X1 port map( A1 => n99129, A2 => n120106, B1 => n120100, B2 
                           => n115090, C1 => n113931, C2 => n120094, ZN => 
                           n115109);
   U85067 : OAI222_X1 port map( A1 => n99128, A2 => n120106, B1 => n120100, B2 
                           => n115062, C1 => n113930, C2 => n120094, ZN => 
                           n115081);
   U85068 : OAI222_X1 port map( A1 => n99127, A2 => n120106, B1 => n120100, B2 
                           => n115034, C1 => n113929, C2 => n120094, ZN => 
                           n115053);
   U85069 : OAI222_X1 port map( A1 => n99126, A2 => n120106, B1 => n120100, B2 
                           => n115006, C1 => n113928, C2 => n120094, ZN => 
                           n115025);
   U85070 : OAI222_X1 port map( A1 => n99125, A2 => n120106, B1 => n120100, B2 
                           => n114978, C1 => n113927, C2 => n120094, ZN => 
                           n114997);
   U85071 : OAI222_X1 port map( A1 => n99124, A2 => n120106, B1 => n120100, B2 
                           => n114950, C1 => n113926, C2 => n120094, ZN => 
                           n114969);
   U85072 : OAI222_X1 port map( A1 => n99123, A2 => n120106, B1 => n120100, B2 
                           => n114922, C1 => n113925, C2 => n120094, ZN => 
                           n114941);
   U85073 : OAI222_X1 port map( A1 => n99122, A2 => n120106, B1 => n120100, B2 
                           => n114894, C1 => n113924, C2 => n120094, ZN => 
                           n114913);
   U85074 : OAI222_X1 port map( A1 => n99121, A2 => n120106, B1 => n120100, B2 
                           => n114866, C1 => n113923, C2 => n120094, ZN => 
                           n114885);
   U85075 : OAI222_X1 port map( A1 => n99120, A2 => n120106, B1 => n120100, B2 
                           => n114838, C1 => n113922, C2 => n120094, ZN => 
                           n114857);
   U85076 : OAI222_X1 port map( A1 => n99119, A2 => n120106, B1 => n120100, B2 
                           => n114810, C1 => n113921, C2 => n120094, ZN => 
                           n114829);
   U85077 : OAI222_X1 port map( A1 => n99118, A2 => n120106, B1 => n120100, B2 
                           => n114782, C1 => n113920, C2 => n120094, ZN => 
                           n114801);
   U85078 : OAI222_X1 port map( A1 => n99177, A2 => n120102, B1 => n120096, B2 
                           => n116434, C1 => n113979, C2 => n120090, ZN => 
                           n116465);
   U85079 : OAI222_X1 port map( A1 => n99176, A2 => n120102, B1 => n120096, B2 
                           => n116406, C1 => n113978, C2 => n120090, ZN => 
                           n116425);
   U85080 : OAI222_X1 port map( A1 => n99175, A2 => n120102, B1 => n120096, B2 
                           => n116378, C1 => n113977, C2 => n120090, ZN => 
                           n116397);
   U85081 : OAI222_X1 port map( A1 => n99174, A2 => n120102, B1 => n120096, B2 
                           => n116350, C1 => n113976, C2 => n120090, ZN => 
                           n116369);
   U85082 : OAI222_X1 port map( A1 => n113972, A2 => n119904, B1 => n90363, B2 
                           => n119898, C1 => n99368, C2 => n119892, ZN => 
                           n117797);
   U85083 : OAI222_X1 port map( A1 => n113971, A2 => n119904, B1 => n90362, B2 
                           => n119898, C1 => n99367, C2 => n119892, ZN => 
                           n117775);
   U85084 : OAI222_X1 port map( A1 => n113970, A2 => n119904, B1 => n90361, B2 
                           => n119898, C1 => n99366, C2 => n119892, ZN => 
                           n117753);
   U85085 : OAI222_X1 port map( A1 => n113969, A2 => n119904, B1 => n90360, B2 
                           => n119898, C1 => n99365, C2 => n119892, ZN => 
                           n117731);
   U85086 : OAI222_X1 port map( A1 => n113979, A2 => n119904, B1 => n90370, B2 
                           => n119898, C1 => n99375, C2 => n119892, ZN => 
                           n117963);
   U85087 : OAI222_X1 port map( A1 => n113978, A2 => n119904, B1 => n90369, B2 
                           => n119898, C1 => n99374, C2 => n119892, ZN => 
                           n117929);
   U85088 : OAI222_X1 port map( A1 => n113977, A2 => n119904, B1 => n90368, B2 
                           => n119898, C1 => n99373, C2 => n119892, ZN => 
                           n117907);
   U85089 : OAI222_X1 port map( A1 => n113976, A2 => n119904, B1 => n90367, B2 
                           => n119898, C1 => n99372, C2 => n119892, ZN => 
                           n117885);
   U85090 : OAI222_X1 port map( A1 => n113975, A2 => n119904, B1 => n90366, B2 
                           => n119898, C1 => n99371, C2 => n119892, ZN => 
                           n117863);
   U85091 : OAI222_X1 port map( A1 => n113974, A2 => n119904, B1 => n90365, B2 
                           => n119898, C1 => n99370, C2 => n119892, ZN => 
                           n117841);
   U85092 : OAI222_X1 port map( A1 => n113973, A2 => n119904, B1 => n90364, B2 
                           => n119898, C1 => n99369, C2 => n119892, ZN => 
                           n117819);
   U85093 : OAI222_X1 port map( A1 => n99173, A2 => n120102, B1 => n120096, B2 
                           => n116322, C1 => n113975, C2 => n120090, ZN => 
                           n116341);
   U85094 : OAI222_X1 port map( A1 => n99172, A2 => n120102, B1 => n120096, B2 
                           => n116294, C1 => n113974, C2 => n120090, ZN => 
                           n116313);
   U85095 : OAI222_X1 port map( A1 => n99171, A2 => n120102, B1 => n120096, B2 
                           => n116266, C1 => n113973, C2 => n120090, ZN => 
                           n116285);
   U85096 : OAI222_X1 port map( A1 => n99170, A2 => n120102, B1 => n120096, B2 
                           => n116238, C1 => n113972, C2 => n120090, ZN => 
                           n116257);
   U85097 : OAI222_X1 port map( A1 => n99169, A2 => n120102, B1 => n120096, B2 
                           => n116210, C1 => n113971, C2 => n120090, ZN => 
                           n116229);
   U85098 : OAI222_X1 port map( A1 => n99168, A2 => n120102, B1 => n120096, B2 
                           => n116182, C1 => n113970, C2 => n120090, ZN => 
                           n116201);
   U85099 : OAI222_X1 port map( A1 => n99167, A2 => n120102, B1 => n120096, B2 
                           => n116154, C1 => n113969, C2 => n120090, ZN => 
                           n116173);
   U85100 : OAI222_X1 port map( A1 => n99166, A2 => n120102, B1 => n120096, B2 
                           => n116126, C1 => n113968, C2 => n120090, ZN => 
                           n116145);
   U85101 : OAI222_X1 port map( A1 => n99165, A2 => n120103, B1 => n120097, B2 
                           => n116098, C1 => n113967, C2 => n120091, ZN => 
                           n116117);
   U85102 : OAI222_X1 port map( A1 => n99164, A2 => n120103, B1 => n120097, B2 
                           => n116070, C1 => n113966, C2 => n120091, ZN => 
                           n116089);
   U85103 : OAI222_X1 port map( A1 => n99163, A2 => n120103, B1 => n120097, B2 
                           => n116042, C1 => n113965, C2 => n120091, ZN => 
                           n116061);
   U85104 : OAI222_X1 port map( A1 => n99162, A2 => n120103, B1 => n120097, B2 
                           => n116014, C1 => n113964, C2 => n120091, ZN => 
                           n116033);
   U85105 : OAI222_X1 port map( A1 => n99161, A2 => n120103, B1 => n120097, B2 
                           => n115986, C1 => n113963, C2 => n120091, ZN => 
                           n116005);
   U85106 : OAI222_X1 port map( A1 => n99160, A2 => n120103, B1 => n120097, B2 
                           => n115958, C1 => n113962, C2 => n120091, ZN => 
                           n115977);
   U85107 : OAI222_X1 port map( A1 => n99159, A2 => n120103, B1 => n120097, B2 
                           => n115930, C1 => n113961, C2 => n120091, ZN => 
                           n115949);
   U85108 : OAI222_X1 port map( A1 => n99158, A2 => n120103, B1 => n120097, B2 
                           => n115902, C1 => n113960, C2 => n120091, ZN => 
                           n115921);
   U85109 : OAI222_X1 port map( A1 => n99157, A2 => n120103, B1 => n120097, B2 
                           => n115874, C1 => n113959, C2 => n120091, ZN => 
                           n115893);
   U85110 : OAI222_X1 port map( A1 => n99156, A2 => n120103, B1 => n120097, B2 
                           => n115846, C1 => n113958, C2 => n120091, ZN => 
                           n115865);
   U85111 : OAI222_X1 port map( A1 => n99155, A2 => n120103, B1 => n120097, B2 
                           => n115818, C1 => n113957, C2 => n120091, ZN => 
                           n115837);
   U85112 : OAI222_X1 port map( A1 => n99154, A2 => n120103, B1 => n120097, B2 
                           => n115790, C1 => n113956, C2 => n120091, ZN => 
                           n115809);
   U85113 : OAI222_X1 port map( A1 => n99153, A2 => n120104, B1 => n120098, B2 
                           => n115762, C1 => n113955, C2 => n120092, ZN => 
                           n115781);
   U85114 : OAI222_X1 port map( A1 => n99152, A2 => n120104, B1 => n120098, B2 
                           => n115734, C1 => n113954, C2 => n120092, ZN => 
                           n115753);
   U85115 : OAI222_X1 port map( A1 => n99151, A2 => n120104, B1 => n120098, B2 
                           => n115706, C1 => n113953, C2 => n120092, ZN => 
                           n115725);
   U85116 : OAI222_X1 port map( A1 => n99150, A2 => n120104, B1 => n120098, B2 
                           => n115678, C1 => n113952, C2 => n120092, ZN => 
                           n115697);
   U85117 : OAI222_X1 port map( A1 => n99149, A2 => n120104, B1 => n120098, B2 
                           => n115650, C1 => n113951, C2 => n120092, ZN => 
                           n115669);
   U85118 : OAI222_X1 port map( A1 => n99148, A2 => n120104, B1 => n120098, B2 
                           => n115622, C1 => n113950, C2 => n120092, ZN => 
                           n115641);
   U85119 : OAI222_X1 port map( A1 => n99147, A2 => n120104, B1 => n120098, B2 
                           => n115594, C1 => n113949, C2 => n120092, ZN => 
                           n115613);
   U85120 : OAI222_X1 port map( A1 => n99146, A2 => n120104, B1 => n120098, B2 
                           => n115566, C1 => n113948, C2 => n120092, ZN => 
                           n115585);
   U85121 : OAI222_X1 port map( A1 => n99145, A2 => n120104, B1 => n120098, B2 
                           => n115538, C1 => n113947, C2 => n120092, ZN => 
                           n115557);
   U85122 : OAI222_X1 port map( A1 => n99144, A2 => n120104, B1 => n120098, B2 
                           => n115510, C1 => n113946, C2 => n120092, ZN => 
                           n115529);
   U85123 : OAI222_X1 port map( A1 => n99143, A2 => n120104, B1 => n120098, B2 
                           => n115482, C1 => n113945, C2 => n120092, ZN => 
                           n115501);
   U85124 : OAI222_X1 port map( A1 => n99142, A2 => n120104, B1 => n120098, B2 
                           => n115454, C1 => n113944, C2 => n120092, ZN => 
                           n115473);
   U85125 : OAI222_X1 port map( A1 => n99141, A2 => n120105, B1 => n120099, B2 
                           => n115426, C1 => n113943, C2 => n120093, ZN => 
                           n115445);
   U85126 : OAI222_X1 port map( A1 => n99140, A2 => n120105, B1 => n120099, B2 
                           => n115398, C1 => n113942, C2 => n120093, ZN => 
                           n115417);
   U85127 : OAI222_X1 port map( A1 => n99139, A2 => n120105, B1 => n120099, B2 
                           => n115370, C1 => n113941, C2 => n120093, ZN => 
                           n115389);
   U85128 : OAI222_X1 port map( A1 => n99138, A2 => n120105, B1 => n120099, B2 
                           => n115342, C1 => n113940, C2 => n120093, ZN => 
                           n115361);
   U85129 : OAI222_X1 port map( A1 => n99137, A2 => n120105, B1 => n120099, B2 
                           => n115314, C1 => n113939, C2 => n120093, ZN => 
                           n115333);
   U85130 : OAI222_X1 port map( A1 => n99136, A2 => n120105, B1 => n120099, B2 
                           => n115286, C1 => n113938, C2 => n120093, ZN => 
                           n115305);
   U85131 : OAI222_X1 port map( A1 => n99135, A2 => n120105, B1 => n120099, B2 
                           => n115258, C1 => n113937, C2 => n120093, ZN => 
                           n115277);
   U85132 : OAI222_X1 port map( A1 => n99134, A2 => n120105, B1 => n120099, B2 
                           => n115230, C1 => n113936, C2 => n120093, ZN => 
                           n115249);
   U85133 : OAI222_X1 port map( A1 => n99133, A2 => n120105, B1 => n120099, B2 
                           => n115202, C1 => n113935, C2 => n120093, ZN => 
                           n115221);
   U85134 : OAI222_X1 port map( A1 => n99132, A2 => n120105, B1 => n120099, B2 
                           => n115174, C1 => n113934, C2 => n120093, ZN => 
                           n115193);
   U85135 : OAI222_X1 port map( A1 => n99117, A2 => n120107, B1 => n120101, B2 
                           => n114756, C1 => n113919, C2 => n120095, ZN => 
                           n114773);
   U85136 : OAI222_X1 port map( A1 => n99116, A2 => n120107, B1 => n120101, B2 
                           => n114730, C1 => n113918, C2 => n120095, ZN => 
                           n114747);
   U85137 : OAI222_X1 port map( A1 => n99115, A2 => n120107, B1 => n120101, B2 
                           => n114704, C1 => n113917, C2 => n120095, ZN => 
                           n114721);
   U85138 : OAI222_X1 port map( A1 => n99113, A2 => n120107, B1 => n114644, B2 
                           => n120101, C1 => n113915, C2 => n120095, ZN => 
                           n114678);
   U85139 : OAI222_X1 port map( A1 => n113919, A2 => n119909, B1 => n90310, B2 
                           => n119903, C1 => n99315, C2 => n119897, ZN => 
                           n116589);
   U85140 : OAI222_X1 port map( A1 => n113918, A2 => n119909, B1 => n90309, B2 
                           => n119903, C1 => n99314, C2 => n119897, ZN => 
                           n116568);
   U85141 : OAI222_X1 port map( A1 => n113917, A2 => n119909, B1 => n90308, B2 
                           => n119903, C1 => n99313, C2 => n119897, ZN => 
                           n116547);
   U85142 : OAI222_X1 port map( A1 => n113915, A2 => n119909, B1 => n90306, B2 
                           => n119903, C1 => n99311, C2 => n119897, ZN => 
                           n116509);
   U85143 : NOR4_X1 port map( A1 => n117697, A2 => n117698, A3 => n117699, A4 
                           => n117700, ZN => n117696);
   U85144 : OAI221_X1 port map( B1 => n99232, B2 => n119964, C1 => n98896, C2 
                           => n119958, A => n117708, ZN => n117697);
   U85145 : OAI221_X1 port map( B1 => n114497, B2 => n120036, C1 => n99298, C2 
                           => n120030, A => n117701, ZN => n117700);
   U85146 : OAI221_X1 port map( B1 => n114563, B2 => n119988, C1 => n114199, C2
                           => n119982, A => n117706, ZN => n117698);
   U85147 : NOR4_X1 port map( A1 => n117675, A2 => n117676, A3 => n117677, A4 
                           => n117678, ZN => n117674);
   U85148 : OAI221_X1 port map( B1 => n99231, B2 => n119965, C1 => n98895, C2 
                           => n119959, A => n117686, ZN => n117675);
   U85149 : OAI221_X1 port map( B1 => n114496, B2 => n120037, C1 => n99297, C2 
                           => n120031, A => n117679, ZN => n117678);
   U85150 : OAI221_X1 port map( B1 => n114562, B2 => n119989, C1 => n114198, C2
                           => n119983, A => n117684, ZN => n117676);
   U85151 : NOR4_X1 port map( A1 => n117653, A2 => n117654, A3 => n117655, A4 
                           => n117656, ZN => n117652);
   U85152 : OAI221_X1 port map( B1 => n99230, B2 => n119965, C1 => n98894, C2 
                           => n119959, A => n117664, ZN => n117653);
   U85153 : OAI221_X1 port map( B1 => n114495, B2 => n120037, C1 => n99296, C2 
                           => n120031, A => n117657, ZN => n117656);
   U85154 : OAI221_X1 port map( B1 => n114561, B2 => n119989, C1 => n114197, C2
                           => n119983, A => n117662, ZN => n117654);
   U85155 : NOR4_X1 port map( A1 => n117631, A2 => n117632, A3 => n117633, A4 
                           => n117634, ZN => n117630);
   U85156 : OAI221_X1 port map( B1 => n99229, B2 => n119965, C1 => n98893, C2 
                           => n119959, A => n117642, ZN => n117631);
   U85157 : OAI221_X1 port map( B1 => n114494, B2 => n120037, C1 => n99295, C2 
                           => n120031, A => n117635, ZN => n117634);
   U85158 : OAI221_X1 port map( B1 => n114560, B2 => n119989, C1 => n114196, C2
                           => n119983, A => n117640, ZN => n117632);
   U85159 : NOR4_X1 port map( A1 => n117609, A2 => n117610, A3 => n117611, A4 
                           => n117612, ZN => n117608);
   U85160 : OAI221_X1 port map( B1 => n99228, B2 => n119965, C1 => n98892, C2 
                           => n119959, A => n117620, ZN => n117609);
   U85161 : OAI221_X1 port map( B1 => n114493, B2 => n120037, C1 => n99294, C2 
                           => n120031, A => n117613, ZN => n117612);
   U85162 : OAI221_X1 port map( B1 => n114559, B2 => n119989, C1 => n114195, C2
                           => n119983, A => n117618, ZN => n117610);
   U85163 : NOR4_X1 port map( A1 => n117587, A2 => n117588, A3 => n117589, A4 
                           => n117590, ZN => n117586);
   U85164 : OAI221_X1 port map( B1 => n99227, B2 => n119965, C1 => n98891, C2 
                           => n119959, A => n117598, ZN => n117587);
   U85165 : OAI221_X1 port map( B1 => n114492, B2 => n120037, C1 => n99293, C2 
                           => n120031, A => n117591, ZN => n117590);
   U85166 : OAI221_X1 port map( B1 => n114558, B2 => n119989, C1 => n114194, C2
                           => n119983, A => n117596, ZN => n117588);
   U85167 : NOR4_X1 port map( A1 => n117565, A2 => n117566, A3 => n117567, A4 
                           => n117568, ZN => n117564);
   U85168 : OAI221_X1 port map( B1 => n99226, B2 => n119965, C1 => n98890, C2 
                           => n119959, A => n117576, ZN => n117565);
   U85169 : OAI221_X1 port map( B1 => n114491, B2 => n120037, C1 => n99292, C2 
                           => n120031, A => n117569, ZN => n117568);
   U85170 : OAI221_X1 port map( B1 => n114557, B2 => n119989, C1 => n114193, C2
                           => n119983, A => n117574, ZN => n117566);
   U85171 : NOR4_X1 port map( A1 => n117543, A2 => n117544, A3 => n117545, A4 
                           => n117546, ZN => n117542);
   U85172 : OAI221_X1 port map( B1 => n99225, B2 => n119965, C1 => n98889, C2 
                           => n119959, A => n117554, ZN => n117543);
   U85173 : OAI221_X1 port map( B1 => n114490, B2 => n120037, C1 => n99291, C2 
                           => n120031, A => n117547, ZN => n117546);
   U85174 : OAI221_X1 port map( B1 => n114556, B2 => n119989, C1 => n114192, C2
                           => n119983, A => n117552, ZN => n117544);
   U85175 : NOR4_X1 port map( A1 => n117520, A2 => n117521, A3 => n117522, A4 
                           => n117523, ZN => n117519);
   U85176 : OAI221_X1 port map( B1 => n99224, B2 => n119965, C1 => n98888, C2 
                           => n119959, A => n117531, ZN => n117520);
   U85177 : OAI221_X1 port map( B1 => n114489, B2 => n120037, C1 => n99290, C2 
                           => n120031, A => n117524, ZN => n117523);
   U85178 : OAI221_X1 port map( B1 => n114555, B2 => n119989, C1 => n114191, C2
                           => n119983, A => n117529, ZN => n117521);
   U85179 : NOR4_X1 port map( A1 => n117497, A2 => n117498, A3 => n117499, A4 
                           => n117500, ZN => n117496);
   U85180 : OAI221_X1 port map( B1 => n99223, B2 => n119965, C1 => n98887, C2 
                           => n119959, A => n117508, ZN => n117497);
   U85181 : OAI221_X1 port map( B1 => n114488, B2 => n120037, C1 => n99289, C2 
                           => n120031, A => n117501, ZN => n117500);
   U85182 : OAI221_X1 port map( B1 => n114554, B2 => n119989, C1 => n114190, C2
                           => n119983, A => n117506, ZN => n117498);
   U85183 : NOR4_X1 port map( A1 => n117474, A2 => n117475, A3 => n117476, A4 
                           => n117477, ZN => n117473);
   U85184 : OAI221_X1 port map( B1 => n99222, B2 => n119965, C1 => n98886, C2 
                           => n119959, A => n117485, ZN => n117474);
   U85185 : OAI221_X1 port map( B1 => n114487, B2 => n120037, C1 => n99288, C2 
                           => n120031, A => n117478, ZN => n117477);
   U85186 : OAI221_X1 port map( B1 => n114553, B2 => n119989, C1 => n114189, C2
                           => n119983, A => n117483, ZN => n117475);
   U85187 : NOR4_X1 port map( A1 => n117451, A2 => n117452, A3 => n117453, A4 
                           => n117454, ZN => n117450);
   U85188 : OAI221_X1 port map( B1 => n99221, B2 => n119965, C1 => n98885, C2 
                           => n119959, A => n117462, ZN => n117451);
   U85189 : OAI221_X1 port map( B1 => n114486, B2 => n120037, C1 => n99287, C2 
                           => n120031, A => n117455, ZN => n117454);
   U85190 : OAI221_X1 port map( B1 => n114552, B2 => n119989, C1 => n114188, C2
                           => n119983, A => n117460, ZN => n117452);
   U85191 : NOR4_X1 port map( A1 => n117428, A2 => n117429, A3 => n117430, A4 
                           => n117431, ZN => n117427);
   U85192 : OAI221_X1 port map( B1 => n99220, B2 => n119965, C1 => n98884, C2 
                           => n119959, A => n117439, ZN => n117428);
   U85193 : OAI221_X1 port map( B1 => n114485, B2 => n120037, C1 => n99286, C2 
                           => n120031, A => n117432, ZN => n117431);
   U85194 : OAI221_X1 port map( B1 => n114551, B2 => n119989, C1 => n114187, C2
                           => n119983, A => n117437, ZN => n117429);
   U85195 : NOR4_X1 port map( A1 => n117405, A2 => n117406, A3 => n117407, A4 
                           => n117408, ZN => n117404);
   U85196 : OAI221_X1 port map( B1 => n99219, B2 => n119966, C1 => n98883, C2 
                           => n119960, A => n117416, ZN => n117405);
   U85197 : OAI221_X1 port map( B1 => n114484, B2 => n120038, C1 => n99285, C2 
                           => n120032, A => n117409, ZN => n117408);
   U85198 : OAI221_X1 port map( B1 => n114550, B2 => n119990, C1 => n114186, C2
                           => n119984, A => n117414, ZN => n117406);
   U85199 : NOR4_X1 port map( A1 => n117382, A2 => n117383, A3 => n117384, A4 
                           => n117385, ZN => n117381);
   U85200 : OAI221_X1 port map( B1 => n99218, B2 => n119966, C1 => n98882, C2 
                           => n119960, A => n117393, ZN => n117382);
   U85201 : OAI221_X1 port map( B1 => n114483, B2 => n120038, C1 => n99284, C2 
                           => n120032, A => n117386, ZN => n117385);
   U85202 : OAI221_X1 port map( B1 => n114549, B2 => n119990, C1 => n114185, C2
                           => n119984, A => n117391, ZN => n117383);
   U85203 : NOR4_X1 port map( A1 => n117359, A2 => n117360, A3 => n117361, A4 
                           => n117362, ZN => n117358);
   U85204 : OAI221_X1 port map( B1 => n99217, B2 => n119966, C1 => n98881, C2 
                           => n119960, A => n117370, ZN => n117359);
   U85205 : OAI221_X1 port map( B1 => n114482, B2 => n120038, C1 => n99283, C2 
                           => n120032, A => n117363, ZN => n117362);
   U85206 : OAI221_X1 port map( B1 => n114548, B2 => n119990, C1 => n114184, C2
                           => n119984, A => n117368, ZN => n117360);
   U85207 : NOR4_X1 port map( A1 => n117336, A2 => n117337, A3 => n117338, A4 
                           => n117339, ZN => n117335);
   U85208 : OAI221_X1 port map( B1 => n99216, B2 => n119966, C1 => n98880, C2 
                           => n119960, A => n117347, ZN => n117336);
   U85209 : OAI221_X1 port map( B1 => n114481, B2 => n120038, C1 => n99282, C2 
                           => n120032, A => n117340, ZN => n117339);
   U85210 : OAI221_X1 port map( B1 => n114547, B2 => n119990, C1 => n114183, C2
                           => n119984, A => n117345, ZN => n117337);
   U85211 : NOR4_X1 port map( A1 => n117313, A2 => n117314, A3 => n117315, A4 
                           => n117316, ZN => n117312);
   U85212 : OAI221_X1 port map( B1 => n99215, B2 => n119966, C1 => n98879, C2 
                           => n119960, A => n117324, ZN => n117313);
   U85213 : OAI221_X1 port map( B1 => n114480, B2 => n120038, C1 => n99281, C2 
                           => n120032, A => n117317, ZN => n117316);
   U85214 : OAI221_X1 port map( B1 => n114546, B2 => n119990, C1 => n114182, C2
                           => n119984, A => n117322, ZN => n117314);
   U85215 : NOR4_X1 port map( A1 => n117290, A2 => n117291, A3 => n117292, A4 
                           => n117293, ZN => n117289);
   U85216 : OAI221_X1 port map( B1 => n99214, B2 => n119966, C1 => n98878, C2 
                           => n119960, A => n117301, ZN => n117290);
   U85217 : OAI221_X1 port map( B1 => n114479, B2 => n120038, C1 => n99280, C2 
                           => n120032, A => n117294, ZN => n117293);
   U85218 : OAI221_X1 port map( B1 => n114545, B2 => n119990, C1 => n114181, C2
                           => n119984, A => n117299, ZN => n117291);
   U85219 : NOR4_X1 port map( A1 => n117267, A2 => n117268, A3 => n117269, A4 
                           => n117270, ZN => n117266);
   U85220 : OAI221_X1 port map( B1 => n99213, B2 => n119966, C1 => n98877, C2 
                           => n119960, A => n117278, ZN => n117267);
   U85221 : OAI221_X1 port map( B1 => n114478, B2 => n120038, C1 => n99279, C2 
                           => n120032, A => n117271, ZN => n117270);
   U85222 : OAI221_X1 port map( B1 => n114544, B2 => n119990, C1 => n114180, C2
                           => n119984, A => n117276, ZN => n117268);
   U85223 : NOR4_X1 port map( A1 => n117244, A2 => n117245, A3 => n117246, A4 
                           => n117247, ZN => n117243);
   U85224 : OAI221_X1 port map( B1 => n99212, B2 => n119966, C1 => n98876, C2 
                           => n119960, A => n117255, ZN => n117244);
   U85225 : OAI221_X1 port map( B1 => n114477, B2 => n120038, C1 => n99278, C2 
                           => n120032, A => n117248, ZN => n117247);
   U85226 : OAI221_X1 port map( B1 => n114543, B2 => n119990, C1 => n114179, C2
                           => n119984, A => n117253, ZN => n117245);
   U85227 : NOR4_X1 port map( A1 => n117221, A2 => n117222, A3 => n117223, A4 
                           => n117224, ZN => n117220);
   U85228 : OAI221_X1 port map( B1 => n99211, B2 => n119966, C1 => n98875, C2 
                           => n119960, A => n117232, ZN => n117221);
   U85229 : OAI221_X1 port map( B1 => n114476, B2 => n120038, C1 => n99277, C2 
                           => n120032, A => n117225, ZN => n117224);
   U85230 : OAI221_X1 port map( B1 => n114542, B2 => n119990, C1 => n114178, C2
                           => n119984, A => n117230, ZN => n117222);
   U85231 : NOR4_X1 port map( A1 => n117198, A2 => n117199, A3 => n117200, A4 
                           => n117201, ZN => n117197);
   U85232 : OAI221_X1 port map( B1 => n99210, B2 => n119966, C1 => n98874, C2 
                           => n119960, A => n117209, ZN => n117198);
   U85233 : OAI221_X1 port map( B1 => n114475, B2 => n120038, C1 => n99276, C2 
                           => n120032, A => n117202, ZN => n117201);
   U85234 : OAI221_X1 port map( B1 => n114541, B2 => n119990, C1 => n114177, C2
                           => n119984, A => n117207, ZN => n117199);
   U85235 : NOR4_X1 port map( A1 => n117175, A2 => n117176, A3 => n117177, A4 
                           => n117178, ZN => n117174);
   U85236 : OAI221_X1 port map( B1 => n99209, B2 => n119966, C1 => n98873, C2 
                           => n119960, A => n117186, ZN => n117175);
   U85237 : OAI221_X1 port map( B1 => n114474, B2 => n120038, C1 => n99275, C2 
                           => n120032, A => n117179, ZN => n117178);
   U85238 : OAI221_X1 port map( B1 => n114540, B2 => n119990, C1 => n114176, C2
                           => n119984, A => n117184, ZN => n117176);
   U85239 : NOR4_X1 port map( A1 => n117152, A2 => n117153, A3 => n117154, A4 
                           => n117155, ZN => n117151);
   U85240 : OAI221_X1 port map( B1 => n99208, B2 => n119966, C1 => n98872, C2 
                           => n119960, A => n117163, ZN => n117152);
   U85241 : OAI221_X1 port map( B1 => n114473, B2 => n120038, C1 => n99274, C2 
                           => n120032, A => n117156, ZN => n117155);
   U85242 : OAI221_X1 port map( B1 => n114539, B2 => n119990, C1 => n114175, C2
                           => n119984, A => n117161, ZN => n117153);
   U85243 : NOR4_X1 port map( A1 => n117129, A2 => n117130, A3 => n117131, A4 
                           => n117132, ZN => n117128);
   U85244 : OAI221_X1 port map( B1 => n99207, B2 => n119967, C1 => n98871, C2 
                           => n119961, A => n117140, ZN => n117129);
   U85245 : OAI221_X1 port map( B1 => n114472, B2 => n120039, C1 => n99273, C2 
                           => n120033, A => n117133, ZN => n117132);
   U85246 : OAI221_X1 port map( B1 => n114538, B2 => n119991, C1 => n114174, C2
                           => n119985, A => n117138, ZN => n117130);
   U85247 : NOR4_X1 port map( A1 => n117106, A2 => n117107, A3 => n117108, A4 
                           => n117109, ZN => n117105);
   U85248 : OAI221_X1 port map( B1 => n99206, B2 => n119967, C1 => n98870, C2 
                           => n119961, A => n117117, ZN => n117106);
   U85249 : OAI221_X1 port map( B1 => n114471, B2 => n120039, C1 => n99272, C2 
                           => n120033, A => n117110, ZN => n117109);
   U85250 : OAI221_X1 port map( B1 => n114537, B2 => n119991, C1 => n114173, C2
                           => n119985, A => n117115, ZN => n117107);
   U85251 : NOR4_X1 port map( A1 => n117083, A2 => n117084, A3 => n117085, A4 
                           => n117086, ZN => n117082);
   U85252 : OAI221_X1 port map( B1 => n99205, B2 => n119967, C1 => n98869, C2 
                           => n119961, A => n117094, ZN => n117083);
   U85253 : OAI221_X1 port map( B1 => n114470, B2 => n120039, C1 => n99271, C2 
                           => n120033, A => n117087, ZN => n117086);
   U85254 : OAI221_X1 port map( B1 => n114536, B2 => n119991, C1 => n114172, C2
                           => n119985, A => n117092, ZN => n117084);
   U85255 : NOR4_X1 port map( A1 => n117060, A2 => n117061, A3 => n117062, A4 
                           => n117063, ZN => n117059);
   U85256 : OAI221_X1 port map( B1 => n99204, B2 => n119967, C1 => n98868, C2 
                           => n119961, A => n117071, ZN => n117060);
   U85257 : OAI221_X1 port map( B1 => n114469, B2 => n120039, C1 => n99270, C2 
                           => n120033, A => n117064, ZN => n117063);
   U85258 : OAI221_X1 port map( B1 => n114535, B2 => n119991, C1 => n114171, C2
                           => n119985, A => n117069, ZN => n117061);
   U85259 : NOR4_X1 port map( A1 => n117037, A2 => n117038, A3 => n117039, A4 
                           => n117040, ZN => n117036);
   U85260 : OAI221_X1 port map( B1 => n99203, B2 => n119967, C1 => n98867, C2 
                           => n119961, A => n117048, ZN => n117037);
   U85261 : OAI221_X1 port map( B1 => n114468, B2 => n120039, C1 => n99269, C2 
                           => n120033, A => n117041, ZN => n117040);
   U85262 : OAI221_X1 port map( B1 => n114534, B2 => n119991, C1 => n114170, C2
                           => n119985, A => n117046, ZN => n117038);
   U85263 : NOR4_X1 port map( A1 => n117014, A2 => n117015, A3 => n117016, A4 
                           => n117017, ZN => n117013);
   U85264 : OAI221_X1 port map( B1 => n99202, B2 => n119967, C1 => n98866, C2 
                           => n119961, A => n117025, ZN => n117014);
   U85265 : OAI221_X1 port map( B1 => n114467, B2 => n120039, C1 => n99268, C2 
                           => n120033, A => n117018, ZN => n117017);
   U85266 : OAI221_X1 port map( B1 => n114533, B2 => n119991, C1 => n114169, C2
                           => n119985, A => n117023, ZN => n117015);
   U85267 : NOR4_X1 port map( A1 => n116991, A2 => n116992, A3 => n116993, A4 
                           => n116994, ZN => n116990);
   U85268 : OAI221_X1 port map( B1 => n99201, B2 => n119967, C1 => n98865, C2 
                           => n119961, A => n117002, ZN => n116991);
   U85269 : OAI221_X1 port map( B1 => n114466, B2 => n120039, C1 => n99267, C2 
                           => n120033, A => n116995, ZN => n116994);
   U85270 : OAI221_X1 port map( B1 => n114532, B2 => n119991, C1 => n114168, C2
                           => n119985, A => n117000, ZN => n116992);
   U85271 : NOR4_X1 port map( A1 => n116968, A2 => n116969, A3 => n116970, A4 
                           => n116971, ZN => n116967);
   U85272 : OAI221_X1 port map( B1 => n99200, B2 => n119967, C1 => n98864, C2 
                           => n119961, A => n116979, ZN => n116968);
   U85273 : OAI221_X1 port map( B1 => n114465, B2 => n120039, C1 => n99266, C2 
                           => n120033, A => n116972, ZN => n116971);
   U85274 : OAI221_X1 port map( B1 => n114531, B2 => n119991, C1 => n114167, C2
                           => n119985, A => n116977, ZN => n116969);
   U85275 : NOR4_X1 port map( A1 => n116945, A2 => n116946, A3 => n116947, A4 
                           => n116948, ZN => n116944);
   U85276 : OAI221_X1 port map( B1 => n99199, B2 => n119967, C1 => n98863, C2 
                           => n119961, A => n116956, ZN => n116945);
   U85277 : OAI221_X1 port map( B1 => n114464, B2 => n120039, C1 => n99265, C2 
                           => n120033, A => n116949, ZN => n116948);
   U85278 : OAI221_X1 port map( B1 => n114530, B2 => n119991, C1 => n114166, C2
                           => n119985, A => n116954, ZN => n116946);
   U85279 : NOR4_X1 port map( A1 => n116922, A2 => n116923, A3 => n116924, A4 
                           => n116925, ZN => n116921);
   U85280 : OAI221_X1 port map( B1 => n99198, B2 => n119967, C1 => n98862, C2 
                           => n119961, A => n116933, ZN => n116922);
   U85281 : OAI221_X1 port map( B1 => n114463, B2 => n120039, C1 => n99264, C2 
                           => n120033, A => n116926, ZN => n116925);
   U85282 : OAI221_X1 port map( B1 => n114529, B2 => n119991, C1 => n114165, C2
                           => n119985, A => n116931, ZN => n116923);
   U85283 : NOR4_X1 port map( A1 => n116899, A2 => n116900, A3 => n116901, A4 
                           => n116902, ZN => n116898);
   U85284 : OAI221_X1 port map( B1 => n99197, B2 => n119967, C1 => n98861, C2 
                           => n119961, A => n116910, ZN => n116899);
   U85285 : OAI221_X1 port map( B1 => n114462, B2 => n120039, C1 => n99263, C2 
                           => n120033, A => n116903, ZN => n116902);
   U85286 : OAI221_X1 port map( B1 => n114528, B2 => n119991, C1 => n114164, C2
                           => n119985, A => n116908, ZN => n116900);
   U85287 : NOR4_X1 port map( A1 => n116876, A2 => n116877, A3 => n116878, A4 
                           => n116879, ZN => n116875);
   U85288 : OAI221_X1 port map( B1 => n99196, B2 => n119967, C1 => n98860, C2 
                           => n119961, A => n116887, ZN => n116876);
   U85289 : OAI221_X1 port map( B1 => n114461, B2 => n120039, C1 => n99262, C2 
                           => n120033, A => n116880, ZN => n116879);
   U85290 : OAI221_X1 port map( B1 => n114527, B2 => n119991, C1 => n114163, C2
                           => n119985, A => n116885, ZN => n116877);
   U85291 : NOR4_X1 port map( A1 => n116853, A2 => n116854, A3 => n116855, A4 
                           => n116856, ZN => n116852);
   U85292 : OAI221_X1 port map( B1 => n99195, B2 => n119968, C1 => n98859, C2 
                           => n119962, A => n116864, ZN => n116853);
   U85293 : OAI221_X1 port map( B1 => n114460, B2 => n120040, C1 => n99261, C2 
                           => n120034, A => n116857, ZN => n116856);
   U85294 : OAI221_X1 port map( B1 => n114526, B2 => n119992, C1 => n114162, C2
                           => n119986, A => n116862, ZN => n116854);
   U85295 : NOR4_X1 port map( A1 => n116830, A2 => n116831, A3 => n116832, A4 
                           => n116833, ZN => n116829);
   U85296 : OAI221_X1 port map( B1 => n99194, B2 => n119968, C1 => n98858, C2 
                           => n119962, A => n116841, ZN => n116830);
   U85297 : OAI221_X1 port map( B1 => n114459, B2 => n120040, C1 => n99260, C2 
                           => n120034, A => n116834, ZN => n116833);
   U85298 : OAI221_X1 port map( B1 => n114525, B2 => n119992, C1 => n114161, C2
                           => n119986, A => n116839, ZN => n116831);
   U85299 : NOR4_X1 port map( A1 => n116807, A2 => n116808, A3 => n116809, A4 
                           => n116810, ZN => n116806);
   U85300 : OAI221_X1 port map( B1 => n99193, B2 => n119968, C1 => n98857, C2 
                           => n119962, A => n116818, ZN => n116807);
   U85301 : OAI221_X1 port map( B1 => n114458, B2 => n120040, C1 => n99259, C2 
                           => n120034, A => n116811, ZN => n116810);
   U85302 : OAI221_X1 port map( B1 => n114524, B2 => n119992, C1 => n114160, C2
                           => n119986, A => n116816, ZN => n116808);
   U85303 : NOR4_X1 port map( A1 => n116784, A2 => n116785, A3 => n116786, A4 
                           => n116787, ZN => n116783);
   U85304 : OAI221_X1 port map( B1 => n99192, B2 => n119968, C1 => n98856, C2 
                           => n119962, A => n116795, ZN => n116784);
   U85305 : OAI221_X1 port map( B1 => n114457, B2 => n120040, C1 => n99258, C2 
                           => n120034, A => n116788, ZN => n116787);
   U85306 : OAI221_X1 port map( B1 => n114523, B2 => n119992, C1 => n114159, C2
                           => n119986, A => n116793, ZN => n116785);
   U85307 : NOR4_X1 port map( A1 => n116761, A2 => n116762, A3 => n116763, A4 
                           => n116764, ZN => n116760);
   U85308 : OAI221_X1 port map( B1 => n99191, B2 => n119968, C1 => n98855, C2 
                           => n119962, A => n116772, ZN => n116761);
   U85309 : OAI221_X1 port map( B1 => n114456, B2 => n120040, C1 => n99257, C2 
                           => n120034, A => n116765, ZN => n116764);
   U85310 : OAI221_X1 port map( B1 => n114522, B2 => n119992, C1 => n114158, C2
                           => n119986, A => n116770, ZN => n116762);
   U85311 : NOR4_X1 port map( A1 => n116738, A2 => n116739, A3 => n116740, A4 
                           => n116741, ZN => n116737);
   U85312 : OAI221_X1 port map( B1 => n99190, B2 => n119968, C1 => n98854, C2 
                           => n119962, A => n116749, ZN => n116738);
   U85313 : OAI221_X1 port map( B1 => n114455, B2 => n120040, C1 => n99256, C2 
                           => n120034, A => n116742, ZN => n116741);
   U85314 : OAI221_X1 port map( B1 => n114521, B2 => n119992, C1 => n114157, C2
                           => n119986, A => n116747, ZN => n116739);
   U85315 : NOR4_X1 port map( A1 => n116715, A2 => n116716, A3 => n116717, A4 
                           => n116718, ZN => n116714);
   U85316 : OAI221_X1 port map( B1 => n99189, B2 => n119968, C1 => n98853, C2 
                           => n119962, A => n116726, ZN => n116715);
   U85317 : OAI221_X1 port map( B1 => n114454, B2 => n120040, C1 => n99255, C2 
                           => n120034, A => n116719, ZN => n116718);
   U85318 : OAI221_X1 port map( B1 => n114520, B2 => n119992, C1 => n114156, C2
                           => n119986, A => n116724, ZN => n116716);
   U85319 : NOR4_X1 port map( A1 => n116692, A2 => n116693, A3 => n116694, A4 
                           => n116695, ZN => n116691);
   U85320 : OAI221_X1 port map( B1 => n99188, B2 => n119968, C1 => n98852, C2 
                           => n119962, A => n116703, ZN => n116692);
   U85321 : OAI221_X1 port map( B1 => n114453, B2 => n120040, C1 => n99254, C2 
                           => n120034, A => n116696, ZN => n116695);
   U85322 : OAI221_X1 port map( B1 => n114519, B2 => n119992, C1 => n114155, C2
                           => n119986, A => n116701, ZN => n116693);
   U85323 : NOR4_X1 port map( A1 => n116669, A2 => n116670, A3 => n116671, A4 
                           => n116672, ZN => n116668);
   U85324 : OAI221_X1 port map( B1 => n99187, B2 => n119968, C1 => n98851, C2 
                           => n119962, A => n116680, ZN => n116669);
   U85325 : OAI221_X1 port map( B1 => n114452, B2 => n120040, C1 => n99253, C2 
                           => n120034, A => n116673, ZN => n116672);
   U85326 : OAI221_X1 port map( B1 => n114518, B2 => n119992, C1 => n114154, C2
                           => n119986, A => n116678, ZN => n116670);
   U85327 : NOR4_X1 port map( A1 => n116646, A2 => n116647, A3 => n116648, A4 
                           => n116649, ZN => n116645);
   U85328 : OAI221_X1 port map( B1 => n99186, B2 => n119968, C1 => n98850, C2 
                           => n119962, A => n116657, ZN => n116646);
   U85329 : OAI221_X1 port map( B1 => n114451, B2 => n120040, C1 => n99252, C2 
                           => n120034, A => n116650, ZN => n116649);
   U85330 : OAI221_X1 port map( B1 => n114517, B2 => n119992, C1 => n114153, C2
                           => n119986, A => n116655, ZN => n116647);
   U85331 : NOR4_X1 port map( A1 => n116623, A2 => n116624, A3 => n116625, A4 
                           => n116626, ZN => n116622);
   U85332 : OAI221_X1 port map( B1 => n99185, B2 => n119968, C1 => n98849, C2 
                           => n119962, A => n116634, ZN => n116623);
   U85333 : OAI221_X1 port map( B1 => n114450, B2 => n120040, C1 => n99251, C2 
                           => n120034, A => n116627, ZN => n116626);
   U85334 : OAI221_X1 port map( B1 => n114516, B2 => n119992, C1 => n114152, C2
                           => n119986, A => n116632, ZN => n116624);
   U85335 : NOR4_X1 port map( A1 => n116600, A2 => n116601, A3 => n116602, A4 
                           => n116603, ZN => n116599);
   U85336 : OAI221_X1 port map( B1 => n99184, B2 => n119968, C1 => n98848, C2 
                           => n119962, A => n116611, ZN => n116600);
   U85337 : OAI221_X1 port map( B1 => n114449, B2 => n120040, C1 => n99250, C2 
                           => n120034, A => n116604, ZN => n116603);
   U85338 : OAI221_X1 port map( B1 => n114515, B2 => n119992, C1 => n114151, C2
                           => n119986, A => n116609, ZN => n116601);
   U85339 : NOR4_X1 port map( A1 => n115151, A2 => n115152, A3 => n115153, A4 
                           => n115154, ZN => n115150);
   U85340 : OAI221_X1 port map( B1 => n114528, B2 => n120165, C1 => n114462, C2
                           => n120159, A => n115162, ZN => n115151);
   U85341 : OAI221_X1 port map( B1 => n98999, B2 => n120189, C1 => n114396, C2 
                           => n120183, A => n115160, ZN => n115152);
   U85342 : OAI221_X1 port map( B1 => n99598, B2 => n120237, C1 => n114005, C2 
                           => n120231, A => n115155, ZN => n115154);
   U85343 : NOR4_X1 port map( A1 => n115123, A2 => n115124, A3 => n115125, A4 
                           => n115126, ZN => n115122);
   U85344 : OAI221_X1 port map( B1 => n114527, B2 => n120165, C1 => n114461, C2
                           => n120159, A => n115134, ZN => n115123);
   U85345 : OAI221_X1 port map( B1 => n98998, B2 => n120189, C1 => n114395, C2 
                           => n120183, A => n115132, ZN => n115124);
   U85346 : OAI221_X1 port map( B1 => n99597, B2 => n120237, C1 => n114004, C2 
                           => n120231, A => n115127, ZN => n115126);
   U85347 : NOR4_X1 port map( A1 => n115095, A2 => n115096, A3 => n115097, A4 
                           => n115098, ZN => n115094);
   U85348 : OAI221_X1 port map( B1 => n114526, B2 => n120166, C1 => n114460, C2
                           => n120160, A => n115106, ZN => n115095);
   U85349 : OAI221_X1 port map( B1 => n98997, B2 => n120190, C1 => n114394, C2 
                           => n120184, A => n115104, ZN => n115096);
   U85350 : OAI221_X1 port map( B1 => n99596, B2 => n120238, C1 => n114003, C2 
                           => n120232, A => n115099, ZN => n115098);
   U85351 : NOR4_X1 port map( A1 => n115067, A2 => n115068, A3 => n115069, A4 
                           => n115070, ZN => n115066);
   U85352 : OAI221_X1 port map( B1 => n114525, B2 => n120166, C1 => n114459, C2
                           => n120160, A => n115078, ZN => n115067);
   U85353 : OAI221_X1 port map( B1 => n98996, B2 => n120190, C1 => n114393, C2 
                           => n120184, A => n115076, ZN => n115068);
   U85354 : OAI221_X1 port map( B1 => n99595, B2 => n120238, C1 => n114002, C2 
                           => n120232, A => n115071, ZN => n115070);
   U85355 : NOR4_X1 port map( A1 => n115039, A2 => n115040, A3 => n115041, A4 
                           => n115042, ZN => n115038);
   U85356 : OAI221_X1 port map( B1 => n114524, B2 => n120166, C1 => n114458, C2
                           => n120160, A => n115050, ZN => n115039);
   U85357 : OAI221_X1 port map( B1 => n98995, B2 => n120190, C1 => n114392, C2 
                           => n120184, A => n115048, ZN => n115040);
   U85358 : OAI221_X1 port map( B1 => n99594, B2 => n120238, C1 => n114001, C2 
                           => n120232, A => n115043, ZN => n115042);
   U85359 : NOR4_X1 port map( A1 => n115011, A2 => n115012, A3 => n115013, A4 
                           => n115014, ZN => n115010);
   U85360 : OAI221_X1 port map( B1 => n114523, B2 => n120166, C1 => n114457, C2
                           => n120160, A => n115022, ZN => n115011);
   U85361 : OAI221_X1 port map( B1 => n98994, B2 => n120190, C1 => n114391, C2 
                           => n120184, A => n115020, ZN => n115012);
   U85362 : OAI221_X1 port map( B1 => n99593, B2 => n120238, C1 => n114000, C2 
                           => n120232, A => n115015, ZN => n115014);
   U85363 : NOR4_X1 port map( A1 => n114983, A2 => n114984, A3 => n114985, A4 
                           => n114986, ZN => n114982);
   U85364 : OAI221_X1 port map( B1 => n114522, B2 => n120166, C1 => n114456, C2
                           => n120160, A => n114994, ZN => n114983);
   U85365 : OAI221_X1 port map( B1 => n98993, B2 => n120190, C1 => n114390, C2 
                           => n120184, A => n114992, ZN => n114984);
   U85366 : OAI221_X1 port map( B1 => n99592, B2 => n120238, C1 => n113999, C2 
                           => n120232, A => n114987, ZN => n114986);
   U85367 : NOR4_X1 port map( A1 => n114955, A2 => n114956, A3 => n114957, A4 
                           => n114958, ZN => n114954);
   U85368 : OAI221_X1 port map( B1 => n114521, B2 => n120166, C1 => n114455, C2
                           => n120160, A => n114966, ZN => n114955);
   U85369 : OAI221_X1 port map( B1 => n98992, B2 => n120190, C1 => n114389, C2 
                           => n120184, A => n114964, ZN => n114956);
   U85370 : OAI221_X1 port map( B1 => n99591, B2 => n120238, C1 => n113998, C2 
                           => n120232, A => n114959, ZN => n114958);
   U85371 : NOR4_X1 port map( A1 => n114927, A2 => n114928, A3 => n114929, A4 
                           => n114930, ZN => n114926);
   U85372 : OAI221_X1 port map( B1 => n114520, B2 => n120166, C1 => n114454, C2
                           => n120160, A => n114938, ZN => n114927);
   U85373 : OAI221_X1 port map( B1 => n98991, B2 => n120190, C1 => n114388, C2 
                           => n120184, A => n114936, ZN => n114928);
   U85374 : OAI221_X1 port map( B1 => n99590, B2 => n120238, C1 => n113997, C2 
                           => n120232, A => n114931, ZN => n114930);
   U85375 : NOR4_X1 port map( A1 => n114899, A2 => n114900, A3 => n114901, A4 
                           => n114902, ZN => n114898);
   U85376 : OAI221_X1 port map( B1 => n114519, B2 => n120166, C1 => n114453, C2
                           => n120160, A => n114910, ZN => n114899);
   U85377 : OAI221_X1 port map( B1 => n98990, B2 => n120190, C1 => n114387, C2 
                           => n120184, A => n114908, ZN => n114900);
   U85378 : OAI221_X1 port map( B1 => n99589, B2 => n120238, C1 => n113996, C2 
                           => n120232, A => n114903, ZN => n114902);
   U85379 : NOR4_X1 port map( A1 => n114871, A2 => n114872, A3 => n114873, A4 
                           => n114874, ZN => n114870);
   U85380 : OAI221_X1 port map( B1 => n114518, B2 => n120166, C1 => n114452, C2
                           => n120160, A => n114882, ZN => n114871);
   U85381 : OAI221_X1 port map( B1 => n98989, B2 => n120190, C1 => n114386, C2 
                           => n120184, A => n114880, ZN => n114872);
   U85382 : OAI221_X1 port map( B1 => n99588, B2 => n120238, C1 => n113995, C2 
                           => n120232, A => n114875, ZN => n114874);
   U85383 : NOR4_X1 port map( A1 => n114843, A2 => n114844, A3 => n114845, A4 
                           => n114846, ZN => n114842);
   U85384 : OAI221_X1 port map( B1 => n114517, B2 => n120166, C1 => n114451, C2
                           => n120160, A => n114854, ZN => n114843);
   U85385 : OAI221_X1 port map( B1 => n98988, B2 => n120190, C1 => n114385, C2 
                           => n120184, A => n114852, ZN => n114844);
   U85386 : OAI221_X1 port map( B1 => n99587, B2 => n120238, C1 => n113994, C2 
                           => n120232, A => n114847, ZN => n114846);
   U85387 : NOR4_X1 port map( A1 => n114815, A2 => n114816, A3 => n114817, A4 
                           => n114818, ZN => n114814);
   U85388 : OAI221_X1 port map( B1 => n114516, B2 => n120166, C1 => n114450, C2
                           => n120160, A => n114826, ZN => n114815);
   U85389 : OAI221_X1 port map( B1 => n98987, B2 => n120190, C1 => n114384, C2 
                           => n120184, A => n114824, ZN => n114816);
   U85390 : OAI221_X1 port map( B1 => n99586, B2 => n120238, C1 => n113993, C2 
                           => n120232, A => n114819, ZN => n114818);
   U85391 : NOR4_X1 port map( A1 => n114787, A2 => n114788, A3 => n114789, A4 
                           => n114790, ZN => n114786);
   U85392 : OAI221_X1 port map( B1 => n114515, B2 => n120166, C1 => n114449, C2
                           => n120160, A => n114798, ZN => n114787);
   U85393 : OAI221_X1 port map( B1 => n98986, B2 => n120190, C1 => n114383, C2 
                           => n120184, A => n114796, ZN => n114788);
   U85394 : OAI221_X1 port map( B1 => n99585, B2 => n120238, C1 => n113992, C2 
                           => n120232, A => n114791, ZN => n114790);
   U85395 : NOR4_X1 port map( A1 => n116439, A2 => n116440, A3 => n116441, A4 
                           => n116442, ZN => n116438);
   U85396 : OAI221_X1 port map( B1 => n114574, B2 => n120162, C1 => n114508, C2
                           => n120156, A => n116460, ZN => n116439);
   U85397 : OAI221_X1 port map( B1 => n99045, B2 => n120186, C1 => n114442, C2 
                           => n120180, A => n116455, ZN => n116440);
   U85398 : OAI221_X1 port map( B1 => n99644, B2 => n120234, C1 => n114051, C2 
                           => n120228, A => n116443, ZN => n116442);
   U85399 : NOR4_X1 port map( A1 => n116411, A2 => n116412, A3 => n116413, A4 
                           => n116414, ZN => n116410);
   U85400 : OAI221_X1 port map( B1 => n114573, B2 => n120162, C1 => n114507, C2
                           => n120156, A => n116422, ZN => n116411);
   U85401 : OAI221_X1 port map( B1 => n99044, B2 => n120186, C1 => n114441, C2 
                           => n120180, A => n116420, ZN => n116412);
   U85402 : OAI221_X1 port map( B1 => n99643, B2 => n120234, C1 => n114050, C2 
                           => n120228, A => n116415, ZN => n116414);
   U85403 : NOR4_X1 port map( A1 => n116383, A2 => n116384, A3 => n116385, A4 
                           => n116386, ZN => n116382);
   U85404 : OAI221_X1 port map( B1 => n114572, B2 => n120162, C1 => n114506, C2
                           => n120156, A => n116394, ZN => n116383);
   U85405 : OAI221_X1 port map( B1 => n99043, B2 => n120186, C1 => n114440, C2 
                           => n120180, A => n116392, ZN => n116384);
   U85406 : OAI221_X1 port map( B1 => n99642, B2 => n120234, C1 => n114049, C2 
                           => n120228, A => n116387, ZN => n116386);
   U85407 : NOR4_X1 port map( A1 => n116355, A2 => n116356, A3 => n116357, A4 
                           => n116358, ZN => n116354);
   U85408 : OAI221_X1 port map( B1 => n114571, B2 => n120162, C1 => n114505, C2
                           => n120156, A => n116366, ZN => n116355);
   U85409 : OAI221_X1 port map( B1 => n99042, B2 => n120186, C1 => n114439, C2 
                           => n120180, A => n116364, ZN => n116356);
   U85410 : OAI221_X1 port map( B1 => n99641, B2 => n120234, C1 => n114048, C2 
                           => n120228, A => n116359, ZN => n116358);
   U85411 : NOR4_X1 port map( A1 => n117785, A2 => n117786, A3 => n117787, A4 
                           => n117788, ZN => n117784);
   U85412 : OAI221_X1 port map( B1 => n99236, B2 => n119964, C1 => n98900, C2 
                           => n119958, A => n117796, ZN => n117785);
   U85413 : OAI221_X1 port map( B1 => n114501, B2 => n120036, C1 => n99302, C2 
                           => n120030, A => n117789, ZN => n117788);
   U85414 : OAI221_X1 port map( B1 => n114567, B2 => n119988, C1 => n114203, C2
                           => n119982, A => n117794, ZN => n117786);
   U85415 : NOR4_X1 port map( A1 => n117763, A2 => n117764, A3 => n117765, A4 
                           => n117766, ZN => n117762);
   U85416 : OAI221_X1 port map( B1 => n99235, B2 => n119964, C1 => n98899, C2 
                           => n119958, A => n117774, ZN => n117763);
   U85417 : OAI221_X1 port map( B1 => n114500, B2 => n120036, C1 => n99301, C2 
                           => n120030, A => n117767, ZN => n117766);
   U85418 : OAI221_X1 port map( B1 => n114566, B2 => n119988, C1 => n114202, C2
                           => n119982, A => n117772, ZN => n117764);
   U85419 : NOR4_X1 port map( A1 => n117741, A2 => n117742, A3 => n117743, A4 
                           => n117744, ZN => n117740);
   U85420 : OAI221_X1 port map( B1 => n99234, B2 => n119964, C1 => n98898, C2 
                           => n119958, A => n117752, ZN => n117741);
   U85421 : OAI221_X1 port map( B1 => n114499, B2 => n120036, C1 => n99300, C2 
                           => n120030, A => n117745, ZN => n117744);
   U85422 : OAI221_X1 port map( B1 => n114565, B2 => n119988, C1 => n114201, C2
                           => n119982, A => n117750, ZN => n117742);
   U85423 : NOR4_X1 port map( A1 => n117719, A2 => n117720, A3 => n117721, A4 
                           => n117722, ZN => n117718);
   U85424 : OAI221_X1 port map( B1 => n99233, B2 => n119964, C1 => n98897, C2 
                           => n119958, A => n117730, ZN => n117719);
   U85425 : OAI221_X1 port map( B1 => n114498, B2 => n120036, C1 => n99299, C2 
                           => n120030, A => n117723, ZN => n117722);
   U85426 : OAI221_X1 port map( B1 => n114564, B2 => n119988, C1 => n114200, C2
                           => n119982, A => n117728, ZN => n117720);
   U85427 : NOR4_X1 port map( A1 => n117939, A2 => n117940, A3 => n117941, A4 
                           => n117942, ZN => n117938);
   U85428 : OAI221_X1 port map( B1 => n99243, B2 => n119964, C1 => n98907, C2 
                           => n119958, A => n117960, ZN => n117939);
   U85429 : OAI221_X1 port map( B1 => n114508, B2 => n120036, C1 => n99309, C2 
                           => n120030, A => n117943, ZN => n117942);
   U85430 : OAI221_X1 port map( B1 => n114574, B2 => n119988, C1 => n114210, C2
                           => n119982, A => n117956, ZN => n117940);
   U85431 : NOR4_X1 port map( A1 => n117917, A2 => n117918, A3 => n117919, A4 
                           => n117920, ZN => n117916);
   U85432 : OAI221_X1 port map( B1 => n99242, B2 => n119964, C1 => n98906, C2 
                           => n119958, A => n117928, ZN => n117917);
   U85433 : OAI221_X1 port map( B1 => n114507, B2 => n120036, C1 => n99308, C2 
                           => n120030, A => n117921, ZN => n117920);
   U85434 : OAI221_X1 port map( B1 => n114573, B2 => n119988, C1 => n114209, C2
                           => n119982, A => n117926, ZN => n117918);
   U85435 : NOR4_X1 port map( A1 => n117895, A2 => n117896, A3 => n117897, A4 
                           => n117898, ZN => n117894);
   U85436 : OAI221_X1 port map( B1 => n99241, B2 => n119964, C1 => n98905, C2 
                           => n119958, A => n117906, ZN => n117895);
   U85437 : OAI221_X1 port map( B1 => n114506, B2 => n120036, C1 => n99307, C2 
                           => n120030, A => n117899, ZN => n117898);
   U85438 : OAI221_X1 port map( B1 => n114572, B2 => n119988, C1 => n114208, C2
                           => n119982, A => n117904, ZN => n117896);
   U85439 : NOR4_X1 port map( A1 => n117873, A2 => n117874, A3 => n117875, A4 
                           => n117876, ZN => n117872);
   U85440 : OAI221_X1 port map( B1 => n99240, B2 => n119964, C1 => n98904, C2 
                           => n119958, A => n117884, ZN => n117873);
   U85441 : OAI221_X1 port map( B1 => n114505, B2 => n120036, C1 => n99306, C2 
                           => n120030, A => n117877, ZN => n117876);
   U85442 : OAI221_X1 port map( B1 => n114571, B2 => n119988, C1 => n114207, C2
                           => n119982, A => n117882, ZN => n117874);
   U85443 : NOR4_X1 port map( A1 => n117851, A2 => n117852, A3 => n117853, A4 
                           => n117854, ZN => n117850);
   U85444 : OAI221_X1 port map( B1 => n99239, B2 => n119964, C1 => n98903, C2 
                           => n119958, A => n117862, ZN => n117851);
   U85445 : OAI221_X1 port map( B1 => n114504, B2 => n120036, C1 => n99305, C2 
                           => n120030, A => n117855, ZN => n117854);
   U85446 : OAI221_X1 port map( B1 => n114570, B2 => n119988, C1 => n114206, C2
                           => n119982, A => n117860, ZN => n117852);
   U85447 : NOR4_X1 port map( A1 => n117829, A2 => n117830, A3 => n117831, A4 
                           => n117832, ZN => n117828);
   U85448 : OAI221_X1 port map( B1 => n99238, B2 => n119964, C1 => n98902, C2 
                           => n119958, A => n117840, ZN => n117829);
   U85449 : OAI221_X1 port map( B1 => n114503, B2 => n120036, C1 => n99304, C2 
                           => n120030, A => n117833, ZN => n117832);
   U85450 : OAI221_X1 port map( B1 => n114569, B2 => n119988, C1 => n114205, C2
                           => n119982, A => n117838, ZN => n117830);
   U85451 : NOR4_X1 port map( A1 => n117807, A2 => n117808, A3 => n117809, A4 
                           => n117810, ZN => n117806);
   U85452 : OAI221_X1 port map( B1 => n99237, B2 => n119964, C1 => n98901, C2 
                           => n119958, A => n117818, ZN => n117807);
   U85453 : OAI221_X1 port map( B1 => n114502, B2 => n120036, C1 => n99303, C2 
                           => n120030, A => n117811, ZN => n117810);
   U85454 : OAI221_X1 port map( B1 => n114568, B2 => n119988, C1 => n114204, C2
                           => n119982, A => n117816, ZN => n117808);
   U85455 : NOR4_X1 port map( A1 => n116327, A2 => n116328, A3 => n116329, A4 
                           => n116330, ZN => n116326);
   U85456 : OAI221_X1 port map( B1 => n114570, B2 => n120162, C1 => n114504, C2
                           => n120156, A => n116338, ZN => n116327);
   U85457 : OAI221_X1 port map( B1 => n99041, B2 => n120186, C1 => n114438, C2 
                           => n120180, A => n116336, ZN => n116328);
   U85458 : OAI221_X1 port map( B1 => n99640, B2 => n120234, C1 => n114047, C2 
                           => n120228, A => n116331, ZN => n116330);
   U85459 : NOR4_X1 port map( A1 => n116299, A2 => n116300, A3 => n116301, A4 
                           => n116302, ZN => n116298);
   U85460 : OAI221_X1 port map( B1 => n114569, B2 => n120162, C1 => n114503, C2
                           => n120156, A => n116310, ZN => n116299);
   U85461 : OAI221_X1 port map( B1 => n99040, B2 => n120186, C1 => n114437, C2 
                           => n120180, A => n116308, ZN => n116300);
   U85462 : OAI221_X1 port map( B1 => n99639, B2 => n120234, C1 => n114046, C2 
                           => n120228, A => n116303, ZN => n116302);
   U85463 : NOR4_X1 port map( A1 => n116271, A2 => n116272, A3 => n116273, A4 
                           => n116274, ZN => n116270);
   U85464 : OAI221_X1 port map( B1 => n114568, B2 => n120162, C1 => n114502, C2
                           => n120156, A => n116282, ZN => n116271);
   U85465 : OAI221_X1 port map( B1 => n99039, B2 => n120186, C1 => n114436, C2 
                           => n120180, A => n116280, ZN => n116272);
   U85466 : OAI221_X1 port map( B1 => n99638, B2 => n120234, C1 => n114045, C2 
                           => n120228, A => n116275, ZN => n116274);
   U85467 : NOR4_X1 port map( A1 => n116243, A2 => n116244, A3 => n116245, A4 
                           => n116246, ZN => n116242);
   U85468 : OAI221_X1 port map( B1 => n114567, B2 => n120162, C1 => n114501, C2
                           => n120156, A => n116254, ZN => n116243);
   U85469 : OAI221_X1 port map( B1 => n99038, B2 => n120186, C1 => n114435, C2 
                           => n120180, A => n116252, ZN => n116244);
   U85470 : OAI221_X1 port map( B1 => n99637, B2 => n120234, C1 => n114044, C2 
                           => n120228, A => n116247, ZN => n116246);
   U85471 : NOR4_X1 port map( A1 => n116215, A2 => n116216, A3 => n116217, A4 
                           => n116218, ZN => n116214);
   U85472 : OAI221_X1 port map( B1 => n114566, B2 => n120162, C1 => n114500, C2
                           => n120156, A => n116226, ZN => n116215);
   U85473 : OAI221_X1 port map( B1 => n99037, B2 => n120186, C1 => n114434, C2 
                           => n120180, A => n116224, ZN => n116216);
   U85474 : OAI221_X1 port map( B1 => n99636, B2 => n120234, C1 => n114043, C2 
                           => n120228, A => n116219, ZN => n116218);
   U85475 : NOR4_X1 port map( A1 => n116187, A2 => n116188, A3 => n116189, A4 
                           => n116190, ZN => n116186);
   U85476 : OAI221_X1 port map( B1 => n114565, B2 => n120162, C1 => n114499, C2
                           => n120156, A => n116198, ZN => n116187);
   U85477 : OAI221_X1 port map( B1 => n99036, B2 => n120186, C1 => n114433, C2 
                           => n120180, A => n116196, ZN => n116188);
   U85478 : OAI221_X1 port map( B1 => n99635, B2 => n120234, C1 => n114042, C2 
                           => n120228, A => n116191, ZN => n116190);
   U85479 : NOR4_X1 port map( A1 => n116159, A2 => n116160, A3 => n116161, A4 
                           => n116162, ZN => n116158);
   U85480 : OAI221_X1 port map( B1 => n114564, B2 => n120162, C1 => n114498, C2
                           => n120156, A => n116170, ZN => n116159);
   U85481 : OAI221_X1 port map( B1 => n99035, B2 => n120186, C1 => n114432, C2 
                           => n120180, A => n116168, ZN => n116160);
   U85482 : OAI221_X1 port map( B1 => n99634, B2 => n120234, C1 => n114041, C2 
                           => n120228, A => n116163, ZN => n116162);
   U85483 : NOR4_X1 port map( A1 => n116131, A2 => n116132, A3 => n116133, A4 
                           => n116134, ZN => n116130);
   U85484 : OAI221_X1 port map( B1 => n114563, B2 => n120162, C1 => n114497, C2
                           => n120156, A => n116142, ZN => n116131);
   U85485 : OAI221_X1 port map( B1 => n99034, B2 => n120186, C1 => n114431, C2 
                           => n120180, A => n116140, ZN => n116132);
   U85486 : OAI221_X1 port map( B1 => n99633, B2 => n120234, C1 => n114040, C2 
                           => n120228, A => n116135, ZN => n116134);
   U85487 : NOR4_X1 port map( A1 => n116103, A2 => n116104, A3 => n116105, A4 
                           => n116106, ZN => n116102);
   U85488 : OAI221_X1 port map( B1 => n114562, B2 => n120163, C1 => n114496, C2
                           => n120157, A => n116114, ZN => n116103);
   U85489 : OAI221_X1 port map( B1 => n99033, B2 => n120187, C1 => n114430, C2 
                           => n120181, A => n116112, ZN => n116104);
   U85490 : OAI221_X1 port map( B1 => n99632, B2 => n120235, C1 => n114039, C2 
                           => n120229, A => n116107, ZN => n116106);
   U85491 : NOR4_X1 port map( A1 => n116075, A2 => n116076, A3 => n116077, A4 
                           => n116078, ZN => n116074);
   U85492 : OAI221_X1 port map( B1 => n114561, B2 => n120163, C1 => n114495, C2
                           => n120157, A => n116086, ZN => n116075);
   U85493 : OAI221_X1 port map( B1 => n99032, B2 => n120187, C1 => n114429, C2 
                           => n120181, A => n116084, ZN => n116076);
   U85494 : OAI221_X1 port map( B1 => n99631, B2 => n120235, C1 => n114038, C2 
                           => n120229, A => n116079, ZN => n116078);
   U85495 : NOR4_X1 port map( A1 => n116047, A2 => n116048, A3 => n116049, A4 
                           => n116050, ZN => n116046);
   U85496 : OAI221_X1 port map( B1 => n114560, B2 => n120163, C1 => n114494, C2
                           => n120157, A => n116058, ZN => n116047);
   U85497 : OAI221_X1 port map( B1 => n99031, B2 => n120187, C1 => n114428, C2 
                           => n120181, A => n116056, ZN => n116048);
   U85498 : OAI221_X1 port map( B1 => n99630, B2 => n120235, C1 => n114037, C2 
                           => n120229, A => n116051, ZN => n116050);
   U85499 : NOR4_X1 port map( A1 => n116019, A2 => n116020, A3 => n116021, A4 
                           => n116022, ZN => n116018);
   U85500 : OAI221_X1 port map( B1 => n114559, B2 => n120163, C1 => n114493, C2
                           => n120157, A => n116030, ZN => n116019);
   U85501 : OAI221_X1 port map( B1 => n99030, B2 => n120187, C1 => n114427, C2 
                           => n120181, A => n116028, ZN => n116020);
   U85502 : OAI221_X1 port map( B1 => n99629, B2 => n120235, C1 => n114036, C2 
                           => n120229, A => n116023, ZN => n116022);
   U85503 : NOR4_X1 port map( A1 => n115991, A2 => n115992, A3 => n115993, A4 
                           => n115994, ZN => n115990);
   U85504 : OAI221_X1 port map( B1 => n114558, B2 => n120163, C1 => n114492, C2
                           => n120157, A => n116002, ZN => n115991);
   U85505 : OAI221_X1 port map( B1 => n99029, B2 => n120187, C1 => n114426, C2 
                           => n120181, A => n116000, ZN => n115992);
   U85506 : OAI221_X1 port map( B1 => n99628, B2 => n120235, C1 => n114035, C2 
                           => n120229, A => n115995, ZN => n115994);
   U85507 : NOR4_X1 port map( A1 => n115963, A2 => n115964, A3 => n115965, A4 
                           => n115966, ZN => n115962);
   U85508 : OAI221_X1 port map( B1 => n114557, B2 => n120163, C1 => n114491, C2
                           => n120157, A => n115974, ZN => n115963);
   U85509 : OAI221_X1 port map( B1 => n99028, B2 => n120187, C1 => n114425, C2 
                           => n120181, A => n115972, ZN => n115964);
   U85510 : OAI221_X1 port map( B1 => n99627, B2 => n120235, C1 => n114034, C2 
                           => n120229, A => n115967, ZN => n115966);
   U85511 : NOR4_X1 port map( A1 => n115935, A2 => n115936, A3 => n115937, A4 
                           => n115938, ZN => n115934);
   U85512 : OAI221_X1 port map( B1 => n114556, B2 => n120163, C1 => n114490, C2
                           => n120157, A => n115946, ZN => n115935);
   U85513 : OAI221_X1 port map( B1 => n99027, B2 => n120187, C1 => n114424, C2 
                           => n120181, A => n115944, ZN => n115936);
   U85514 : OAI221_X1 port map( B1 => n99626, B2 => n120235, C1 => n114033, C2 
                           => n120229, A => n115939, ZN => n115938);
   U85515 : NOR4_X1 port map( A1 => n115907, A2 => n115908, A3 => n115909, A4 
                           => n115910, ZN => n115906);
   U85516 : OAI221_X1 port map( B1 => n114555, B2 => n120163, C1 => n114489, C2
                           => n120157, A => n115918, ZN => n115907);
   U85517 : OAI221_X1 port map( B1 => n99026, B2 => n120187, C1 => n114423, C2 
                           => n120181, A => n115916, ZN => n115908);
   U85518 : OAI221_X1 port map( B1 => n99625, B2 => n120235, C1 => n114032, C2 
                           => n120229, A => n115911, ZN => n115910);
   U85519 : NOR4_X1 port map( A1 => n115879, A2 => n115880, A3 => n115881, A4 
                           => n115882, ZN => n115878);
   U85520 : OAI221_X1 port map( B1 => n114554, B2 => n120163, C1 => n114488, C2
                           => n120157, A => n115890, ZN => n115879);
   U85521 : OAI221_X1 port map( B1 => n99025, B2 => n120187, C1 => n114422, C2 
                           => n120181, A => n115888, ZN => n115880);
   U85522 : OAI221_X1 port map( B1 => n99624, B2 => n120235, C1 => n114031, C2 
                           => n120229, A => n115883, ZN => n115882);
   U85523 : NOR4_X1 port map( A1 => n115851, A2 => n115852, A3 => n115853, A4 
                           => n115854, ZN => n115850);
   U85524 : OAI221_X1 port map( B1 => n114553, B2 => n120163, C1 => n114487, C2
                           => n120157, A => n115862, ZN => n115851);
   U85525 : OAI221_X1 port map( B1 => n99024, B2 => n120187, C1 => n114421, C2 
                           => n120181, A => n115860, ZN => n115852);
   U85526 : OAI221_X1 port map( B1 => n99623, B2 => n120235, C1 => n114030, C2 
                           => n120229, A => n115855, ZN => n115854);
   U85527 : NOR4_X1 port map( A1 => n115823, A2 => n115824, A3 => n115825, A4 
                           => n115826, ZN => n115822);
   U85528 : OAI221_X1 port map( B1 => n114552, B2 => n120163, C1 => n114486, C2
                           => n120157, A => n115834, ZN => n115823);
   U85529 : OAI221_X1 port map( B1 => n99023, B2 => n120187, C1 => n114420, C2 
                           => n120181, A => n115832, ZN => n115824);
   U85530 : OAI221_X1 port map( B1 => n99622, B2 => n120235, C1 => n114029, C2 
                           => n120229, A => n115827, ZN => n115826);
   U85531 : NOR4_X1 port map( A1 => n115795, A2 => n115796, A3 => n115797, A4 
                           => n115798, ZN => n115794);
   U85532 : OAI221_X1 port map( B1 => n114551, B2 => n120163, C1 => n114485, C2
                           => n120157, A => n115806, ZN => n115795);
   U85533 : OAI221_X1 port map( B1 => n99022, B2 => n120187, C1 => n114419, C2 
                           => n120181, A => n115804, ZN => n115796);
   U85534 : OAI221_X1 port map( B1 => n99621, B2 => n120235, C1 => n114028, C2 
                           => n120229, A => n115799, ZN => n115798);
   U85535 : NOR4_X1 port map( A1 => n115767, A2 => n115768, A3 => n115769, A4 
                           => n115770, ZN => n115766);
   U85536 : OAI221_X1 port map( B1 => n114550, B2 => n120164, C1 => n114484, C2
                           => n120158, A => n115778, ZN => n115767);
   U85537 : OAI221_X1 port map( B1 => n99021, B2 => n120188, C1 => n114418, C2 
                           => n120182, A => n115776, ZN => n115768);
   U85538 : OAI221_X1 port map( B1 => n99620, B2 => n120236, C1 => n114027, C2 
                           => n120230, A => n115771, ZN => n115770);
   U85539 : NOR4_X1 port map( A1 => n115739, A2 => n115740, A3 => n115741, A4 
                           => n115742, ZN => n115738);
   U85540 : OAI221_X1 port map( B1 => n114549, B2 => n120164, C1 => n114483, C2
                           => n120158, A => n115750, ZN => n115739);
   U85541 : OAI221_X1 port map( B1 => n99020, B2 => n120188, C1 => n114417, C2 
                           => n120182, A => n115748, ZN => n115740);
   U85542 : OAI221_X1 port map( B1 => n99619, B2 => n120236, C1 => n114026, C2 
                           => n120230, A => n115743, ZN => n115742);
   U85543 : NOR4_X1 port map( A1 => n115711, A2 => n115712, A3 => n115713, A4 
                           => n115714, ZN => n115710);
   U85544 : OAI221_X1 port map( B1 => n114548, B2 => n120164, C1 => n114482, C2
                           => n120158, A => n115722, ZN => n115711);
   U85545 : OAI221_X1 port map( B1 => n99019, B2 => n120188, C1 => n114416, C2 
                           => n120182, A => n115720, ZN => n115712);
   U85546 : OAI221_X1 port map( B1 => n99618, B2 => n120236, C1 => n114025, C2 
                           => n120230, A => n115715, ZN => n115714);
   U85547 : NOR4_X1 port map( A1 => n115683, A2 => n115684, A3 => n115685, A4 
                           => n115686, ZN => n115682);
   U85548 : OAI221_X1 port map( B1 => n114547, B2 => n120164, C1 => n114481, C2
                           => n120158, A => n115694, ZN => n115683);
   U85549 : OAI221_X1 port map( B1 => n99018, B2 => n120188, C1 => n114415, C2 
                           => n120182, A => n115692, ZN => n115684);
   U85550 : OAI221_X1 port map( B1 => n99617, B2 => n120236, C1 => n114024, C2 
                           => n120230, A => n115687, ZN => n115686);
   U85551 : NOR4_X1 port map( A1 => n115655, A2 => n115656, A3 => n115657, A4 
                           => n115658, ZN => n115654);
   U85552 : OAI221_X1 port map( B1 => n114546, B2 => n120164, C1 => n114480, C2
                           => n120158, A => n115666, ZN => n115655);
   U85553 : OAI221_X1 port map( B1 => n99017, B2 => n120188, C1 => n114414, C2 
                           => n120182, A => n115664, ZN => n115656);
   U85554 : OAI221_X1 port map( B1 => n99616, B2 => n120236, C1 => n114023, C2 
                           => n120230, A => n115659, ZN => n115658);
   U85555 : NOR4_X1 port map( A1 => n115627, A2 => n115628, A3 => n115629, A4 
                           => n115630, ZN => n115626);
   U85556 : OAI221_X1 port map( B1 => n114545, B2 => n120164, C1 => n114479, C2
                           => n120158, A => n115638, ZN => n115627);
   U85557 : OAI221_X1 port map( B1 => n99016, B2 => n120188, C1 => n114413, C2 
                           => n120182, A => n115636, ZN => n115628);
   U85558 : OAI221_X1 port map( B1 => n99615, B2 => n120236, C1 => n114022, C2 
                           => n120230, A => n115631, ZN => n115630);
   U85559 : NOR4_X1 port map( A1 => n115599, A2 => n115600, A3 => n115601, A4 
                           => n115602, ZN => n115598);
   U85560 : OAI221_X1 port map( B1 => n114544, B2 => n120164, C1 => n114478, C2
                           => n120158, A => n115610, ZN => n115599);
   U85561 : OAI221_X1 port map( B1 => n99015, B2 => n120188, C1 => n114412, C2 
                           => n120182, A => n115608, ZN => n115600);
   U85562 : OAI221_X1 port map( B1 => n99614, B2 => n120236, C1 => n114021, C2 
                           => n120230, A => n115603, ZN => n115602);
   U85563 : NOR4_X1 port map( A1 => n115571, A2 => n115572, A3 => n115573, A4 
                           => n115574, ZN => n115570);
   U85564 : OAI221_X1 port map( B1 => n114543, B2 => n120164, C1 => n114477, C2
                           => n120158, A => n115582, ZN => n115571);
   U85565 : OAI221_X1 port map( B1 => n99014, B2 => n120188, C1 => n114411, C2 
                           => n120182, A => n115580, ZN => n115572);
   U85566 : OAI221_X1 port map( B1 => n99613, B2 => n120236, C1 => n114020, C2 
                           => n120230, A => n115575, ZN => n115574);
   U85567 : NOR4_X1 port map( A1 => n115543, A2 => n115544, A3 => n115545, A4 
                           => n115546, ZN => n115542);
   U85568 : OAI221_X1 port map( B1 => n114542, B2 => n120164, C1 => n114476, C2
                           => n120158, A => n115554, ZN => n115543);
   U85569 : OAI221_X1 port map( B1 => n99013, B2 => n120188, C1 => n114410, C2 
                           => n120182, A => n115552, ZN => n115544);
   U85570 : OAI221_X1 port map( B1 => n99612, B2 => n120236, C1 => n114019, C2 
                           => n120230, A => n115547, ZN => n115546);
   U85571 : NOR4_X1 port map( A1 => n115515, A2 => n115516, A3 => n115517, A4 
                           => n115518, ZN => n115514);
   U85572 : OAI221_X1 port map( B1 => n114541, B2 => n120164, C1 => n114475, C2
                           => n120158, A => n115526, ZN => n115515);
   U85573 : OAI221_X1 port map( B1 => n99012, B2 => n120188, C1 => n114409, C2 
                           => n120182, A => n115524, ZN => n115516);
   U85574 : OAI221_X1 port map( B1 => n99611, B2 => n120236, C1 => n114018, C2 
                           => n120230, A => n115519, ZN => n115518);
   U85575 : NOR4_X1 port map( A1 => n115487, A2 => n115488, A3 => n115489, A4 
                           => n115490, ZN => n115486);
   U85576 : OAI221_X1 port map( B1 => n114540, B2 => n120164, C1 => n114474, C2
                           => n120158, A => n115498, ZN => n115487);
   U85577 : OAI221_X1 port map( B1 => n99011, B2 => n120188, C1 => n114408, C2 
                           => n120182, A => n115496, ZN => n115488);
   U85578 : OAI221_X1 port map( B1 => n99610, B2 => n120236, C1 => n114017, C2 
                           => n120230, A => n115491, ZN => n115490);
   U85579 : NOR4_X1 port map( A1 => n115459, A2 => n115460, A3 => n115461, A4 
                           => n115462, ZN => n115458);
   U85580 : OAI221_X1 port map( B1 => n114539, B2 => n120164, C1 => n114473, C2
                           => n120158, A => n115470, ZN => n115459);
   U85581 : OAI221_X1 port map( B1 => n99010, B2 => n120188, C1 => n114407, C2 
                           => n120182, A => n115468, ZN => n115460);
   U85582 : OAI221_X1 port map( B1 => n99609, B2 => n120236, C1 => n114016, C2 
                           => n120230, A => n115463, ZN => n115462);
   U85583 : NOR4_X1 port map( A1 => n115431, A2 => n115432, A3 => n115433, A4 
                           => n115434, ZN => n115430);
   U85584 : OAI221_X1 port map( B1 => n114538, B2 => n120165, C1 => n114472, C2
                           => n120159, A => n115442, ZN => n115431);
   U85585 : OAI221_X1 port map( B1 => n99009, B2 => n120189, C1 => n114406, C2 
                           => n120183, A => n115440, ZN => n115432);
   U85586 : OAI221_X1 port map( B1 => n99608, B2 => n120237, C1 => n114015, C2 
                           => n120231, A => n115435, ZN => n115434);
   U85587 : NOR4_X1 port map( A1 => n115403, A2 => n115404, A3 => n115405, A4 
                           => n115406, ZN => n115402);
   U85588 : OAI221_X1 port map( B1 => n114537, B2 => n120165, C1 => n114471, C2
                           => n120159, A => n115414, ZN => n115403);
   U85589 : OAI221_X1 port map( B1 => n99008, B2 => n120189, C1 => n114405, C2 
                           => n120183, A => n115412, ZN => n115404);
   U85590 : OAI221_X1 port map( B1 => n99607, B2 => n120237, C1 => n114014, C2 
                           => n120231, A => n115407, ZN => n115406);
   U85591 : NOR4_X1 port map( A1 => n115375, A2 => n115376, A3 => n115377, A4 
                           => n115378, ZN => n115374);
   U85592 : OAI221_X1 port map( B1 => n114536, B2 => n120165, C1 => n114470, C2
                           => n120159, A => n115386, ZN => n115375);
   U85593 : OAI221_X1 port map( B1 => n99007, B2 => n120189, C1 => n114404, C2 
                           => n120183, A => n115384, ZN => n115376);
   U85594 : OAI221_X1 port map( B1 => n99606, B2 => n120237, C1 => n114013, C2 
                           => n120231, A => n115379, ZN => n115378);
   U85595 : NOR4_X1 port map( A1 => n115347, A2 => n115348, A3 => n115349, A4 
                           => n115350, ZN => n115346);
   U85596 : OAI221_X1 port map( B1 => n114535, B2 => n120165, C1 => n114469, C2
                           => n120159, A => n115358, ZN => n115347);
   U85597 : OAI221_X1 port map( B1 => n99006, B2 => n120189, C1 => n114403, C2 
                           => n120183, A => n115356, ZN => n115348);
   U85598 : OAI221_X1 port map( B1 => n99605, B2 => n120237, C1 => n114012, C2 
                           => n120231, A => n115351, ZN => n115350);
   U85599 : NOR4_X1 port map( A1 => n115319, A2 => n115320, A3 => n115321, A4 
                           => n115322, ZN => n115318);
   U85600 : OAI221_X1 port map( B1 => n114534, B2 => n120165, C1 => n114468, C2
                           => n120159, A => n115330, ZN => n115319);
   U85601 : OAI221_X1 port map( B1 => n99005, B2 => n120189, C1 => n114402, C2 
                           => n120183, A => n115328, ZN => n115320);
   U85602 : OAI221_X1 port map( B1 => n99604, B2 => n120237, C1 => n114011, C2 
                           => n120231, A => n115323, ZN => n115322);
   U85603 : NOR4_X1 port map( A1 => n115291, A2 => n115292, A3 => n115293, A4 
                           => n115294, ZN => n115290);
   U85604 : OAI221_X1 port map( B1 => n114533, B2 => n120165, C1 => n114467, C2
                           => n120159, A => n115302, ZN => n115291);
   U85605 : OAI221_X1 port map( B1 => n99004, B2 => n120189, C1 => n114401, C2 
                           => n120183, A => n115300, ZN => n115292);
   U85606 : OAI221_X1 port map( B1 => n99603, B2 => n120237, C1 => n114010, C2 
                           => n120231, A => n115295, ZN => n115294);
   U85607 : NOR4_X1 port map( A1 => n115263, A2 => n115264, A3 => n115265, A4 
                           => n115266, ZN => n115262);
   U85608 : OAI221_X1 port map( B1 => n114532, B2 => n120165, C1 => n114466, C2
                           => n120159, A => n115274, ZN => n115263);
   U85609 : OAI221_X1 port map( B1 => n99003, B2 => n120189, C1 => n114400, C2 
                           => n120183, A => n115272, ZN => n115264);
   U85610 : OAI221_X1 port map( B1 => n99602, B2 => n120237, C1 => n114009, C2 
                           => n120231, A => n115267, ZN => n115266);
   U85611 : NOR4_X1 port map( A1 => n115235, A2 => n115236, A3 => n115237, A4 
                           => n115238, ZN => n115234);
   U85612 : OAI221_X1 port map( B1 => n114531, B2 => n120165, C1 => n114465, C2
                           => n120159, A => n115246, ZN => n115235);
   U85613 : OAI221_X1 port map( B1 => n99002, B2 => n120189, C1 => n114399, C2 
                           => n120183, A => n115244, ZN => n115236);
   U85614 : OAI221_X1 port map( B1 => n99601, B2 => n120237, C1 => n114008, C2 
                           => n120231, A => n115239, ZN => n115238);
   U85615 : NOR4_X1 port map( A1 => n115207, A2 => n115208, A3 => n115209, A4 
                           => n115210, ZN => n115206);
   U85616 : OAI221_X1 port map( B1 => n114530, B2 => n120165, C1 => n114464, C2
                           => n120159, A => n115218, ZN => n115207);
   U85617 : OAI221_X1 port map( B1 => n99001, B2 => n120189, C1 => n114398, C2 
                           => n120183, A => n115216, ZN => n115208);
   U85618 : OAI221_X1 port map( B1 => n99600, B2 => n120237, C1 => n114007, C2 
                           => n120231, A => n115211, ZN => n115210);
   U85619 : NOR4_X1 port map( A1 => n115179, A2 => n115180, A3 => n115181, A4 
                           => n115182, ZN => n115178);
   U85620 : OAI221_X1 port map( B1 => n114529, B2 => n120165, C1 => n114463, C2
                           => n120159, A => n115190, ZN => n115179);
   U85621 : OAI221_X1 port map( B1 => n99000, B2 => n120189, C1 => n114397, C2 
                           => n120183, A => n115188, ZN => n115180);
   U85622 : OAI221_X1 port map( B1 => n99599, B2 => n120237, C1 => n114006, C2 
                           => n120231, A => n115183, ZN => n115182);
   U85623 : AOI221_X1 port map( B1 => n120089, B2 => n118982, C1 => n120083, C2
                           => n118546, A => n114779, ZN => n114758);
   U85624 : OAI22_X1 port map( A1 => n98718, A2 => n120077, B1 => n99918, B2 =>
                           n120071, ZN => n114779);
   U85625 : AOI221_X1 port map( B1 => n120089, B2 => n118983, C1 => n120083, C2
                           => n118547, A => n114753, ZN => n114732);
   U85626 : OAI22_X1 port map( A1 => n98717, A2 => n120077, B1 => n99917, B2 =>
                           n120071, ZN => n114753);
   U85627 : AOI221_X1 port map( B1 => n120089, B2 => n118984, C1 => n120083, C2
                           => n118548, A => n114727, ZN => n114706);
   U85628 : OAI22_X1 port map( A1 => n98716, A2 => n120077, B1 => n99916, B2 =>
                           n120071, ZN => n114727);
   U85629 : AOI221_X1 port map( B1 => n120089, B2 => n118985, C1 => n120083, C2
                           => n118549, A => n114695, ZN => n114647);
   U85630 : OAI22_X1 port map( A1 => n98714, A2 => n120077, B1 => n99914, B2 =>
                           n120071, ZN => n114695);
   U85631 : AOI221_X1 port map( B1 => n119867, B2 => n95525, C1 => n119861, C2 
                           => n117985, A => n116595, ZN => n116575);
   U85632 : OAI22_X1 port map( A1 => n98652, A2 => n119855, B1 => n99584, B2 =>
                           n119849, ZN => n116595);
   U85633 : AOI221_X1 port map( B1 => n119867, B2 => n95526, C1 => n119861, C2 
                           => n117986, A => n116574, ZN => n116554);
   U85634 : OAI22_X1 port map( A1 => n98651, A2 => n119855, B1 => n99583, B2 =>
                           n119849, ZN => n116574);
   U85635 : AOI221_X1 port map( B1 => n119867, B2 => n95527, C1 => n119861, C2 
                           => n117987, A => n116553, ZN => n116533);
   U85636 : OAI22_X1 port map( A1 => n98650, A2 => n119855, B1 => n99582, B2 =>
                           n119849, ZN => n116553);
   U85637 : AOI221_X1 port map( B1 => n119867, B2 => n95528, C1 => n119861, C2 
                           => n117988, A => n116530, ZN => n116479);
   U85638 : OAI22_X1 port map( A1 => n98648, A2 => n119855, B1 => n99580, B2 =>
                           n119849, ZN => n116530);
   U85639 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), ZN => n113986)
                           ;
   U85640 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n114375, ZN => n113908);
   U85641 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => n114376, ZN => n113913);
   U85642 : OAI221_X1 port map( B1 => n99584, B2 => n120239, C1 => n89969, C2 
                           => n120233, A => n114765, ZN => n114764);
   U85643 : AOI22_X1 port map( A1 => n120227, A2 => n109895, B1 => n120216, B2 
                           => OUT1_60_port, ZN => n114765);
   U85644 : OAI221_X1 port map( B1 => n99583, B2 => n120239, C1 => n89968, C2 
                           => n120233, A => n114739, ZN => n114738);
   U85645 : AOI22_X1 port map( A1 => n120227, A2 => n109896, B1 => n120216, B2 
                           => OUT1_61_port, ZN => n114739);
   U85646 : OAI221_X1 port map( B1 => n99582, B2 => n120239, C1 => n89967, C2 
                           => n120233, A => n114713, ZN => n114712);
   U85647 : AOI22_X1 port map( A1 => n120227, A2 => n109897, B1 => n120216, B2 
                           => OUT1_62_port, ZN => n114713);
   U85648 : OAI221_X1 port map( B1 => n99580, B2 => n120239, C1 => n89965, C2 
                           => n120233, A => n114656, ZN => n114653);
   U85649 : AOI22_X1 port map( A1 => n120227, A2 => n109898, B1 => n120218, B2 
                           => OUT1_63_port, ZN => n114656);
   U85650 : OAI221_X1 port map( B1 => n114448, B2 => n120041, C1 => n99249, C2 
                           => n120035, A => n116583, ZN => n116582);
   U85651 : AOI22_X1 port map( A1 => n120029, A2 => n109903, B1 => n120018, B2 
                           => OUT2_60_port, ZN => n116583);
   U85652 : OAI221_X1 port map( B1 => n114447, B2 => n120041, C1 => n99248, C2 
                           => n120035, A => n116562, ZN => n116561);
   U85653 : AOI22_X1 port map( A1 => n120029, A2 => n109904, B1 => n120018, B2 
                           => OUT2_61_port, ZN => n116562);
   U85654 : OAI221_X1 port map( B1 => n114446, B2 => n120041, C1 => n99247, C2 
                           => n120035, A => n116541, ZN => n116540);
   U85655 : AOI22_X1 port map( A1 => n120029, A2 => n109905, B1 => n120018, B2 
                           => OUT2_62_port, ZN => n116541);
   U85656 : OAI221_X1 port map( B1 => n114444, B2 => n120041, C1 => n99245, C2 
                           => n120035, A => n116489, ZN => n116486);
   U85657 : AOI22_X1 port map( A1 => n120029, A2 => n109906, B1 => n120020, B2 
                           => OUT2_63_port, ZN => n116489);
   U85658 : OAI221_X1 port map( B1 => n114164, B2 => n120213, C1 => n98666, C2 
                           => n120207, A => n115157, ZN => n115153);
   U85659 : AOI22_X1 port map( A1 => n120201, A2 => n118610, B1 => n120195, B2 
                           => n119238, ZN => n115157);
   U85660 : OAI221_X1 port map( B1 => n114163, B2 => n120213, C1 => n98665, C2 
                           => n120207, A => n115129, ZN => n115125);
   U85661 : AOI22_X1 port map( A1 => n120201, A2 => n118611, B1 => n120195, B2 
                           => n119239, ZN => n115129);
   U85662 : OAI221_X1 port map( B1 => n114162, B2 => n120214, C1 => n98664, C2 
                           => n120208, A => n115101, ZN => n115097);
   U85663 : AOI22_X1 port map( A1 => n120202, A2 => n118612, B1 => n120196, B2 
                           => n119240, ZN => n115101);
   U85664 : OAI221_X1 port map( B1 => n114161, B2 => n120214, C1 => n98663, C2 
                           => n120208, A => n115073, ZN => n115069);
   U85665 : AOI22_X1 port map( A1 => n120202, A2 => n118613, B1 => n120196, B2 
                           => n119241, ZN => n115073);
   U85666 : OAI221_X1 port map( B1 => n114160, B2 => n120214, C1 => n98662, C2 
                           => n120208, A => n115045, ZN => n115041);
   U85667 : AOI22_X1 port map( A1 => n120202, A2 => n118614, B1 => n120196, B2 
                           => n119242, ZN => n115045);
   U85668 : OAI221_X1 port map( B1 => n114159, B2 => n120214, C1 => n98661, C2 
                           => n120208, A => n115017, ZN => n115013);
   U85669 : AOI22_X1 port map( A1 => n120202, A2 => n118615, B1 => n120196, B2 
                           => n119243, ZN => n115017);
   U85670 : OAI221_X1 port map( B1 => n114158, B2 => n120214, C1 => n98660, C2 
                           => n120208, A => n114989, ZN => n114985);
   U85671 : AOI22_X1 port map( A1 => n120202, A2 => n118616, B1 => n120196, B2 
                           => n119244, ZN => n114989);
   U85672 : OAI221_X1 port map( B1 => n114157, B2 => n120214, C1 => n98659, C2 
                           => n120208, A => n114961, ZN => n114957);
   U85673 : AOI22_X1 port map( A1 => n120202, A2 => n118617, B1 => n120196, B2 
                           => n119245, ZN => n114961);
   U85674 : OAI221_X1 port map( B1 => n114156, B2 => n120214, C1 => n98658, C2 
                           => n120208, A => n114933, ZN => n114929);
   U85675 : AOI22_X1 port map( A1 => n120202, A2 => n118618, B1 => n120196, B2 
                           => n119246, ZN => n114933);
   U85676 : OAI221_X1 port map( B1 => n114155, B2 => n120214, C1 => n98657, C2 
                           => n120208, A => n114905, ZN => n114901);
   U85677 : AOI22_X1 port map( A1 => n120202, A2 => n118619, B1 => n120196, B2 
                           => n119247, ZN => n114905);
   U85678 : OAI221_X1 port map( B1 => n114154, B2 => n120214, C1 => n98656, C2 
                           => n120208, A => n114877, ZN => n114873);
   U85679 : AOI22_X1 port map( A1 => n120202, A2 => n118620, B1 => n120196, B2 
                           => n119248, ZN => n114877);
   U85680 : OAI221_X1 port map( B1 => n114153, B2 => n120214, C1 => n98655, C2 
                           => n120208, A => n114849, ZN => n114845);
   U85681 : AOI22_X1 port map( A1 => n120202, A2 => n118621, B1 => n120196, B2 
                           => n119249, ZN => n114849);
   U85682 : OAI221_X1 port map( B1 => n114152, B2 => n120214, C1 => n98654, C2 
                           => n120208, A => n114821, ZN => n114817);
   U85683 : AOI22_X1 port map( A1 => n120202, A2 => n118622, B1 => n120196, B2 
                           => n119250, ZN => n114821);
   U85684 : OAI221_X1 port map( B1 => n114151, B2 => n120214, C1 => n98653, C2 
                           => n120208, A => n114793, ZN => n114789);
   U85685 : AOI22_X1 port map( A1 => n120202, A2 => n118623, B1 => n120196, B2 
                           => n119251, ZN => n114793);
   U85686 : OAI221_X1 port map( B1 => n114198, B2 => n120211, C1 => n98700, C2 
                           => n120205, A => n116109, ZN => n116105);
   U85687 : AOI22_X1 port map( A1 => n120199, A2 => n118624, B1 => n120193, B2 
                           => n119252, ZN => n116109);
   U85688 : OAI221_X1 port map( B1 => n114197, B2 => n120211, C1 => n98699, C2 
                           => n120205, A => n116081, ZN => n116077);
   U85689 : AOI22_X1 port map( A1 => n120199, A2 => n118625, B1 => n120193, B2 
                           => n119253, ZN => n116081);
   U85690 : OAI221_X1 port map( B1 => n114196, B2 => n120211, C1 => n98698, C2 
                           => n120205, A => n116053, ZN => n116049);
   U85691 : AOI22_X1 port map( A1 => n120199, A2 => n118626, B1 => n120193, B2 
                           => n119254, ZN => n116053);
   U85692 : OAI221_X1 port map( B1 => n114195, B2 => n120211, C1 => n98697, C2 
                           => n120205, A => n116025, ZN => n116021);
   U85693 : AOI22_X1 port map( A1 => n120199, A2 => n118627, B1 => n120193, B2 
                           => n119255, ZN => n116025);
   U85694 : OAI221_X1 port map( B1 => n114194, B2 => n120211, C1 => n98696, C2 
                           => n120205, A => n115997, ZN => n115993);
   U85695 : AOI22_X1 port map( A1 => n120199, A2 => n118628, B1 => n120193, B2 
                           => n119256, ZN => n115997);
   U85696 : OAI221_X1 port map( B1 => n114193, B2 => n120211, C1 => n98695, C2 
                           => n120205, A => n115969, ZN => n115965);
   U85697 : AOI22_X1 port map( A1 => n120199, A2 => n118629, B1 => n120193, B2 
                           => n119257, ZN => n115969);
   U85698 : OAI221_X1 port map( B1 => n114192, B2 => n120211, C1 => n98694, C2 
                           => n120205, A => n115941, ZN => n115937);
   U85699 : AOI22_X1 port map( A1 => n120199, A2 => n118630, B1 => n120193, B2 
                           => n119258, ZN => n115941);
   U85700 : OAI221_X1 port map( B1 => n114191, B2 => n120211, C1 => n98693, C2 
                           => n120205, A => n115913, ZN => n115909);
   U85701 : AOI22_X1 port map( A1 => n120199, A2 => n118631, B1 => n120193, B2 
                           => n119259, ZN => n115913);
   U85702 : OAI221_X1 port map( B1 => n114190, B2 => n120211, C1 => n98692, C2 
                           => n120205, A => n115885, ZN => n115881);
   U85703 : AOI22_X1 port map( A1 => n120199, A2 => n118632, B1 => n120193, B2 
                           => n119260, ZN => n115885);
   U85704 : OAI221_X1 port map( B1 => n114189, B2 => n120211, C1 => n98691, C2 
                           => n120205, A => n115857, ZN => n115853);
   U85705 : AOI22_X1 port map( A1 => n120199, A2 => n118633, B1 => n120193, B2 
                           => n119261, ZN => n115857);
   U85706 : OAI221_X1 port map( B1 => n114188, B2 => n120211, C1 => n98690, C2 
                           => n120205, A => n115829, ZN => n115825);
   U85707 : AOI22_X1 port map( A1 => n120199, A2 => n118634, B1 => n120193, B2 
                           => n119262, ZN => n115829);
   U85708 : OAI221_X1 port map( B1 => n114187, B2 => n120211, C1 => n98689, C2 
                           => n120205, A => n115801, ZN => n115797);
   U85709 : AOI22_X1 port map( A1 => n120199, A2 => n118635, B1 => n120193, B2 
                           => n119263, ZN => n115801);
   U85710 : OAI221_X1 port map( B1 => n114186, B2 => n120212, C1 => n98688, C2 
                           => n120206, A => n115773, ZN => n115769);
   U85711 : AOI22_X1 port map( A1 => n120200, A2 => n118636, B1 => n120194, B2 
                           => n119264, ZN => n115773);
   U85712 : OAI221_X1 port map( B1 => n114185, B2 => n120212, C1 => n98687, C2 
                           => n120206, A => n115745, ZN => n115741);
   U85713 : AOI22_X1 port map( A1 => n120200, A2 => n118637, B1 => n120194, B2 
                           => n119265, ZN => n115745);
   U85714 : OAI221_X1 port map( B1 => n114184, B2 => n120212, C1 => n98686, C2 
                           => n120206, A => n115717, ZN => n115713);
   U85715 : AOI22_X1 port map( A1 => n120200, A2 => n118638, B1 => n120194, B2 
                           => n119266, ZN => n115717);
   U85716 : OAI221_X1 port map( B1 => n114183, B2 => n120212, C1 => n98685, C2 
                           => n120206, A => n115689, ZN => n115685);
   U85717 : AOI22_X1 port map( A1 => n120200, A2 => n118639, B1 => n120194, B2 
                           => n119267, ZN => n115689);
   U85718 : OAI221_X1 port map( B1 => n114182, B2 => n120212, C1 => n98684, C2 
                           => n120206, A => n115661, ZN => n115657);
   U85719 : AOI22_X1 port map( A1 => n120200, A2 => n118640, B1 => n120194, B2 
                           => n119268, ZN => n115661);
   U85720 : OAI221_X1 port map( B1 => n114181, B2 => n120212, C1 => n98683, C2 
                           => n120206, A => n115633, ZN => n115629);
   U85721 : AOI22_X1 port map( A1 => n120200, A2 => n118641, B1 => n120194, B2 
                           => n119269, ZN => n115633);
   U85722 : OAI221_X1 port map( B1 => n114180, B2 => n120212, C1 => n98682, C2 
                           => n120206, A => n115605, ZN => n115601);
   U85723 : AOI22_X1 port map( A1 => n120200, A2 => n118642, B1 => n120194, B2 
                           => n119270, ZN => n115605);
   U85724 : OAI221_X1 port map( B1 => n114179, B2 => n120212, C1 => n98681, C2 
                           => n120206, A => n115577, ZN => n115573);
   U85725 : AOI22_X1 port map( A1 => n120200, A2 => n118643, B1 => n120194, B2 
                           => n119271, ZN => n115577);
   U85726 : OAI221_X1 port map( B1 => n114178, B2 => n120212, C1 => n98680, C2 
                           => n120206, A => n115549, ZN => n115545);
   U85727 : AOI22_X1 port map( A1 => n120200, A2 => n118644, B1 => n120194, B2 
                           => n119272, ZN => n115549);
   U85728 : OAI221_X1 port map( B1 => n114177, B2 => n120212, C1 => n98679, C2 
                           => n120206, A => n115521, ZN => n115517);
   U85729 : AOI22_X1 port map( A1 => n120200, A2 => n118645, B1 => n120194, B2 
                           => n119273, ZN => n115521);
   U85730 : OAI221_X1 port map( B1 => n114176, B2 => n120212, C1 => n98678, C2 
                           => n120206, A => n115493, ZN => n115489);
   U85731 : AOI22_X1 port map( A1 => n120200, A2 => n118646, B1 => n120194, B2 
                           => n119274, ZN => n115493);
   U85732 : OAI221_X1 port map( B1 => n114175, B2 => n120212, C1 => n98677, C2 
                           => n120206, A => n115465, ZN => n115461);
   U85733 : AOI22_X1 port map( A1 => n120200, A2 => n118647, B1 => n120194, B2 
                           => n119275, ZN => n115465);
   U85734 : OAI221_X1 port map( B1 => n114174, B2 => n120213, C1 => n98676, C2 
                           => n120207, A => n115437, ZN => n115433);
   U85735 : AOI22_X1 port map( A1 => n120201, A2 => n118648, B1 => n120195, B2 
                           => n119276, ZN => n115437);
   U85736 : OAI221_X1 port map( B1 => n114173, B2 => n120213, C1 => n98675, C2 
                           => n120207, A => n115409, ZN => n115405);
   U85737 : AOI22_X1 port map( A1 => n120201, A2 => n118649, B1 => n120195, B2 
                           => n119277, ZN => n115409);
   U85738 : OAI221_X1 port map( B1 => n114172, B2 => n120213, C1 => n98674, C2 
                           => n120207, A => n115381, ZN => n115377);
   U85739 : AOI22_X1 port map( A1 => n120201, A2 => n118650, B1 => n120195, B2 
                           => n119278, ZN => n115381);
   U85740 : OAI221_X1 port map( B1 => n114171, B2 => n120213, C1 => n98673, C2 
                           => n120207, A => n115353, ZN => n115349);
   U85741 : AOI22_X1 port map( A1 => n120201, A2 => n118651, B1 => n120195, B2 
                           => n119279, ZN => n115353);
   U85742 : OAI221_X1 port map( B1 => n114170, B2 => n120213, C1 => n98672, C2 
                           => n120207, A => n115325, ZN => n115321);
   U85743 : AOI22_X1 port map( A1 => n120201, A2 => n118652, B1 => n120195, B2 
                           => n119280, ZN => n115325);
   U85744 : OAI221_X1 port map( B1 => n114169, B2 => n120213, C1 => n98671, C2 
                           => n120207, A => n115297, ZN => n115293);
   U85745 : AOI22_X1 port map( A1 => n120201, A2 => n118653, B1 => n120195, B2 
                           => n119281, ZN => n115297);
   U85746 : OAI221_X1 port map( B1 => n114168, B2 => n120213, C1 => n98670, C2 
                           => n120207, A => n115269, ZN => n115265);
   U85747 : AOI22_X1 port map( A1 => n120201, A2 => n118654, B1 => n120195, B2 
                           => n119282, ZN => n115269);
   U85748 : OAI221_X1 port map( B1 => n114167, B2 => n120213, C1 => n98669, C2 
                           => n120207, A => n115241, ZN => n115237);
   U85749 : AOI22_X1 port map( A1 => n120201, A2 => n118655, B1 => n120195, B2 
                           => n119283, ZN => n115241);
   U85750 : OAI221_X1 port map( B1 => n114166, B2 => n120213, C1 => n98668, C2 
                           => n120207, A => n115213, ZN => n115209);
   U85751 : AOI22_X1 port map( A1 => n120201, A2 => n118656, B1 => n120195, B2 
                           => n119284, ZN => n115213);
   U85752 : OAI221_X1 port map( B1 => n114165, B2 => n120213, C1 => n98667, C2 
                           => n120207, A => n115185, ZN => n115181);
   U85753 : AOI22_X1 port map( A1 => n120201, A2 => n118657, B1 => n120195, B2 
                           => n119285, ZN => n115185);
   U85754 : OAI221_X1 port map( B1 => n114210, B2 => n120210, C1 => n98712, C2 
                           => n120204, A => n116449, ZN => n116441);
   U85755 : AOI22_X1 port map( A1 => n120198, A2 => n118658, B1 => n120192, B2 
                           => n119286, ZN => n116449);
   U85756 : OAI221_X1 port map( B1 => n114209, B2 => n120210, C1 => n98711, C2 
                           => n120204, A => n116417, ZN => n116413);
   U85757 : AOI22_X1 port map( A1 => n120198, A2 => n118659, B1 => n120192, B2 
                           => n119287, ZN => n116417);
   U85758 : OAI221_X1 port map( B1 => n114208, B2 => n120210, C1 => n98710, C2 
                           => n120204, A => n116389, ZN => n116385);
   U85759 : AOI22_X1 port map( A1 => n120198, A2 => n118660, B1 => n120192, B2 
                           => n119288, ZN => n116389);
   U85760 : OAI221_X1 port map( B1 => n114207, B2 => n120210, C1 => n98709, C2 
                           => n120204, A => n116361, ZN => n116357);
   U85761 : AOI22_X1 port map( A1 => n120198, A2 => n118661, B1 => n120192, B2 
                           => n119289, ZN => n116361);
   U85762 : OAI221_X1 port map( B1 => n114206, B2 => n120210, C1 => n98708, C2 
                           => n120204, A => n116333, ZN => n116329);
   U85763 : AOI22_X1 port map( A1 => n120198, A2 => n118662, B1 => n120192, B2 
                           => n119290, ZN => n116333);
   U85764 : OAI221_X1 port map( B1 => n114205, B2 => n120210, C1 => n98707, C2 
                           => n120204, A => n116305, ZN => n116301);
   U85765 : AOI22_X1 port map( A1 => n120198, A2 => n118663, B1 => n120192, B2 
                           => n119291, ZN => n116305);
   U85766 : OAI221_X1 port map( B1 => n114204, B2 => n120210, C1 => n98706, C2 
                           => n120204, A => n116277, ZN => n116273);
   U85767 : AOI22_X1 port map( A1 => n120198, A2 => n118664, B1 => n120192, B2 
                           => n119292, ZN => n116277);
   U85768 : OAI221_X1 port map( B1 => n114203, B2 => n120210, C1 => n98705, C2 
                           => n120204, A => n116249, ZN => n116245);
   U85769 : AOI22_X1 port map( A1 => n120198, A2 => n118665, B1 => n120192, B2 
                           => n119293, ZN => n116249);
   U85770 : OAI221_X1 port map( B1 => n114202, B2 => n120210, C1 => n98704, C2 
                           => n120204, A => n116221, ZN => n116217);
   U85771 : AOI22_X1 port map( A1 => n120198, A2 => n118666, B1 => n120192, B2 
                           => n119294, ZN => n116221);
   U85772 : OAI221_X1 port map( B1 => n114201, B2 => n120210, C1 => n98703, C2 
                           => n120204, A => n116193, ZN => n116189);
   U85773 : AOI22_X1 port map( A1 => n120198, A2 => n118667, B1 => n120192, B2 
                           => n119295, ZN => n116193);
   U85774 : OAI221_X1 port map( B1 => n114200, B2 => n120210, C1 => n98702, C2 
                           => n120204, A => n116165, ZN => n116161);
   U85775 : AOI22_X1 port map( A1 => n120198, A2 => n118668, B1 => n120192, B2 
                           => n119296, ZN => n116165);
   U85776 : OAI221_X1 port map( B1 => n114199, B2 => n120210, C1 => n98701, C2 
                           => n120204, A => n116137, ZN => n116133);
   U85777 : AOI22_X1 port map( A1 => n120198, A2 => n118669, B1 => n120192, B2 
                           => n119297, ZN => n116137);
   U85778 : OAI221_X1 port map( B1 => n114127, B2 => n120191, C1 => n114382, C2
                           => n120185, A => n114769, ZN => n114762);
   U85779 : AOI22_X1 port map( A1 => n120179, A2 => n117974, B1 => n120173, B2 
                           => n119110, ZN => n114769);
   U85780 : OAI221_X1 port map( B1 => n114126, B2 => n120191, C1 => n114381, C2
                           => n120185, A => n114743, ZN => n114736);
   U85781 : AOI22_X1 port map( A1 => n120179, A2 => n117975, B1 => n120173, B2 
                           => n119111, ZN => n114743);
   U85782 : OAI221_X1 port map( B1 => n114125, B2 => n120191, C1 => n114380, C2
                           => n120185, A => n114717, ZN => n114710);
   U85783 : AOI22_X1 port map( A1 => n120179, A2 => n117976, B1 => n120173, B2 
                           => n119112, ZN => n114717);
   U85784 : OAI221_X1 port map( B1 => n114123, B2 => n120191, C1 => n114378, C2
                           => n120185, A => n114668, ZN => n114651);
   U85785 : AOI22_X1 port map( A1 => n120179, A2 => n117977, B1 => n120173, B2 
                           => n119113, ZN => n114668);
   U85786 : OAI221_X1 port map( B1 => n114514, B2 => n119993, C1 => n114150, C2
                           => n119987, A => n116587, ZN => n116580);
   U85787 : AOI22_X1 port map( A1 => n119981, A2 => n111041, B1 => n119975, B2 
                           => n117993, ZN => n116587);
   U85788 : OAI221_X1 port map( B1 => n114513, B2 => n119993, C1 => n114149, C2
                           => n119987, A => n116566, ZN => n116559);
   U85789 : AOI22_X1 port map( A1 => n119981, A2 => n111042, B1 => n119975, B2 
                           => n117994, ZN => n116566);
   U85790 : OAI221_X1 port map( B1 => n114512, B2 => n119993, C1 => n114148, C2
                           => n119987, A => n116545, ZN => n116538);
   U85791 : AOI22_X1 port map( A1 => n119981, A2 => n111043, B1 => n119975, B2 
                           => n117995, ZN => n116545);
   U85792 : OAI221_X1 port map( B1 => n114510, B2 => n119993, C1 => n114146, C2
                           => n119987, A => n116501, ZN => n116484);
   U85793 : AOI22_X1 port map( A1 => n119981, A2 => n111044, B1 => n119975, B2 
                           => n117996, ZN => n116501);
   U85794 : OAI221_X1 port map( B1 => n114514, B2 => n120167, C1 => n114448, C2
                           => n120161, A => n114771, ZN => n114761);
   U85795 : AOI22_X1 port map( A1 => n120155, A2 => n111045, B1 => n120149, B2 
                           => n119046, ZN => n114771);
   U85796 : OAI221_X1 port map( B1 => n114513, B2 => n120167, C1 => n114447, C2
                           => n120161, A => n114745, ZN => n114735);
   U85797 : AOI22_X1 port map( A1 => n120155, A2 => n111046, B1 => n120149, B2 
                           => n119047, ZN => n114745);
   U85798 : OAI221_X1 port map( B1 => n114512, B2 => n120167, C1 => n114446, C2
                           => n120161, A => n114719, ZN => n114709);
   U85799 : AOI22_X1 port map( A1 => n120155, A2 => n111047, B1 => n120149, B2 
                           => n119048, ZN => n114719);
   U85800 : OAI221_X1 port map( B1 => n114510, B2 => n120167, C1 => n114444, C2
                           => n120161, A => n114674, ZN => n114650);
   U85801 : AOI22_X1 port map( A1 => n120155, A2 => n111048, B1 => n120149, B2 
                           => n119049, ZN => n114674);
   U85802 : OAI221_X1 port map( B1 => n99183, B2 => n119969, C1 => n113985, C2 
                           => n119963, A => n116588, ZN => n116579);
   U85803 : AOI22_X1 port map( A1 => n119957, A2 => n117981, B1 => n119951, B2 
                           => n117974, ZN => n116588);
   U85804 : OAI221_X1 port map( B1 => n99182, B2 => n119969, C1 => n113984, C2 
                           => n119963, A => n116567, ZN => n116558);
   U85805 : AOI22_X1 port map( A1 => n119957, A2 => n117982, B1 => n119951, B2 
                           => n117975, ZN => n116567);
   U85806 : OAI221_X1 port map( B1 => n99181, B2 => n119969, C1 => n113983, C2 
                           => n119963, A => n116546, ZN => n116537);
   U85807 : AOI22_X1 port map( A1 => n119957, A2 => n117983, B1 => n119951, B2 
                           => n117976, ZN => n116546);
   U85808 : OAI221_X1 port map( B1 => n99179, B2 => n119969, C1 => n113981, C2 
                           => n119963, A => n116506, ZN => n116483);
   U85809 : AOI22_X1 port map( A1 => n119957, A2 => n117984, B1 => n119951, B2 
                           => n117977, ZN => n116506);
   U85810 : OAI22_X1 port map( A1 => n99051, A2 => n120143, B1 => n89500, B2 =>
                           n120137, ZN => n114776);
   U85811 : OAI22_X1 port map( A1 => n99050, A2 => n120143, B1 => n89498, B2 =>
                           n120137, ZN => n114750);
   U85812 : OAI22_X1 port map( A1 => n99049, A2 => n120143, B1 => n89496, B2 =>
                           n120137, ZN => n114724);
   U85813 : OAI22_X1 port map( A1 => n99047, A2 => n120143, B1 => n89493, B2 =>
                           n120137, ZN => n114681);
   U85814 : OAI22_X1 port map( A1 => n99720, A2 => n119945, B1 => n89500, B2 =>
                           n119939, ZN => n116592);
   U85815 : OAI22_X1 port map( A1 => n99719, A2 => n119945, B1 => n89498, B2 =>
                           n119939, ZN => n116571);
   U85816 : OAI22_X1 port map( A1 => n99718, A2 => n119945, B1 => n89496, B2 =>
                           n119939, ZN => n116550);
   U85817 : OAI22_X1 port map( A1 => n99716, A2 => n119945, B1 => n89493, B2 =>
                           n119939, ZN => n116512);
   U85818 : OAI22_X1 port map( A1 => n90310, A2 => n120131, B1 => n114239, B2 
                           => n120125, ZN => n114775);
   U85819 : OAI22_X1 port map( A1 => n90309, A2 => n120131, B1 => n114238, B2 
                           => n120125, ZN => n114749);
   U85820 : OAI22_X1 port map( A1 => n90308, A2 => n120131, B1 => n114237, B2 
                           => n120125, ZN => n114723);
   U85821 : OAI22_X1 port map( A1 => n90306, A2 => n120131, B1 => n114235, B2 
                           => n120125, ZN => n114680);
   U85822 : OAI22_X1 port map( A1 => n90715, A2 => n119933, B1 => n99051, B2 =>
                           n119927, ZN => n116591);
   U85823 : OAI22_X1 port map( A1 => n90714, A2 => n119933, B1 => n99050, B2 =>
                           n119927, ZN => n116570);
   U85824 : OAI22_X1 port map( A1 => n90713, A2 => n119933, B1 => n99049, B2 =>
                           n119927, ZN => n116549);
   U85825 : OAI22_X1 port map( A1 => n90711, A2 => n119933, B1 => n99047, B2 =>
                           n119927, ZN => n116511);
   U85826 : OAI22_X1 port map( A1 => n89969, A2 => n119879, B1 => n99450, B2 =>
                           n119873, ZN => n116594);
   U85827 : OAI22_X1 port map( A1 => n89968, A2 => n119879, B1 => n99449, B2 =>
                           n119873, ZN => n116573);
   U85828 : OAI22_X1 port map( A1 => n89967, A2 => n119879, B1 => n99448, B2 =>
                           n119873, ZN => n116552);
   U85829 : OAI22_X1 port map( A1 => n89965, A2 => n119879, B1 => n99446, B2 =>
                           n119873, ZN => n116525);
   U85830 : OAI22_X1 port map( A1 => n90516, A2 => n120119, B1 => n90035, B2 =>
                           n120113, ZN => n114774);
   U85831 : OAI22_X1 port map( A1 => n90515, A2 => n120119, B1 => n90034, B2 =>
                           n120113, ZN => n114748);
   U85832 : OAI22_X1 port map( A1 => n90514, A2 => n120119, B1 => n90033, B2 =>
                           n120113, ZN => n114722);
   U85833 : OAI22_X1 port map( A1 => n90512, A2 => n120119, B1 => n90031, B2 =>
                           n120113, ZN => n114679);
   U85834 : OAI22_X1 port map( A1 => n98718, A2 => n119921, B1 => n90377, B2 =>
                           n119915, ZN => n116590);
   U85835 : OAI22_X1 port map( A1 => n98717, A2 => n119921, B1 => n90376, B2 =>
                           n119915, ZN => n116569);
   U85836 : OAI22_X1 port map( A1 => n98716, A2 => n119921, B1 => n90375, B2 =>
                           n119915, ZN => n116548);
   U85837 : OAI22_X1 port map( A1 => n98714, A2 => n119921, B1 => n90373, B2 =>
                           n119915, ZN => n116510);
   U85838 : OAI22_X1 port map( A1 => n90764, A2 => n119928, B1 => n99100, B2 =>
                           n119922, ZN => n117711);
   U85839 : OAI22_X1 port map( A1 => n90763, A2 => n119929, B1 => n99099, B2 =>
                           n119923, ZN => n117689);
   U85840 : OAI22_X1 port map( A1 => n90762, A2 => n119929, B1 => n99098, B2 =>
                           n119923, ZN => n117667);
   U85841 : OAI22_X1 port map( A1 => n90761, A2 => n119929, B1 => n99097, B2 =>
                           n119923, ZN => n117645);
   U85842 : OAI22_X1 port map( A1 => n90760, A2 => n119929, B1 => n99096, B2 =>
                           n119923, ZN => n117623);
   U85843 : OAI22_X1 port map( A1 => n90759, A2 => n119929, B1 => n99095, B2 =>
                           n119923, ZN => n117601);
   U85844 : OAI22_X1 port map( A1 => n90758, A2 => n119929, B1 => n99094, B2 =>
                           n119923, ZN => n117579);
   U85845 : OAI22_X1 port map( A1 => n90757, A2 => n119929, B1 => n99093, B2 =>
                           n119923, ZN => n117557);
   U85846 : OAI22_X1 port map( A1 => n90756, A2 => n119929, B1 => n99092, B2 =>
                           n119923, ZN => n117534);
   U85847 : OAI22_X1 port map( A1 => n90755, A2 => n119929, B1 => n99091, B2 =>
                           n119923, ZN => n117511);
   U85848 : OAI22_X1 port map( A1 => n90754, A2 => n119929, B1 => n99090, B2 =>
                           n119923, ZN => n117488);
   U85849 : OAI22_X1 port map( A1 => n90753, A2 => n119929, B1 => n99089, B2 =>
                           n119923, ZN => n117465);
   U85850 : OAI22_X1 port map( A1 => n90752, A2 => n119929, B1 => n99088, B2 =>
                           n119923, ZN => n117442);
   U85851 : OAI22_X1 port map( A1 => n90751, A2 => n119930, B1 => n99087, B2 =>
                           n119924, ZN => n117419);
   U85852 : OAI22_X1 port map( A1 => n90750, A2 => n119930, B1 => n99086, B2 =>
                           n119924, ZN => n117396);
   U85853 : OAI22_X1 port map( A1 => n90749, A2 => n119930, B1 => n99085, B2 =>
                           n119924, ZN => n117373);
   U85854 : OAI22_X1 port map( A1 => n90748, A2 => n119930, B1 => n99084, B2 =>
                           n119924, ZN => n117350);
   U85855 : OAI22_X1 port map( A1 => n90747, A2 => n119930, B1 => n99083, B2 =>
                           n119924, ZN => n117327);
   U85856 : OAI22_X1 port map( A1 => n90746, A2 => n119930, B1 => n99082, B2 =>
                           n119924, ZN => n117304);
   U85857 : OAI22_X1 port map( A1 => n90745, A2 => n119930, B1 => n99081, B2 =>
                           n119924, ZN => n117281);
   U85858 : OAI22_X1 port map( A1 => n90744, A2 => n119930, B1 => n99080, B2 =>
                           n119924, ZN => n117258);
   U85859 : OAI22_X1 port map( A1 => n90743, A2 => n119930, B1 => n99079, B2 =>
                           n119924, ZN => n117235);
   U85860 : OAI22_X1 port map( A1 => n90742, A2 => n119930, B1 => n99078, B2 =>
                           n119924, ZN => n117212);
   U85861 : OAI22_X1 port map( A1 => n90741, A2 => n119930, B1 => n99077, B2 =>
                           n119924, ZN => n117189);
   U85862 : OAI22_X1 port map( A1 => n90740, A2 => n119930, B1 => n99076, B2 =>
                           n119924, ZN => n117166);
   U85863 : OAI22_X1 port map( A1 => n90739, A2 => n119931, B1 => n99075, B2 =>
                           n119925, ZN => n117143);
   U85864 : OAI22_X1 port map( A1 => n90738, A2 => n119931, B1 => n99074, B2 =>
                           n119925, ZN => n117120);
   U85865 : OAI22_X1 port map( A1 => n90737, A2 => n119931, B1 => n99073, B2 =>
                           n119925, ZN => n117097);
   U85866 : OAI22_X1 port map( A1 => n90736, A2 => n119931, B1 => n99072, B2 =>
                           n119925, ZN => n117074);
   U85867 : OAI22_X1 port map( A1 => n90735, A2 => n119931, B1 => n99071, B2 =>
                           n119925, ZN => n117051);
   U85868 : OAI22_X1 port map( A1 => n90734, A2 => n119931, B1 => n99070, B2 =>
                           n119925, ZN => n117028);
   U85869 : OAI22_X1 port map( A1 => n90733, A2 => n119931, B1 => n99069, B2 =>
                           n119925, ZN => n117005);
   U85870 : OAI22_X1 port map( A1 => n90732, A2 => n119931, B1 => n99068, B2 =>
                           n119925, ZN => n116982);
   U85871 : OAI22_X1 port map( A1 => n90731, A2 => n119931, B1 => n99067, B2 =>
                           n119925, ZN => n116959);
   U85872 : OAI22_X1 port map( A1 => n90730, A2 => n119931, B1 => n99066, B2 =>
                           n119925, ZN => n116936);
   U85873 : OAI22_X1 port map( A1 => n90729, A2 => n119931, B1 => n99065, B2 =>
                           n119925, ZN => n116913);
   U85874 : OAI22_X1 port map( A1 => n90728, A2 => n119931, B1 => n99064, B2 =>
                           n119925, ZN => n116890);
   U85875 : OAI22_X1 port map( A1 => n90727, A2 => n119932, B1 => n99063, B2 =>
                           n119926, ZN => n116867);
   U85876 : OAI22_X1 port map( A1 => n90726, A2 => n119932, B1 => n99062, B2 =>
                           n119926, ZN => n116844);
   U85877 : OAI22_X1 port map( A1 => n90725, A2 => n119932, B1 => n99061, B2 =>
                           n119926, ZN => n116821);
   U85878 : OAI22_X1 port map( A1 => n90724, A2 => n119932, B1 => n99060, B2 =>
                           n119926, ZN => n116798);
   U85879 : OAI22_X1 port map( A1 => n90723, A2 => n119932, B1 => n99059, B2 =>
                           n119926, ZN => n116775);
   U85880 : OAI22_X1 port map( A1 => n90722, A2 => n119932, B1 => n99058, B2 =>
                           n119926, ZN => n116752);
   U85881 : OAI22_X1 port map( A1 => n90721, A2 => n119932, B1 => n99057, B2 =>
                           n119926, ZN => n116729);
   U85882 : OAI22_X1 port map( A1 => n90720, A2 => n119932, B1 => n99056, B2 =>
                           n119926, ZN => n116706);
   U85883 : OAI22_X1 port map( A1 => n90719, A2 => n119932, B1 => n99055, B2 =>
                           n119926, ZN => n116683);
   U85884 : OAI22_X1 port map( A1 => n90718, A2 => n119932, B1 => n99054, B2 =>
                           n119926, ZN => n116660);
   U85885 : OAI22_X1 port map( A1 => n90717, A2 => n119932, B1 => n99053, B2 =>
                           n119926, ZN => n116637);
   U85886 : OAI22_X1 port map( A1 => n90716, A2 => n119932, B1 => n99052, B2 =>
                           n119926, ZN => n116614);
   U85887 : OAI22_X1 port map( A1 => n90768, A2 => n119928, B1 => n99104, B2 =>
                           n119922, ZN => n117799);
   U85888 : OAI22_X1 port map( A1 => n90767, A2 => n119928, B1 => n99103, B2 =>
                           n119922, ZN => n117777);
   U85889 : OAI22_X1 port map( A1 => n90766, A2 => n119928, B1 => n99102, B2 =>
                           n119922, ZN => n117755);
   U85890 : OAI22_X1 port map( A1 => n90765, A2 => n119928, B1 => n99101, B2 =>
                           n119922, ZN => n117733);
   U85891 : OAI22_X1 port map( A1 => n90775, A2 => n119928, B1 => n99111, B2 =>
                           n119922, ZN => n117965);
   U85892 : OAI22_X1 port map( A1 => n90774, A2 => n119928, B1 => n99110, B2 =>
                           n119922, ZN => n117931);
   U85893 : OAI22_X1 port map( A1 => n90773, A2 => n119928, B1 => n99109, B2 =>
                           n119922, ZN => n117909);
   U85894 : OAI22_X1 port map( A1 => n90772, A2 => n119928, B1 => n99108, B2 =>
                           n119922, ZN => n117887);
   U85895 : OAI22_X1 port map( A1 => n90771, A2 => n119928, B1 => n99107, B2 =>
                           n119922, ZN => n117865);
   U85896 : OAI22_X1 port map( A1 => n90770, A2 => n119928, B1 => n99106, B2 =>
                           n119922, ZN => n117843);
   U85897 : OAI22_X1 port map( A1 => n90769, A2 => n119928, B1 => n99105, B2 =>
                           n119922, ZN => n117821);
   U85898 : OAI22_X1 port map( A1 => n98701, A2 => n119850, B1 => n99633, B2 =>
                           n119844, ZN => n117714);
   U85899 : OAI22_X1 port map( A1 => n98700, A2 => n119851, B1 => n99632, B2 =>
                           n119845, ZN => n117692);
   U85900 : OAI22_X1 port map( A1 => n98699, A2 => n119851, B1 => n99631, B2 =>
                           n119845, ZN => n117670);
   U85901 : OAI22_X1 port map( A1 => n98698, A2 => n119851, B1 => n99630, B2 =>
                           n119845, ZN => n117648);
   U85902 : OAI22_X1 port map( A1 => n98697, A2 => n119851, B1 => n99629, B2 =>
                           n119845, ZN => n117626);
   U85903 : OAI22_X1 port map( A1 => n98696, A2 => n119851, B1 => n99628, B2 =>
                           n119845, ZN => n117604);
   U85904 : OAI22_X1 port map( A1 => n98695, A2 => n119851, B1 => n99627, B2 =>
                           n119845, ZN => n117582);
   U85905 : OAI22_X1 port map( A1 => n98694, A2 => n119851, B1 => n99626, B2 =>
                           n119845, ZN => n117560);
   U85906 : OAI22_X1 port map( A1 => n98693, A2 => n119851, B1 => n99625, B2 =>
                           n119845, ZN => n117538);
   U85907 : OAI22_X1 port map( A1 => n98692, A2 => n119851, B1 => n99624, B2 =>
                           n119845, ZN => n117515);
   U85908 : OAI22_X1 port map( A1 => n98691, A2 => n119851, B1 => n99623, B2 =>
                           n119845, ZN => n117492);
   U85909 : OAI22_X1 port map( A1 => n98690, A2 => n119851, B1 => n99622, B2 =>
                           n119845, ZN => n117469);
   U85910 : OAI22_X1 port map( A1 => n98689, A2 => n119851, B1 => n99621, B2 =>
                           n119845, ZN => n117446);
   U85911 : OAI22_X1 port map( A1 => n98688, A2 => n119852, B1 => n99620, B2 =>
                           n119846, ZN => n117423);
   U85912 : OAI22_X1 port map( A1 => n98687, A2 => n119852, B1 => n99619, B2 =>
                           n119846, ZN => n117400);
   U85913 : OAI22_X1 port map( A1 => n98686, A2 => n119852, B1 => n99618, B2 =>
                           n119846, ZN => n117377);
   U85914 : OAI22_X1 port map( A1 => n98685, A2 => n119852, B1 => n99617, B2 =>
                           n119846, ZN => n117354);
   U85915 : OAI22_X1 port map( A1 => n98684, A2 => n119852, B1 => n99616, B2 =>
                           n119846, ZN => n117331);
   U85916 : OAI22_X1 port map( A1 => n98683, A2 => n119852, B1 => n99615, B2 =>
                           n119846, ZN => n117308);
   U85917 : OAI22_X1 port map( A1 => n98682, A2 => n119852, B1 => n99614, B2 =>
                           n119846, ZN => n117285);
   U85918 : OAI22_X1 port map( A1 => n98681, A2 => n119852, B1 => n99613, B2 =>
                           n119846, ZN => n117262);
   U85919 : OAI22_X1 port map( A1 => n98680, A2 => n119852, B1 => n99612, B2 =>
                           n119846, ZN => n117239);
   U85920 : OAI22_X1 port map( A1 => n98679, A2 => n119852, B1 => n99611, B2 =>
                           n119846, ZN => n117216);
   U85921 : OAI22_X1 port map( A1 => n98678, A2 => n119852, B1 => n99610, B2 =>
                           n119846, ZN => n117193);
   U85922 : OAI22_X1 port map( A1 => n98677, A2 => n119852, B1 => n99609, B2 =>
                           n119846, ZN => n117170);
   U85923 : OAI22_X1 port map( A1 => n98676, A2 => n119853, B1 => n99608, B2 =>
                           n119847, ZN => n117147);
   U85924 : OAI22_X1 port map( A1 => n98675, A2 => n119853, B1 => n99607, B2 =>
                           n119847, ZN => n117124);
   U85925 : OAI22_X1 port map( A1 => n98674, A2 => n119853, B1 => n99606, B2 =>
                           n119847, ZN => n117101);
   U85926 : OAI22_X1 port map( A1 => n98673, A2 => n119853, B1 => n99605, B2 =>
                           n119847, ZN => n117078);
   U85927 : OAI22_X1 port map( A1 => n98672, A2 => n119853, B1 => n99604, B2 =>
                           n119847, ZN => n117055);
   U85928 : OAI22_X1 port map( A1 => n98671, A2 => n119853, B1 => n99603, B2 =>
                           n119847, ZN => n117032);
   U85929 : OAI22_X1 port map( A1 => n98670, A2 => n119853, B1 => n99602, B2 =>
                           n119847, ZN => n117009);
   U85930 : OAI22_X1 port map( A1 => n98669, A2 => n119853, B1 => n99601, B2 =>
                           n119847, ZN => n116986);
   U85931 : OAI22_X1 port map( A1 => n98668, A2 => n119853, B1 => n99600, B2 =>
                           n119847, ZN => n116963);
   U85932 : OAI22_X1 port map( A1 => n98667, A2 => n119853, B1 => n99599, B2 =>
                           n119847, ZN => n116940);
   U85933 : OAI22_X1 port map( A1 => n98666, A2 => n119853, B1 => n99598, B2 =>
                           n119847, ZN => n116917);
   U85934 : OAI22_X1 port map( A1 => n98665, A2 => n119853, B1 => n99597, B2 =>
                           n119847, ZN => n116894);
   U85935 : OAI22_X1 port map( A1 => n98664, A2 => n119854, B1 => n99596, B2 =>
                           n119848, ZN => n116871);
   U85936 : OAI22_X1 port map( A1 => n98663, A2 => n119854, B1 => n99595, B2 =>
                           n119848, ZN => n116848);
   U85937 : OAI22_X1 port map( A1 => n98662, A2 => n119854, B1 => n99594, B2 =>
                           n119848, ZN => n116825);
   U85938 : OAI22_X1 port map( A1 => n98661, A2 => n119854, B1 => n99593, B2 =>
                           n119848, ZN => n116802);
   U85939 : OAI22_X1 port map( A1 => n98660, A2 => n119854, B1 => n99592, B2 =>
                           n119848, ZN => n116779);
   U85940 : OAI22_X1 port map( A1 => n98659, A2 => n119854, B1 => n99591, B2 =>
                           n119848, ZN => n116756);
   U85941 : OAI22_X1 port map( A1 => n98658, A2 => n119854, B1 => n99590, B2 =>
                           n119848, ZN => n116733);
   U85942 : OAI22_X1 port map( A1 => n98657, A2 => n119854, B1 => n99589, B2 =>
                           n119848, ZN => n116710);
   U85943 : OAI22_X1 port map( A1 => n98656, A2 => n119854, B1 => n99588, B2 =>
                           n119848, ZN => n116687);
   U85944 : OAI22_X1 port map( A1 => n98655, A2 => n119854, B1 => n99587, B2 =>
                           n119848, ZN => n116664);
   U85945 : OAI22_X1 port map( A1 => n98654, A2 => n119854, B1 => n99586, B2 =>
                           n119848, ZN => n116641);
   U85946 : OAI22_X1 port map( A1 => n98653, A2 => n119854, B1 => n99585, B2 =>
                           n119848, ZN => n116618);
   U85947 : OAI22_X1 port map( A1 => n98732, A2 => n120075, B1 => n99932, B2 =>
                           n120069, ZN => n115171);
   U85948 : OAI22_X1 port map( A1 => n98731, A2 => n120075, B1 => n99931, B2 =>
                           n120069, ZN => n115143);
   U85949 : OAI22_X1 port map( A1 => n98730, A2 => n120076, B1 => n99930, B2 =>
                           n120070, ZN => n115115);
   U85950 : OAI22_X1 port map( A1 => n98729, A2 => n120076, B1 => n99929, B2 =>
                           n120070, ZN => n115087);
   U85951 : OAI22_X1 port map( A1 => n98728, A2 => n120076, B1 => n99928, B2 =>
                           n120070, ZN => n115059);
   U85952 : OAI22_X1 port map( A1 => n98727, A2 => n120076, B1 => n99927, B2 =>
                           n120070, ZN => n115031);
   U85953 : OAI22_X1 port map( A1 => n98726, A2 => n120076, B1 => n99926, B2 =>
                           n120070, ZN => n115003);
   U85954 : OAI22_X1 port map( A1 => n98725, A2 => n120076, B1 => n99925, B2 =>
                           n120070, ZN => n114975);
   U85955 : OAI22_X1 port map( A1 => n98724, A2 => n120076, B1 => n99924, B2 =>
                           n120070, ZN => n114947);
   U85956 : OAI22_X1 port map( A1 => n98723, A2 => n120076, B1 => n99923, B2 =>
                           n120070, ZN => n114919);
   U85957 : OAI22_X1 port map( A1 => n98722, A2 => n120076, B1 => n99922, B2 =>
                           n120070, ZN => n114891);
   U85958 : OAI22_X1 port map( A1 => n98721, A2 => n120076, B1 => n99921, B2 =>
                           n120070, ZN => n114863);
   U85959 : OAI22_X1 port map( A1 => n98720, A2 => n120076, B1 => n99920, B2 =>
                           n120070, ZN => n114835);
   U85960 : OAI22_X1 port map( A1 => n98719, A2 => n120076, B1 => n99919, B2 =>
                           n120070, ZN => n114807);
   U85961 : OAI22_X1 port map( A1 => n98778, A2 => n120072, B1 => n99978, B2 =>
                           n120066, ZN => n116474);
   U85962 : OAI22_X1 port map( A1 => n98777, A2 => n120072, B1 => n99977, B2 =>
                           n120066, ZN => n116431);
   U85963 : OAI22_X1 port map( A1 => n98776, A2 => n120072, B1 => n99976, B2 =>
                           n120066, ZN => n116403);
   U85964 : OAI22_X1 port map( A1 => n98775, A2 => n120072, B1 => n99975, B2 =>
                           n120066, ZN => n116375);
   U85965 : OAI22_X1 port map( A1 => n98705, A2 => n119850, B1 => n99637, B2 =>
                           n119844, ZN => n117802);
   U85966 : OAI22_X1 port map( A1 => n98704, A2 => n119850, B1 => n99636, B2 =>
                           n119844, ZN => n117780);
   U85967 : OAI22_X1 port map( A1 => n98703, A2 => n119850, B1 => n99635, B2 =>
                           n119844, ZN => n117758);
   U85968 : OAI22_X1 port map( A1 => n98702, A2 => n119850, B1 => n99634, B2 =>
                           n119844, ZN => n117736);
   U85969 : OAI22_X1 port map( A1 => n98712, A2 => n119850, B1 => n99644, B2 =>
                           n119844, ZN => n117972);
   U85970 : OAI22_X1 port map( A1 => n98711, A2 => n119850, B1 => n99643, B2 =>
                           n119844, ZN => n117934);
   U85971 : OAI22_X1 port map( A1 => n98710, A2 => n119850, B1 => n99642, B2 =>
                           n119844, ZN => n117912);
   U85972 : OAI22_X1 port map( A1 => n98709, A2 => n119850, B1 => n99641, B2 =>
                           n119844, ZN => n117890);
   U85973 : OAI22_X1 port map( A1 => n98708, A2 => n119850, B1 => n99640, B2 =>
                           n119844, ZN => n117868);
   U85974 : OAI22_X1 port map( A1 => n98707, A2 => n119850, B1 => n99639, B2 =>
                           n119844, ZN => n117846);
   U85975 : OAI22_X1 port map( A1 => n98706, A2 => n119850, B1 => n99638, B2 =>
                           n119844, ZN => n117824);
   U85976 : OAI22_X1 port map( A1 => n98774, A2 => n120072, B1 => n99974, B2 =>
                           n120066, ZN => n116347);
   U85977 : OAI22_X1 port map( A1 => n98773, A2 => n120072, B1 => n99973, B2 =>
                           n120066, ZN => n116319);
   U85978 : OAI22_X1 port map( A1 => n98772, A2 => n120072, B1 => n99972, B2 =>
                           n120066, ZN => n116291);
   U85979 : OAI22_X1 port map( A1 => n98771, A2 => n120072, B1 => n99971, B2 =>
                           n120066, ZN => n116263);
   U85980 : OAI22_X1 port map( A1 => n98770, A2 => n120072, B1 => n99970, B2 =>
                           n120066, ZN => n116235);
   U85981 : OAI22_X1 port map( A1 => n98769, A2 => n120072, B1 => n99969, B2 =>
                           n120066, ZN => n116207);
   U85982 : OAI22_X1 port map( A1 => n98768, A2 => n120072, B1 => n99968, B2 =>
                           n120066, ZN => n116179);
   U85983 : OAI22_X1 port map( A1 => n98767, A2 => n120072, B1 => n99967, B2 =>
                           n120066, ZN => n116151);
   U85984 : OAI22_X1 port map( A1 => n98766, A2 => n120073, B1 => n99966, B2 =>
                           n120067, ZN => n116123);
   U85985 : OAI22_X1 port map( A1 => n98765, A2 => n120073, B1 => n99965, B2 =>
                           n120067, ZN => n116095);
   U85986 : OAI22_X1 port map( A1 => n98764, A2 => n120073, B1 => n99964, B2 =>
                           n120067, ZN => n116067);
   U85987 : OAI22_X1 port map( A1 => n98763, A2 => n120073, B1 => n99963, B2 =>
                           n120067, ZN => n116039);
   U85988 : OAI22_X1 port map( A1 => n98762, A2 => n120073, B1 => n99962, B2 =>
                           n120067, ZN => n116011);
   U85989 : OAI22_X1 port map( A1 => n98761, A2 => n120073, B1 => n99961, B2 =>
                           n120067, ZN => n115983);
   U85990 : OAI22_X1 port map( A1 => n98760, A2 => n120073, B1 => n99960, B2 =>
                           n120067, ZN => n115955);
   U85991 : OAI22_X1 port map( A1 => n98759, A2 => n120073, B1 => n99959, B2 =>
                           n120067, ZN => n115927);
   U85992 : OAI22_X1 port map( A1 => n98758, A2 => n120073, B1 => n99958, B2 =>
                           n120067, ZN => n115899);
   U85993 : OAI22_X1 port map( A1 => n98757, A2 => n120073, B1 => n99957, B2 =>
                           n120067, ZN => n115871);
   U85994 : OAI22_X1 port map( A1 => n98756, A2 => n120073, B1 => n99956, B2 =>
                           n120067, ZN => n115843);
   U85995 : OAI22_X1 port map( A1 => n98755, A2 => n120073, B1 => n99955, B2 =>
                           n120067, ZN => n115815);
   U85996 : OAI22_X1 port map( A1 => n98754, A2 => n120074, B1 => n99954, B2 =>
                           n120068, ZN => n115787);
   U85997 : OAI22_X1 port map( A1 => n98753, A2 => n120074, B1 => n99953, B2 =>
                           n120068, ZN => n115759);
   U85998 : OAI22_X1 port map( A1 => n98752, A2 => n120074, B1 => n99952, B2 =>
                           n120068, ZN => n115731);
   U85999 : OAI22_X1 port map( A1 => n98751, A2 => n120074, B1 => n99951, B2 =>
                           n120068, ZN => n115703);
   U86000 : OAI22_X1 port map( A1 => n98750, A2 => n120074, B1 => n99950, B2 =>
                           n120068, ZN => n115675);
   U86001 : OAI22_X1 port map( A1 => n98749, A2 => n120074, B1 => n99949, B2 =>
                           n120068, ZN => n115647);
   U86002 : OAI22_X1 port map( A1 => n98748, A2 => n120074, B1 => n99948, B2 =>
                           n120068, ZN => n115619);
   U86003 : OAI22_X1 port map( A1 => n98747, A2 => n120074, B1 => n99947, B2 =>
                           n120068, ZN => n115591);
   U86004 : OAI22_X1 port map( A1 => n98746, A2 => n120074, B1 => n99946, B2 =>
                           n120068, ZN => n115563);
   U86005 : OAI22_X1 port map( A1 => n98745, A2 => n120074, B1 => n99945, B2 =>
                           n120068, ZN => n115535);
   U86006 : OAI22_X1 port map( A1 => n98744, A2 => n120074, B1 => n99944, B2 =>
                           n120068, ZN => n115507);
   U86007 : OAI22_X1 port map( A1 => n98743, A2 => n120074, B1 => n99943, B2 =>
                           n120068, ZN => n115479);
   U86008 : OAI22_X1 port map( A1 => n98742, A2 => n120075, B1 => n99942, B2 =>
                           n120069, ZN => n115451);
   U86009 : OAI22_X1 port map( A1 => n98741, A2 => n120075, B1 => n99941, B2 =>
                           n120069, ZN => n115423);
   U86010 : OAI22_X1 port map( A1 => n98740, A2 => n120075, B1 => n99940, B2 =>
                           n120069, ZN => n115395);
   U86011 : OAI22_X1 port map( A1 => n98739, A2 => n120075, B1 => n99939, B2 =>
                           n120069, ZN => n115367);
   U86012 : OAI22_X1 port map( A1 => n98738, A2 => n120075, B1 => n99938, B2 =>
                           n120069, ZN => n115339);
   U86013 : OAI22_X1 port map( A1 => n98737, A2 => n120075, B1 => n99937, B2 =>
                           n120069, ZN => n115311);
   U86014 : OAI22_X1 port map( A1 => n98736, A2 => n120075, B1 => n99936, B2 =>
                           n120069, ZN => n115283);
   U86015 : OAI22_X1 port map( A1 => n98735, A2 => n120075, B1 => n99935, B2 =>
                           n120069, ZN => n115255);
   U86016 : OAI22_X1 port map( A1 => n98734, A2 => n120075, B1 => n99934, B2 =>
                           n120069, ZN => n115227);
   U86017 : OAI22_X1 port map( A1 => n98733, A2 => n120075, B1 => n99933, B2 =>
                           n120069, ZN => n115199);
   U86018 : OAI22_X1 port map( A1 => n114040, A2 => n119874, B1 => n99499, B2 
                           => n119868, ZN => n117713);
   U86019 : OAI22_X1 port map( A1 => n114039, A2 => n119875, B1 => n99498, B2 
                           => n119869, ZN => n117691);
   U86020 : OAI22_X1 port map( A1 => n114038, A2 => n119875, B1 => n99497, B2 
                           => n119869, ZN => n117669);
   U86021 : OAI22_X1 port map( A1 => n114037, A2 => n119875, B1 => n99496, B2 
                           => n119869, ZN => n117647);
   U86022 : OAI22_X1 port map( A1 => n114036, A2 => n119875, B1 => n99495, B2 
                           => n119869, ZN => n117625);
   U86023 : OAI22_X1 port map( A1 => n114035, A2 => n119875, B1 => n99494, B2 
                           => n119869, ZN => n117603);
   U86024 : OAI22_X1 port map( A1 => n114034, A2 => n119875, B1 => n99493, B2 
                           => n119869, ZN => n117581);
   U86025 : OAI22_X1 port map( A1 => n114033, A2 => n119875, B1 => n99492, B2 
                           => n119869, ZN => n117559);
   U86026 : OAI22_X1 port map( A1 => n114032, A2 => n119875, B1 => n99491, B2 
                           => n119869, ZN => n117537);
   U86027 : OAI22_X1 port map( A1 => n114031, A2 => n119875, B1 => n99490, B2 
                           => n119869, ZN => n117514);
   U86028 : OAI22_X1 port map( A1 => n114030, A2 => n119875, B1 => n99489, B2 
                           => n119869, ZN => n117491);
   U86029 : OAI22_X1 port map( A1 => n114029, A2 => n119875, B1 => n99488, B2 
                           => n119869, ZN => n117468);
   U86030 : OAI22_X1 port map( A1 => n114028, A2 => n119875, B1 => n99487, B2 
                           => n119869, ZN => n117445);
   U86031 : OAI22_X1 port map( A1 => n114027, A2 => n119876, B1 => n99486, B2 
                           => n119870, ZN => n117422);
   U86032 : OAI22_X1 port map( A1 => n114026, A2 => n119876, B1 => n99485, B2 
                           => n119870, ZN => n117399);
   U86033 : OAI22_X1 port map( A1 => n114025, A2 => n119876, B1 => n99484, B2 
                           => n119870, ZN => n117376);
   U86034 : OAI22_X1 port map( A1 => n114024, A2 => n119876, B1 => n99483, B2 
                           => n119870, ZN => n117353);
   U86035 : OAI22_X1 port map( A1 => n114023, A2 => n119876, B1 => n99482, B2 
                           => n119870, ZN => n117330);
   U86036 : OAI22_X1 port map( A1 => n114022, A2 => n119876, B1 => n99481, B2 
                           => n119870, ZN => n117307);
   U86037 : OAI22_X1 port map( A1 => n114021, A2 => n119876, B1 => n99480, B2 
                           => n119870, ZN => n117284);
   U86038 : OAI22_X1 port map( A1 => n114020, A2 => n119876, B1 => n99479, B2 
                           => n119870, ZN => n117261);
   U86039 : OAI22_X1 port map( A1 => n114019, A2 => n119876, B1 => n99478, B2 
                           => n119870, ZN => n117238);
   U86040 : OAI22_X1 port map( A1 => n114018, A2 => n119876, B1 => n99477, B2 
                           => n119870, ZN => n117215);
   U86041 : OAI22_X1 port map( A1 => n114017, A2 => n119876, B1 => n99476, B2 
                           => n119870, ZN => n117192);
   U86042 : OAI22_X1 port map( A1 => n114016, A2 => n119876, B1 => n99475, B2 
                           => n119870, ZN => n117169);
   U86043 : OAI22_X1 port map( A1 => n114015, A2 => n119877, B1 => n99474, B2 
                           => n119871, ZN => n117146);
   U86044 : OAI22_X1 port map( A1 => n114014, A2 => n119877, B1 => n99473, B2 
                           => n119871, ZN => n117123);
   U86045 : OAI22_X1 port map( A1 => n114013, A2 => n119877, B1 => n99472, B2 
                           => n119871, ZN => n117100);
   U86046 : OAI22_X1 port map( A1 => n114012, A2 => n119877, B1 => n99471, B2 
                           => n119871, ZN => n117077);
   U86047 : OAI22_X1 port map( A1 => n114011, A2 => n119877, B1 => n99470, B2 
                           => n119871, ZN => n117054);
   U86048 : OAI22_X1 port map( A1 => n114010, A2 => n119877, B1 => n99469, B2 
                           => n119871, ZN => n117031);
   U86049 : OAI22_X1 port map( A1 => n114009, A2 => n119877, B1 => n99468, B2 
                           => n119871, ZN => n117008);
   U86050 : OAI22_X1 port map( A1 => n114008, A2 => n119877, B1 => n99467, B2 
                           => n119871, ZN => n116985);
   U86051 : OAI22_X1 port map( A1 => n114007, A2 => n119877, B1 => n99466, B2 
                           => n119871, ZN => n116962);
   U86052 : OAI22_X1 port map( A1 => n114006, A2 => n119877, B1 => n99465, B2 
                           => n119871, ZN => n116939);
   U86053 : OAI22_X1 port map( A1 => n114005, A2 => n119877, B1 => n99464, B2 
                           => n119871, ZN => n116916);
   U86054 : OAI22_X1 port map( A1 => n114004, A2 => n119877, B1 => n99463, B2 
                           => n119871, ZN => n116893);
   U86055 : OAI22_X1 port map( A1 => n114003, A2 => n119878, B1 => n99462, B2 
                           => n119872, ZN => n116870);
   U86056 : OAI22_X1 port map( A1 => n114002, A2 => n119878, B1 => n99461, B2 
                           => n119872, ZN => n116847);
   U86057 : OAI22_X1 port map( A1 => n114001, A2 => n119878, B1 => n99460, B2 
                           => n119872, ZN => n116824);
   U86058 : OAI22_X1 port map( A1 => n114000, A2 => n119878, B1 => n99459, B2 
                           => n119872, ZN => n116801);
   U86059 : OAI22_X1 port map( A1 => n113999, A2 => n119878, B1 => n99458, B2 
                           => n119872, ZN => n116778);
   U86060 : OAI22_X1 port map( A1 => n113998, A2 => n119878, B1 => n99457, B2 
                           => n119872, ZN => n116755);
   U86061 : OAI22_X1 port map( A1 => n113997, A2 => n119878, B1 => n99456, B2 
                           => n119872, ZN => n116732);
   U86062 : OAI22_X1 port map( A1 => n113996, A2 => n119878, B1 => n99455, B2 
                           => n119872, ZN => n116709);
   U86063 : OAI22_X1 port map( A1 => n113995, A2 => n119878, B1 => n99454, B2 
                           => n119872, ZN => n116686);
   U86064 : OAI22_X1 port map( A1 => n113994, A2 => n119878, B1 => n99453, B2 
                           => n119872, ZN => n116663);
   U86065 : OAI22_X1 port map( A1 => n113993, A2 => n119878, B1 => n99452, B2 
                           => n119872, ZN => n116640);
   U86066 : OAI22_X1 port map( A1 => n113992, A2 => n119878, B1 => n99451, B2 
                           => n119872, ZN => n116617);
   U86067 : OAI22_X1 port map( A1 => n114044, A2 => n119874, B1 => n99503, B2 
                           => n119868, ZN => n117801);
   U86068 : OAI22_X1 port map( A1 => n114043, A2 => n119874, B1 => n99502, B2 
                           => n119868, ZN => n117779);
   U86069 : OAI22_X1 port map( A1 => n114042, A2 => n119874, B1 => n99501, B2 
                           => n119868, ZN => n117757);
   U86070 : OAI22_X1 port map( A1 => n114041, A2 => n119874, B1 => n99500, B2 
                           => n119868, ZN => n117735);
   U86071 : OAI22_X1 port map( A1 => n114051, A2 => n119874, B1 => n99510, B2 
                           => n119868, ZN => n117969);
   U86072 : OAI22_X1 port map( A1 => n114050, A2 => n119874, B1 => n99509, B2 
                           => n119868, ZN => n117933);
   U86073 : OAI22_X1 port map( A1 => n114049, A2 => n119874, B1 => n99508, B2 
                           => n119868, ZN => n117911);
   U86074 : OAI22_X1 port map( A1 => n114048, A2 => n119874, B1 => n99507, B2 
                           => n119868, ZN => n117889);
   U86075 : OAI22_X1 port map( A1 => n114047, A2 => n119874, B1 => n99506, B2 
                           => n119868, ZN => n117867);
   U86076 : OAI22_X1 port map( A1 => n114046, A2 => n119874, B1 => n99505, B2 
                           => n119868, ZN => n117845);
   U86077 : OAI22_X1 port map( A1 => n114045, A2 => n119874, B1 => n99504, B2 
                           => n119868, ZN => n117823);
   U86078 : OAI22_X1 port map( A1 => n99769, A2 => n119940, B1 => n113868, B2 
                           => n119934, ZN => n117712);
   U86079 : OAI22_X1 port map( A1 => n99768, A2 => n119941, B1 => n113866, B2 
                           => n119935, ZN => n117690);
   U86080 : OAI22_X1 port map( A1 => n99767, A2 => n119941, B1 => n113864, B2 
                           => n119935, ZN => n117668);
   U86081 : OAI22_X1 port map( A1 => n99766, A2 => n119941, B1 => n113862, B2 
                           => n119935, ZN => n117646);
   U86082 : OAI22_X1 port map( A1 => n99765, A2 => n119941, B1 => n113860, B2 
                           => n119935, ZN => n117624);
   U86083 : OAI22_X1 port map( A1 => n99764, A2 => n119941, B1 => n113858, B2 
                           => n119935, ZN => n117602);
   U86084 : OAI22_X1 port map( A1 => n99763, A2 => n119941, B1 => n113856, B2 
                           => n119935, ZN => n117580);
   U86085 : OAI22_X1 port map( A1 => n99762, A2 => n119941, B1 => n113854, B2 
                           => n119935, ZN => n117558);
   U86086 : OAI22_X1 port map( A1 => n99761, A2 => n119941, B1 => n113852, B2 
                           => n119935, ZN => n117535);
   U86087 : OAI22_X1 port map( A1 => n99760, A2 => n119941, B1 => n113850, B2 
                           => n119935, ZN => n117512);
   U86088 : OAI22_X1 port map( A1 => n99759, A2 => n119941, B1 => n113848, B2 
                           => n119935, ZN => n117489);
   U86089 : OAI22_X1 port map( A1 => n99758, A2 => n119941, B1 => n113846, B2 
                           => n119935, ZN => n117466);
   U86090 : OAI22_X1 port map( A1 => n99757, A2 => n119941, B1 => n113844, B2 
                           => n119935, ZN => n117443);
   U86091 : OAI22_X1 port map( A1 => n99756, A2 => n119942, B1 => n113842, B2 
                           => n119936, ZN => n117420);
   U86092 : OAI22_X1 port map( A1 => n99755, A2 => n119942, B1 => n113840, B2 
                           => n119936, ZN => n117397);
   U86093 : OAI22_X1 port map( A1 => n99754, A2 => n119942, B1 => n113838, B2 
                           => n119936, ZN => n117374);
   U86094 : OAI22_X1 port map( A1 => n99753, A2 => n119942, B1 => n113836, B2 
                           => n119936, ZN => n117351);
   U86095 : OAI22_X1 port map( A1 => n99752, A2 => n119942, B1 => n113834, B2 
                           => n119936, ZN => n117328);
   U86096 : OAI22_X1 port map( A1 => n99751, A2 => n119942, B1 => n113832, B2 
                           => n119936, ZN => n117305);
   U86097 : OAI22_X1 port map( A1 => n99750, A2 => n119942, B1 => n113830, B2 
                           => n119936, ZN => n117282);
   U86098 : OAI22_X1 port map( A1 => n99749, A2 => n119942, B1 => n113828, B2 
                           => n119936, ZN => n117259);
   U86099 : OAI22_X1 port map( A1 => n99748, A2 => n119942, B1 => n113826, B2 
                           => n119936, ZN => n117236);
   U86100 : OAI22_X1 port map( A1 => n99747, A2 => n119942, B1 => n113824, B2 
                           => n119936, ZN => n117213);
   U86101 : OAI22_X1 port map( A1 => n99746, A2 => n119942, B1 => n113822, B2 
                           => n119936, ZN => n117190);
   U86102 : OAI22_X1 port map( A1 => n99745, A2 => n119942, B1 => n113820, B2 
                           => n119936, ZN => n117167);
   U86103 : OAI22_X1 port map( A1 => n99744, A2 => n119943, B1 => n113818, B2 
                           => n119937, ZN => n117144);
   U86104 : OAI22_X1 port map( A1 => n99743, A2 => n119943, B1 => n113816, B2 
                           => n119937, ZN => n117121);
   U86105 : OAI22_X1 port map( A1 => n99742, A2 => n119943, B1 => n113814, B2 
                           => n119937, ZN => n117098);
   U86106 : OAI22_X1 port map( A1 => n99741, A2 => n119943, B1 => n113812, B2 
                           => n119937, ZN => n117075);
   U86107 : OAI22_X1 port map( A1 => n99740, A2 => n119943, B1 => n113810, B2 
                           => n119937, ZN => n117052);
   U86108 : OAI22_X1 port map( A1 => n99739, A2 => n119943, B1 => n113808, B2 
                           => n119937, ZN => n117029);
   U86109 : OAI22_X1 port map( A1 => n99738, A2 => n119943, B1 => n113806, B2 
                           => n119937, ZN => n117006);
   U86110 : OAI22_X1 port map( A1 => n99737, A2 => n119943, B1 => n113804, B2 
                           => n119937, ZN => n116983);
   U86111 : OAI22_X1 port map( A1 => n99736, A2 => n119943, B1 => n113802, B2 
                           => n119937, ZN => n116960);
   U86112 : OAI22_X1 port map( A1 => n99735, A2 => n119943, B1 => n113800, B2 
                           => n119937, ZN => n116937);
   U86113 : OAI22_X1 port map( A1 => n99734, A2 => n119943, B1 => n113798, B2 
                           => n119937, ZN => n116914);
   U86114 : OAI22_X1 port map( A1 => n99733, A2 => n119943, B1 => n113796, B2 
                           => n119937, ZN => n116891);
   U86115 : OAI22_X1 port map( A1 => n99732, A2 => n119944, B1 => n113794, B2 
                           => n119938, ZN => n116868);
   U86116 : OAI22_X1 port map( A1 => n99731, A2 => n119944, B1 => n113792, B2 
                           => n119938, ZN => n116845);
   U86117 : OAI22_X1 port map( A1 => n99730, A2 => n119944, B1 => n113790, B2 
                           => n119938, ZN => n116822);
   U86118 : OAI22_X1 port map( A1 => n99729, A2 => n119944, B1 => n113788, B2 
                           => n119938, ZN => n116799);
   U86119 : OAI22_X1 port map( A1 => n99728, A2 => n119944, B1 => n113786, B2 
                           => n119938, ZN => n116776);
   U86120 : OAI22_X1 port map( A1 => n99727, A2 => n119944, B1 => n113784, B2 
                           => n119938, ZN => n116753);
   U86121 : OAI22_X1 port map( A1 => n99726, A2 => n119944, B1 => n113782, B2 
                           => n119938, ZN => n116730);
   U86122 : OAI22_X1 port map( A1 => n99725, A2 => n119944, B1 => n113780, B2 
                           => n119938, ZN => n116707);
   U86123 : OAI22_X1 port map( A1 => n99724, A2 => n119944, B1 => n113778, B2 
                           => n119938, ZN => n116684);
   U86124 : OAI22_X1 port map( A1 => n99723, A2 => n119944, B1 => n113776, B2 
                           => n119938, ZN => n116661);
   U86125 : OAI22_X1 port map( A1 => n99722, A2 => n119944, B1 => n113774, B2 
                           => n119938, ZN => n116638);
   U86126 : OAI22_X1 port map( A1 => n99721, A2 => n119944, B1 => n113772, B2 
                           => n119938, ZN => n116615);
   U86127 : OAI22_X1 port map( A1 => n99065, A2 => n120141, B1 => n113798, B2 
                           => n120135, ZN => n115168);
   U86128 : OAI22_X1 port map( A1 => n99064, A2 => n120141, B1 => n113796, B2 
                           => n120135, ZN => n115140);
   U86129 : OAI22_X1 port map( A1 => n99063, A2 => n120142, B1 => n113794, B2 
                           => n120136, ZN => n115112);
   U86130 : OAI22_X1 port map( A1 => n99062, A2 => n120142, B1 => n113792, B2 
                           => n120136, ZN => n115084);
   U86131 : OAI22_X1 port map( A1 => n99061, A2 => n120142, B1 => n113790, B2 
                           => n120136, ZN => n115056);
   U86132 : OAI22_X1 port map( A1 => n99060, A2 => n120142, B1 => n113788, B2 
                           => n120136, ZN => n115028);
   U86133 : OAI22_X1 port map( A1 => n99059, A2 => n120142, B1 => n113786, B2 
                           => n120136, ZN => n115000);
   U86134 : OAI22_X1 port map( A1 => n99058, A2 => n120142, B1 => n113784, B2 
                           => n120136, ZN => n114972);
   U86135 : OAI22_X1 port map( A1 => n99057, A2 => n120142, B1 => n113782, B2 
                           => n120136, ZN => n114944);
   U86136 : OAI22_X1 port map( A1 => n99056, A2 => n120142, B1 => n113780, B2 
                           => n120136, ZN => n114916);
   U86137 : OAI22_X1 port map( A1 => n99055, A2 => n120142, B1 => n113778, B2 
                           => n120136, ZN => n114888);
   U86138 : OAI22_X1 port map( A1 => n99054, A2 => n120142, B1 => n113776, B2 
                           => n120136, ZN => n114860);
   U86139 : OAI22_X1 port map( A1 => n99053, A2 => n120142, B1 => n113774, B2 
                           => n120136, ZN => n114832);
   U86140 : OAI22_X1 port map( A1 => n99052, A2 => n120142, B1 => n113772, B2 
                           => n120136, ZN => n114804);
   U86141 : OAI22_X1 port map( A1 => n99111, A2 => n120138, B1 => n113890, B2 
                           => n120132, ZN => n116468);
   U86142 : OAI22_X1 port map( A1 => n99110, A2 => n120138, B1 => n113888, B2 
                           => n120132, ZN => n116428);
   U86143 : OAI22_X1 port map( A1 => n99109, A2 => n120138, B1 => n113886, B2 
                           => n120132, ZN => n116400);
   U86144 : OAI22_X1 port map( A1 => n99108, A2 => n120138, B1 => n113884, B2 
                           => n120132, ZN => n116372);
   U86145 : OAI22_X1 port map( A1 => n99773, A2 => n119940, B1 => n113876, B2 
                           => n119934, ZN => n117800);
   U86146 : OAI22_X1 port map( A1 => n99772, A2 => n119940, B1 => n113874, B2 
                           => n119934, ZN => n117778);
   U86147 : OAI22_X1 port map( A1 => n99771, A2 => n119940, B1 => n113872, B2 
                           => n119934, ZN => n117756);
   U86148 : OAI22_X1 port map( A1 => n99770, A2 => n119940, B1 => n113870, B2 
                           => n119934, ZN => n117734);
   U86149 : OAI22_X1 port map( A1 => n99780, A2 => n119940, B1 => n113890, B2 
                           => n119934, ZN => n117966);
   U86150 : OAI22_X1 port map( A1 => n99779, A2 => n119940, B1 => n113888, B2 
                           => n119934, ZN => n117932);
   U86151 : OAI22_X1 port map( A1 => n99778, A2 => n119940, B1 => n113886, B2 
                           => n119934, ZN => n117910);
   U86152 : OAI22_X1 port map( A1 => n99777, A2 => n119940, B1 => n113884, B2 
                           => n119934, ZN => n117888);
   U86153 : OAI22_X1 port map( A1 => n99776, A2 => n119940, B1 => n113882, B2 
                           => n119934, ZN => n117866);
   U86154 : OAI22_X1 port map( A1 => n99775, A2 => n119940, B1 => n113880, B2 
                           => n119934, ZN => n117844);
   U86155 : OAI22_X1 port map( A1 => n99774, A2 => n119940, B1 => n113878, B2 
                           => n119934, ZN => n117822);
   U86156 : OAI22_X1 port map( A1 => n99107, A2 => n120138, B1 => n113882, B2 
                           => n120132, ZN => n116344);
   U86157 : OAI22_X1 port map( A1 => n99106, A2 => n120138, B1 => n113880, B2 
                           => n120132, ZN => n116316);
   U86158 : OAI22_X1 port map( A1 => n99105, A2 => n120138, B1 => n113878, B2 
                           => n120132, ZN => n116288);
   U86159 : OAI22_X1 port map( A1 => n99104, A2 => n120138, B1 => n113876, B2 
                           => n120132, ZN => n116260);
   U86160 : OAI22_X1 port map( A1 => n99103, A2 => n120138, B1 => n113874, B2 
                           => n120132, ZN => n116232);
   U86161 : OAI22_X1 port map( A1 => n99102, A2 => n120138, B1 => n113872, B2 
                           => n120132, ZN => n116204);
   U86162 : OAI22_X1 port map( A1 => n99101, A2 => n120138, B1 => n113870, B2 
                           => n120132, ZN => n116176);
   U86163 : OAI22_X1 port map( A1 => n99100, A2 => n120138, B1 => n113868, B2 
                           => n120132, ZN => n116148);
   U86164 : OAI22_X1 port map( A1 => n99099, A2 => n120139, B1 => n113866, B2 
                           => n120133, ZN => n116120);
   U86165 : OAI22_X1 port map( A1 => n99098, A2 => n120139, B1 => n113864, B2 
                           => n120133, ZN => n116092);
   U86166 : OAI22_X1 port map( A1 => n99097, A2 => n120139, B1 => n113862, B2 
                           => n120133, ZN => n116064);
   U86167 : OAI22_X1 port map( A1 => n99096, A2 => n120139, B1 => n113860, B2 
                           => n120133, ZN => n116036);
   U86168 : OAI22_X1 port map( A1 => n99095, A2 => n120139, B1 => n113858, B2 
                           => n120133, ZN => n116008);
   U86169 : OAI22_X1 port map( A1 => n99094, A2 => n120139, B1 => n113856, B2 
                           => n120133, ZN => n115980);
   U86170 : OAI22_X1 port map( A1 => n99093, A2 => n120139, B1 => n113854, B2 
                           => n120133, ZN => n115952);
   U86171 : OAI22_X1 port map( A1 => n99092, A2 => n120139, B1 => n113852, B2 
                           => n120133, ZN => n115924);
   U86172 : OAI22_X1 port map( A1 => n99091, A2 => n120139, B1 => n113850, B2 
                           => n120133, ZN => n115896);
   U86173 : OAI22_X1 port map( A1 => n99090, A2 => n120139, B1 => n113848, B2 
                           => n120133, ZN => n115868);
   U86174 : OAI22_X1 port map( A1 => n99089, A2 => n120139, B1 => n113846, B2 
                           => n120133, ZN => n115840);
   U86175 : OAI22_X1 port map( A1 => n99088, A2 => n120139, B1 => n113844, B2 
                           => n120133, ZN => n115812);
   U86176 : OAI22_X1 port map( A1 => n99087, A2 => n120140, B1 => n113842, B2 
                           => n120134, ZN => n115784);
   U86177 : OAI22_X1 port map( A1 => n99086, A2 => n120140, B1 => n113840, B2 
                           => n120134, ZN => n115756);
   U86178 : OAI22_X1 port map( A1 => n99085, A2 => n120140, B1 => n113838, B2 
                           => n120134, ZN => n115728);
   U86179 : OAI22_X1 port map( A1 => n99084, A2 => n120140, B1 => n113836, B2 
                           => n120134, ZN => n115700);
   U86180 : OAI22_X1 port map( A1 => n99083, A2 => n120140, B1 => n113834, B2 
                           => n120134, ZN => n115672);
   U86181 : OAI22_X1 port map( A1 => n99082, A2 => n120140, B1 => n113832, B2 
                           => n120134, ZN => n115644);
   U86182 : OAI22_X1 port map( A1 => n99081, A2 => n120140, B1 => n113830, B2 
                           => n120134, ZN => n115616);
   U86183 : OAI22_X1 port map( A1 => n99080, A2 => n120140, B1 => n113828, B2 
                           => n120134, ZN => n115588);
   U86184 : OAI22_X1 port map( A1 => n99079, A2 => n120140, B1 => n113826, B2 
                           => n120134, ZN => n115560);
   U86185 : OAI22_X1 port map( A1 => n99078, A2 => n120140, B1 => n113824, B2 
                           => n120134, ZN => n115532);
   U86186 : OAI22_X1 port map( A1 => n99077, A2 => n120140, B1 => n113822, B2 
                           => n120134, ZN => n115504);
   U86187 : OAI22_X1 port map( A1 => n99076, A2 => n120140, B1 => n113820, B2 
                           => n120134, ZN => n115476);
   U86188 : OAI22_X1 port map( A1 => n99075, A2 => n120141, B1 => n113818, B2 
                           => n120135, ZN => n115448);
   U86189 : OAI22_X1 port map( A1 => n99074, A2 => n120141, B1 => n113816, B2 
                           => n120135, ZN => n115420);
   U86190 : OAI22_X1 port map( A1 => n99073, A2 => n120141, B1 => n113814, B2 
                           => n120135, ZN => n115392);
   U86191 : OAI22_X1 port map( A1 => n99072, A2 => n120141, B1 => n113812, B2 
                           => n120135, ZN => n115364);
   U86192 : OAI22_X1 port map( A1 => n99071, A2 => n120141, B1 => n113810, B2 
                           => n120135, ZN => n115336);
   U86193 : OAI22_X1 port map( A1 => n99070, A2 => n120141, B1 => n113808, B2 
                           => n120135, ZN => n115308);
   U86194 : OAI22_X1 port map( A1 => n99069, A2 => n120141, B1 => n113806, B2 
                           => n120135, ZN => n115280);
   U86195 : OAI22_X1 port map( A1 => n99068, A2 => n120141, B1 => n113804, B2 
                           => n120135, ZN => n115252);
   U86196 : OAI22_X1 port map( A1 => n99067, A2 => n120141, B1 => n113802, B2 
                           => n120135, ZN => n115224);
   U86197 : OAI22_X1 port map( A1 => n99066, A2 => n120141, B1 => n113800, B2 
                           => n120135, ZN => n115196);
   U86198 : OAI22_X1 port map( A1 => n98767, A2 => n119916, B1 => n90426, B2 =>
                           n119910, ZN => n117710);
   U86199 : OAI22_X1 port map( A1 => n98766, A2 => n119917, B1 => n90425, B2 =>
                           n119911, ZN => n117688);
   U86200 : OAI22_X1 port map( A1 => n98765, A2 => n119917, B1 => n90424, B2 =>
                           n119911, ZN => n117666);
   U86201 : OAI22_X1 port map( A1 => n98764, A2 => n119917, B1 => n90423, B2 =>
                           n119911, ZN => n117644);
   U86202 : OAI22_X1 port map( A1 => n98763, A2 => n119917, B1 => n90422, B2 =>
                           n119911, ZN => n117622);
   U86203 : OAI22_X1 port map( A1 => n98762, A2 => n119917, B1 => n90421, B2 =>
                           n119911, ZN => n117600);
   U86204 : OAI22_X1 port map( A1 => n98761, A2 => n119917, B1 => n90420, B2 =>
                           n119911, ZN => n117578);
   U86205 : OAI22_X1 port map( A1 => n98760, A2 => n119917, B1 => n90419, B2 =>
                           n119911, ZN => n117556);
   U86206 : OAI22_X1 port map( A1 => n98759, A2 => n119917, B1 => n90418, B2 =>
                           n119911, ZN => n117533);
   U86207 : OAI22_X1 port map( A1 => n98758, A2 => n119917, B1 => n90417, B2 =>
                           n119911, ZN => n117510);
   U86208 : OAI22_X1 port map( A1 => n98757, A2 => n119917, B1 => n90416, B2 =>
                           n119911, ZN => n117487);
   U86209 : OAI22_X1 port map( A1 => n98756, A2 => n119917, B1 => n90415, B2 =>
                           n119911, ZN => n117464);
   U86210 : OAI22_X1 port map( A1 => n98755, A2 => n119917, B1 => n90414, B2 =>
                           n119911, ZN => n117441);
   U86211 : OAI22_X1 port map( A1 => n98754, A2 => n119918, B1 => n90413, B2 =>
                           n119912, ZN => n117418);
   U86212 : OAI22_X1 port map( A1 => n98753, A2 => n119918, B1 => n90412, B2 =>
                           n119912, ZN => n117395);
   U86213 : OAI22_X1 port map( A1 => n98752, A2 => n119918, B1 => n90411, B2 =>
                           n119912, ZN => n117372);
   U86214 : OAI22_X1 port map( A1 => n98751, A2 => n119918, B1 => n90410, B2 =>
                           n119912, ZN => n117349);
   U86215 : OAI22_X1 port map( A1 => n98750, A2 => n119918, B1 => n90409, B2 =>
                           n119912, ZN => n117326);
   U86216 : OAI22_X1 port map( A1 => n98749, A2 => n119918, B1 => n90408, B2 =>
                           n119912, ZN => n117303);
   U86217 : OAI22_X1 port map( A1 => n98748, A2 => n119918, B1 => n90407, B2 =>
                           n119912, ZN => n117280);
   U86218 : OAI22_X1 port map( A1 => n98747, A2 => n119918, B1 => n90406, B2 =>
                           n119912, ZN => n117257);
   U86219 : OAI22_X1 port map( A1 => n98746, A2 => n119918, B1 => n90405, B2 =>
                           n119912, ZN => n117234);
   U86220 : OAI22_X1 port map( A1 => n98745, A2 => n119918, B1 => n90404, B2 =>
                           n119912, ZN => n117211);
   U86221 : OAI22_X1 port map( A1 => n98744, A2 => n119918, B1 => n90403, B2 =>
                           n119912, ZN => n117188);
   U86222 : OAI22_X1 port map( A1 => n98743, A2 => n119918, B1 => n90402, B2 =>
                           n119912, ZN => n117165);
   U86223 : OAI22_X1 port map( A1 => n98742, A2 => n119919, B1 => n90401, B2 =>
                           n119913, ZN => n117142);
   U86224 : OAI22_X1 port map( A1 => n98741, A2 => n119919, B1 => n90400, B2 =>
                           n119913, ZN => n117119);
   U86225 : OAI22_X1 port map( A1 => n98740, A2 => n119919, B1 => n90399, B2 =>
                           n119913, ZN => n117096);
   U86226 : OAI22_X1 port map( A1 => n98739, A2 => n119919, B1 => n90398, B2 =>
                           n119913, ZN => n117073);
   U86227 : OAI22_X1 port map( A1 => n98738, A2 => n119919, B1 => n90397, B2 =>
                           n119913, ZN => n117050);
   U86228 : OAI22_X1 port map( A1 => n98737, A2 => n119919, B1 => n90396, B2 =>
                           n119913, ZN => n117027);
   U86229 : OAI22_X1 port map( A1 => n98736, A2 => n119919, B1 => n90395, B2 =>
                           n119913, ZN => n117004);
   U86230 : OAI22_X1 port map( A1 => n98735, A2 => n119919, B1 => n90394, B2 =>
                           n119913, ZN => n116981);
   U86231 : OAI22_X1 port map( A1 => n98734, A2 => n119919, B1 => n90393, B2 =>
                           n119913, ZN => n116958);
   U86232 : OAI22_X1 port map( A1 => n98733, A2 => n119919, B1 => n90392, B2 =>
                           n119913, ZN => n116935);
   U86233 : OAI22_X1 port map( A1 => n98732, A2 => n119919, B1 => n90391, B2 =>
                           n119913, ZN => n116912);
   U86234 : OAI22_X1 port map( A1 => n98731, A2 => n119919, B1 => n90390, B2 =>
                           n119913, ZN => n116889);
   U86235 : OAI22_X1 port map( A1 => n98730, A2 => n119920, B1 => n90389, B2 =>
                           n119914, ZN => n116866);
   U86236 : OAI22_X1 port map( A1 => n98729, A2 => n119920, B1 => n90388, B2 =>
                           n119914, ZN => n116843);
   U86237 : OAI22_X1 port map( A1 => n98728, A2 => n119920, B1 => n90387, B2 =>
                           n119914, ZN => n116820);
   U86238 : OAI22_X1 port map( A1 => n98727, A2 => n119920, B1 => n90386, B2 =>
                           n119914, ZN => n116797);
   U86239 : OAI22_X1 port map( A1 => n98726, A2 => n119920, B1 => n90385, B2 =>
                           n119914, ZN => n116774);
   U86240 : OAI22_X1 port map( A1 => n98725, A2 => n119920, B1 => n90384, B2 =>
                           n119914, ZN => n116751);
   U86241 : OAI22_X1 port map( A1 => n98724, A2 => n119920, B1 => n90383, B2 =>
                           n119914, ZN => n116728);
   U86242 : OAI22_X1 port map( A1 => n98723, A2 => n119920, B1 => n90382, B2 =>
                           n119914, ZN => n116705);
   U86243 : OAI22_X1 port map( A1 => n98722, A2 => n119920, B1 => n90381, B2 =>
                           n119914, ZN => n116682);
   U86244 : OAI22_X1 port map( A1 => n98721, A2 => n119920, B1 => n90380, B2 =>
                           n119914, ZN => n116659);
   U86245 : OAI22_X1 port map( A1 => n98720, A2 => n119920, B1 => n90379, B2 =>
                           n119914, ZN => n116636);
   U86246 : OAI22_X1 port map( A1 => n98719, A2 => n119920, B1 => n90378, B2 =>
                           n119914, ZN => n116613);
   U86247 : OAI22_X1 port map( A1 => n90530, A2 => n120117, B1 => n90049, B2 =>
                           n120111, ZN => n115166);
   U86248 : OAI22_X1 port map( A1 => n90529, A2 => n120117, B1 => n90048, B2 =>
                           n120111, ZN => n115138);
   U86249 : OAI22_X1 port map( A1 => n90528, A2 => n120118, B1 => n90047, B2 =>
                           n120112, ZN => n115110);
   U86250 : OAI22_X1 port map( A1 => n90527, A2 => n120118, B1 => n90046, B2 =>
                           n120112, ZN => n115082);
   U86251 : OAI22_X1 port map( A1 => n90526, A2 => n120118, B1 => n90045, B2 =>
                           n120112, ZN => n115054);
   U86252 : OAI22_X1 port map( A1 => n90525, A2 => n120118, B1 => n90044, B2 =>
                           n120112, ZN => n115026);
   U86253 : OAI22_X1 port map( A1 => n90524, A2 => n120118, B1 => n90043, B2 =>
                           n120112, ZN => n114998);
   U86254 : OAI22_X1 port map( A1 => n90523, A2 => n120118, B1 => n90042, B2 =>
                           n120112, ZN => n114970);
   U86255 : OAI22_X1 port map( A1 => n90522, A2 => n120118, B1 => n90041, B2 =>
                           n120112, ZN => n114942);
   U86256 : OAI22_X1 port map( A1 => n90521, A2 => n120118, B1 => n90040, B2 =>
                           n120112, ZN => n114914);
   U86257 : OAI22_X1 port map( A1 => n90520, A2 => n120118, B1 => n90039, B2 =>
                           n120112, ZN => n114886);
   U86258 : OAI22_X1 port map( A1 => n90519, A2 => n120118, B1 => n90038, B2 =>
                           n120112, ZN => n114858);
   U86259 : OAI22_X1 port map( A1 => n90518, A2 => n120118, B1 => n90037, B2 =>
                           n120112, ZN => n114830);
   U86260 : OAI22_X1 port map( A1 => n90517, A2 => n120118, B1 => n90036, B2 =>
                           n120112, ZN => n114802);
   U86261 : OAI22_X1 port map( A1 => n114233, A2 => n120114, B1 => n90095, B2 
                           => n120108, ZN => n116466);
   U86262 : OAI22_X1 port map( A1 => n114232, A2 => n120114, B1 => n90094, B2 
                           => n120108, ZN => n116426);
   U86263 : OAI22_X1 port map( A1 => n114231, A2 => n120114, B1 => n90093, B2 
                           => n120108, ZN => n116398);
   U86264 : OAI22_X1 port map( A1 => n114230, A2 => n120114, B1 => n90092, B2 
                           => n120108, ZN => n116370);
   U86265 : OAI22_X1 port map( A1 => n98771, A2 => n119916, B1 => n90430, B2 =>
                           n119910, ZN => n117798);
   U86266 : OAI22_X1 port map( A1 => n98770, A2 => n119916, B1 => n90429, B2 =>
                           n119910, ZN => n117776);
   U86267 : OAI22_X1 port map( A1 => n98769, A2 => n119916, B1 => n90428, B2 =>
                           n119910, ZN => n117754);
   U86268 : OAI22_X1 port map( A1 => n98768, A2 => n119916, B1 => n90427, B2 =>
                           n119910, ZN => n117732);
   U86269 : OAI22_X1 port map( A1 => n98778, A2 => n119916, B1 => n90437, B2 =>
                           n119910, ZN => n117964);
   U86270 : OAI22_X1 port map( A1 => n98777, A2 => n119916, B1 => n90436, B2 =>
                           n119910, ZN => n117930);
   U86271 : OAI22_X1 port map( A1 => n98776, A2 => n119916, B1 => n90435, B2 =>
                           n119910, ZN => n117908);
   U86272 : OAI22_X1 port map( A1 => n98775, A2 => n119916, B1 => n90434, B2 =>
                           n119910, ZN => n117886);
   U86273 : OAI22_X1 port map( A1 => n98774, A2 => n119916, B1 => n90433, B2 =>
                           n119910, ZN => n117864);
   U86274 : OAI22_X1 port map( A1 => n98773, A2 => n119916, B1 => n90432, B2 =>
                           n119910, ZN => n117842);
   U86275 : OAI22_X1 port map( A1 => n98772, A2 => n119916, B1 => n90431, B2 =>
                           n119910, ZN => n117820);
   U86276 : OAI22_X1 port map( A1 => n114229, A2 => n120114, B1 => n90091, B2 
                           => n120108, ZN => n116342);
   U86277 : OAI22_X1 port map( A1 => n114228, A2 => n120114, B1 => n90090, B2 
                           => n120108, ZN => n116314);
   U86278 : OAI22_X1 port map( A1 => n114227, A2 => n120114, B1 => n90089, B2 
                           => n120108, ZN => n116286);
   U86279 : OAI22_X1 port map( A1 => n114226, A2 => n120114, B1 => n90088, B2 
                           => n120108, ZN => n116258);
   U86280 : OAI22_X1 port map( A1 => n114225, A2 => n120114, B1 => n90087, B2 
                           => n120108, ZN => n116230);
   U86281 : OAI22_X1 port map( A1 => n114224, A2 => n120114, B1 => n90086, B2 
                           => n120108, ZN => n116202);
   U86282 : OAI22_X1 port map( A1 => n114223, A2 => n120114, B1 => n90085, B2 
                           => n120108, ZN => n116174);
   U86283 : OAI22_X1 port map( A1 => n114222, A2 => n120114, B1 => n90084, B2 
                           => n120108, ZN => n116146);
   U86284 : OAI22_X1 port map( A1 => n114221, A2 => n120115, B1 => n90083, B2 
                           => n120109, ZN => n116118);
   U86285 : OAI22_X1 port map( A1 => n114220, A2 => n120115, B1 => n90082, B2 
                           => n120109, ZN => n116090);
   U86286 : OAI22_X1 port map( A1 => n114219, A2 => n120115, B1 => n90081, B2 
                           => n120109, ZN => n116062);
   U86287 : OAI22_X1 port map( A1 => n114218, A2 => n120115, B1 => n90080, B2 
                           => n120109, ZN => n116034);
   U86288 : OAI22_X1 port map( A1 => n114217, A2 => n120115, B1 => n90079, B2 
                           => n120109, ZN => n116006);
   U86289 : OAI22_X1 port map( A1 => n114216, A2 => n120115, B1 => n90078, B2 
                           => n120109, ZN => n115978);
   U86290 : OAI22_X1 port map( A1 => n114215, A2 => n120115, B1 => n90077, B2 
                           => n120109, ZN => n115950);
   U86291 : OAI22_X1 port map( A1 => n90557, A2 => n120115, B1 => n90076, B2 =>
                           n120109, ZN => n115922);
   U86292 : OAI22_X1 port map( A1 => n90556, A2 => n120115, B1 => n90075, B2 =>
                           n120109, ZN => n115894);
   U86293 : OAI22_X1 port map( A1 => n90555, A2 => n120115, B1 => n90074, B2 =>
                           n120109, ZN => n115866);
   U86294 : OAI22_X1 port map( A1 => n90554, A2 => n120115, B1 => n90073, B2 =>
                           n120109, ZN => n115838);
   U86295 : OAI22_X1 port map( A1 => n90553, A2 => n120115, B1 => n90072, B2 =>
                           n120109, ZN => n115810);
   U86296 : OAI22_X1 port map( A1 => n90552, A2 => n120116, B1 => n90071, B2 =>
                           n120110, ZN => n115782);
   U86297 : OAI22_X1 port map( A1 => n90551, A2 => n120116, B1 => n90070, B2 =>
                           n120110, ZN => n115754);
   U86298 : OAI22_X1 port map( A1 => n90550, A2 => n120116, B1 => n90069, B2 =>
                           n120110, ZN => n115726);
   U86299 : OAI22_X1 port map( A1 => n90549, A2 => n120116, B1 => n90068, B2 =>
                           n120110, ZN => n115698);
   U86300 : OAI22_X1 port map( A1 => n90548, A2 => n120116, B1 => n90067, B2 =>
                           n120110, ZN => n115670);
   U86301 : OAI22_X1 port map( A1 => n90547, A2 => n120116, B1 => n90066, B2 =>
                           n120110, ZN => n115642);
   U86302 : OAI22_X1 port map( A1 => n90546, A2 => n120116, B1 => n90065, B2 =>
                           n120110, ZN => n115614);
   U86303 : OAI22_X1 port map( A1 => n90545, A2 => n120116, B1 => n90064, B2 =>
                           n120110, ZN => n115586);
   U86304 : OAI22_X1 port map( A1 => n90544, A2 => n120116, B1 => n90063, B2 =>
                           n120110, ZN => n115558);
   U86305 : OAI22_X1 port map( A1 => n90543, A2 => n120116, B1 => n90062, B2 =>
                           n120110, ZN => n115530);
   U86306 : OAI22_X1 port map( A1 => n90542, A2 => n120116, B1 => n90061, B2 =>
                           n120110, ZN => n115502);
   U86307 : OAI22_X1 port map( A1 => n90541, A2 => n120116, B1 => n90060, B2 =>
                           n120110, ZN => n115474);
   U86308 : OAI22_X1 port map( A1 => n90540, A2 => n120117, B1 => n90059, B2 =>
                           n120111, ZN => n115446);
   U86309 : OAI22_X1 port map( A1 => n90539, A2 => n120117, B1 => n90058, B2 =>
                           n120111, ZN => n115418);
   U86310 : OAI22_X1 port map( A1 => n90538, A2 => n120117, B1 => n90057, B2 =>
                           n120111, ZN => n115390);
   U86311 : OAI22_X1 port map( A1 => n90537, A2 => n120117, B1 => n90056, B2 =>
                           n120111, ZN => n115362);
   U86312 : OAI22_X1 port map( A1 => n90536, A2 => n120117, B1 => n90055, B2 =>
                           n120111, ZN => n115334);
   U86313 : OAI22_X1 port map( A1 => n90535, A2 => n120117, B1 => n90054, B2 =>
                           n120111, ZN => n115306);
   U86314 : OAI22_X1 port map( A1 => n90534, A2 => n120117, B1 => n90053, B2 =>
                           n120111, ZN => n115278);
   U86315 : OAI22_X1 port map( A1 => n90533, A2 => n120117, B1 => n90052, B2 =>
                           n120111, ZN => n115250);
   U86316 : OAI22_X1 port map( A1 => n90532, A2 => n120117, B1 => n90051, B2 =>
                           n120111, ZN => n115222);
   U86317 : OAI22_X1 port map( A1 => n90531, A2 => n120117, B1 => n90050, B2 =>
                           n120111, ZN => n115194);
   U86318 : OAI22_X1 port map( A1 => n90324, A2 => n120129, B1 => n114253, B2 
                           => n120123, ZN => n115167);
   U86319 : OAI22_X1 port map( A1 => n90323, A2 => n120129, B1 => n114252, B2 
                           => n120123, ZN => n115139);
   U86320 : OAI22_X1 port map( A1 => n90322, A2 => n120130, B1 => n114251, B2 
                           => n120124, ZN => n115111);
   U86321 : OAI22_X1 port map( A1 => n90321, A2 => n120130, B1 => n114250, B2 
                           => n120124, ZN => n115083);
   U86322 : OAI22_X1 port map( A1 => n90320, A2 => n120130, B1 => n114249, B2 
                           => n120124, ZN => n115055);
   U86323 : OAI22_X1 port map( A1 => n90319, A2 => n120130, B1 => n114248, B2 
                           => n120124, ZN => n115027);
   U86324 : OAI22_X1 port map( A1 => n90318, A2 => n120130, B1 => n114247, B2 
                           => n120124, ZN => n114999);
   U86325 : OAI22_X1 port map( A1 => n90317, A2 => n120130, B1 => n114246, B2 
                           => n120124, ZN => n114971);
   U86326 : OAI22_X1 port map( A1 => n90316, A2 => n120130, B1 => n114245, B2 
                           => n120124, ZN => n114943);
   U86327 : OAI22_X1 port map( A1 => n90315, A2 => n120130, B1 => n114244, B2 
                           => n120124, ZN => n114915);
   U86328 : OAI22_X1 port map( A1 => n90314, A2 => n120130, B1 => n114243, B2 
                           => n120124, ZN => n114887);
   U86329 : OAI22_X1 port map( A1 => n90313, A2 => n120130, B1 => n114242, B2 
                           => n120124, ZN => n114859);
   U86330 : OAI22_X1 port map( A1 => n90312, A2 => n120130, B1 => n114241, B2 
                           => n120124, ZN => n114831);
   U86331 : OAI22_X1 port map( A1 => n90311, A2 => n120130, B1 => n114240, B2 
                           => n120124, ZN => n114803);
   U86332 : OAI22_X1 port map( A1 => n90370, A2 => n120126, B1 => n114299, B2 
                           => n120120, ZN => n116467);
   U86333 : OAI22_X1 port map( A1 => n90369, A2 => n120126, B1 => n114298, B2 
                           => n120120, ZN => n116427);
   U86334 : OAI22_X1 port map( A1 => n90368, A2 => n120126, B1 => n114297, B2 
                           => n120120, ZN => n116399);
   U86335 : OAI22_X1 port map( A1 => n90367, A2 => n120126, B1 => n114296, B2 
                           => n120120, ZN => n116371);
   U86336 : OAI22_X1 port map( A1 => n90366, A2 => n120126, B1 => n114295, B2 
                           => n120120, ZN => n116343);
   U86337 : OAI22_X1 port map( A1 => n90365, A2 => n120126, B1 => n114294, B2 
                           => n120120, ZN => n116315);
   U86338 : OAI22_X1 port map( A1 => n90364, A2 => n120126, B1 => n114293, B2 
                           => n120120, ZN => n116287);
   U86339 : OAI22_X1 port map( A1 => n90363, A2 => n120126, B1 => n114292, B2 
                           => n120120, ZN => n116259);
   U86340 : OAI22_X1 port map( A1 => n90362, A2 => n120126, B1 => n114291, B2 
                           => n120120, ZN => n116231);
   U86341 : OAI22_X1 port map( A1 => n90361, A2 => n120126, B1 => n114290, B2 
                           => n120120, ZN => n116203);
   U86342 : OAI22_X1 port map( A1 => n90360, A2 => n120126, B1 => n114289, B2 
                           => n120120, ZN => n116175);
   U86343 : OAI22_X1 port map( A1 => n90359, A2 => n120126, B1 => n114288, B2 
                           => n120120, ZN => n116147);
   U86344 : OAI22_X1 port map( A1 => n90358, A2 => n120127, B1 => n114287, B2 
                           => n120121, ZN => n116119);
   U86345 : OAI22_X1 port map( A1 => n90357, A2 => n120127, B1 => n114286, B2 
                           => n120121, ZN => n116091);
   U86346 : OAI22_X1 port map( A1 => n90356, A2 => n120127, B1 => n114285, B2 
                           => n120121, ZN => n116063);
   U86347 : OAI22_X1 port map( A1 => n90355, A2 => n120127, B1 => n114284, B2 
                           => n120121, ZN => n116035);
   U86348 : OAI22_X1 port map( A1 => n90354, A2 => n120127, B1 => n114283, B2 
                           => n120121, ZN => n116007);
   U86349 : OAI22_X1 port map( A1 => n90353, A2 => n120127, B1 => n114282, B2 
                           => n120121, ZN => n115979);
   U86350 : OAI22_X1 port map( A1 => n90352, A2 => n120127, B1 => n114281, B2 
                           => n120121, ZN => n115951);
   U86351 : OAI22_X1 port map( A1 => n90351, A2 => n120127, B1 => n114280, B2 
                           => n120121, ZN => n115923);
   U86352 : OAI22_X1 port map( A1 => n90350, A2 => n120127, B1 => n114279, B2 
                           => n120121, ZN => n115895);
   U86353 : OAI22_X1 port map( A1 => n90349, A2 => n120127, B1 => n114278, B2 
                           => n120121, ZN => n115867);
   U86354 : OAI22_X1 port map( A1 => n90348, A2 => n120127, B1 => n114277, B2 
                           => n120121, ZN => n115839);
   U86355 : OAI22_X1 port map( A1 => n90347, A2 => n120127, B1 => n114276, B2 
                           => n120121, ZN => n115811);
   U86356 : OAI22_X1 port map( A1 => n90346, A2 => n120128, B1 => n114275, B2 
                           => n120122, ZN => n115783);
   U86357 : OAI22_X1 port map( A1 => n90345, A2 => n120128, B1 => n114274, B2 
                           => n120122, ZN => n115755);
   U86358 : OAI22_X1 port map( A1 => n90344, A2 => n120128, B1 => n114273, B2 
                           => n120122, ZN => n115727);
   U86359 : OAI22_X1 port map( A1 => n90343, A2 => n120128, B1 => n114272, B2 
                           => n120122, ZN => n115699);
   U86360 : OAI22_X1 port map( A1 => n90342, A2 => n120128, B1 => n114271, B2 
                           => n120122, ZN => n115671);
   U86361 : OAI22_X1 port map( A1 => n90341, A2 => n120128, B1 => n114270, B2 
                           => n120122, ZN => n115643);
   U86362 : OAI22_X1 port map( A1 => n90340, A2 => n120128, B1 => n114269, B2 
                           => n120122, ZN => n115615);
   U86363 : OAI22_X1 port map( A1 => n90339, A2 => n120128, B1 => n114268, B2 
                           => n120122, ZN => n115587);
   U86364 : OAI22_X1 port map( A1 => n90338, A2 => n120128, B1 => n114267, B2 
                           => n120122, ZN => n115559);
   U86365 : OAI22_X1 port map( A1 => n90337, A2 => n120128, B1 => n114266, B2 
                           => n120122, ZN => n115531);
   U86366 : OAI22_X1 port map( A1 => n90336, A2 => n120128, B1 => n114265, B2 
                           => n120122, ZN => n115503);
   U86367 : OAI22_X1 port map( A1 => n90335, A2 => n120128, B1 => n114264, B2 
                           => n120122, ZN => n115475);
   U86368 : OAI22_X1 port map( A1 => n90334, A2 => n120129, B1 => n114263, B2 
                           => n120123, ZN => n115447);
   U86369 : OAI22_X1 port map( A1 => n90333, A2 => n120129, B1 => n114262, B2 
                           => n120123, ZN => n115419);
   U86370 : OAI22_X1 port map( A1 => n90332, A2 => n120129, B1 => n114261, B2 
                           => n120123, ZN => n115391);
   U86371 : OAI22_X1 port map( A1 => n90331, A2 => n120129, B1 => n114260, B2 
                           => n120123, ZN => n115363);
   U86372 : OAI22_X1 port map( A1 => n90330, A2 => n120129, B1 => n114259, B2 
                           => n120123, ZN => n115335);
   U86373 : OAI22_X1 port map( A1 => n90329, A2 => n120129, B1 => n114258, B2 
                           => n120123, ZN => n115307);
   U86374 : OAI22_X1 port map( A1 => n90328, A2 => n120129, B1 => n114257, B2 
                           => n120123, ZN => n115279);
   U86375 : OAI22_X1 port map( A1 => n90327, A2 => n120129, B1 => n114256, B2 
                           => n120123, ZN => n115251);
   U86376 : OAI22_X1 port map( A1 => n90326, A2 => n120129, B1 => n114255, B2 
                           => n120123, ZN => n115223);
   U86377 : OAI22_X1 port map( A1 => n90325, A2 => n120129, B1 => n114254, B2 
                           => n120123, ZN => n115195);
   U86378 : OAI22_X1 port map( A1 => n98599, A2 => n120051, B1 => n114596, B2 
                           => n120045, ZN => n115173);
   U86379 : OAI22_X1 port map( A1 => n98598, A2 => n120051, B1 => n114595, B2 
                           => n120045, ZN => n115145);
   U86380 : OAI22_X1 port map( A1 => n98597, A2 => n120052, B1 => n114594, B2 
                           => n120046, ZN => n115117);
   U86381 : OAI22_X1 port map( A1 => n98596, A2 => n120052, B1 => n114593, B2 
                           => n120046, ZN => n115089);
   U86382 : OAI22_X1 port map( A1 => n98595, A2 => n120052, B1 => n114592, B2 
                           => n120046, ZN => n115061);
   U86383 : OAI22_X1 port map( A1 => n98594, A2 => n120052, B1 => n114591, B2 
                           => n120046, ZN => n115033);
   U86384 : OAI22_X1 port map( A1 => n98593, A2 => n120052, B1 => n114590, B2 
                           => n120046, ZN => n115005);
   U86385 : OAI22_X1 port map( A1 => n98592, A2 => n120052, B1 => n114589, B2 
                           => n120046, ZN => n114977);
   U86386 : OAI22_X1 port map( A1 => n98591, A2 => n120052, B1 => n114588, B2 
                           => n120046, ZN => n114949);
   U86387 : OAI22_X1 port map( A1 => n98590, A2 => n120052, B1 => n114587, B2 
                           => n120046, ZN => n114921);
   U86388 : OAI22_X1 port map( A1 => n98589, A2 => n120052, B1 => n114586, B2 
                           => n120046, ZN => n114893);
   U86389 : OAI22_X1 port map( A1 => n98588, A2 => n120052, B1 => n114585, B2 
                           => n120046, ZN => n114865);
   U86390 : OAI22_X1 port map( A1 => n98587, A2 => n120052, B1 => n114584, B2 
                           => n120046, ZN => n114837);
   U86391 : OAI22_X1 port map( A1 => n98586, A2 => n120052, B1 => n114583, B2 
                           => n120046, ZN => n114809);
   U86392 : OAI22_X1 port map( A1 => n98645, A2 => n120048, B1 => n114642, B2 
                           => n120042, ZN => n116477);
   U86393 : OAI22_X1 port map( A1 => n98644, A2 => n120048, B1 => n114641, B2 
                           => n120042, ZN => n116433);
   U86394 : OAI22_X1 port map( A1 => n98643, A2 => n120048, B1 => n114640, B2 
                           => n120042, ZN => n116405);
   U86395 : OAI22_X1 port map( A1 => n98642, A2 => n120048, B1 => n114639, B2 
                           => n120042, ZN => n116377);
   U86396 : OAI22_X1 port map( A1 => n98641, A2 => n120048, B1 => n114638, B2 
                           => n120042, ZN => n116349);
   U86397 : OAI22_X1 port map( A1 => n98640, A2 => n120048, B1 => n114637, B2 
                           => n120042, ZN => n116321);
   U86398 : OAI22_X1 port map( A1 => n98639, A2 => n120048, B1 => n114636, B2 
                           => n120042, ZN => n116293);
   U86399 : OAI22_X1 port map( A1 => n98638, A2 => n120048, B1 => n114635, B2 
                           => n120042, ZN => n116265);
   U86400 : OAI22_X1 port map( A1 => n98637, A2 => n120048, B1 => n114634, B2 
                           => n120042, ZN => n116237);
   U86401 : OAI22_X1 port map( A1 => n98636, A2 => n120048, B1 => n114633, B2 
                           => n120042, ZN => n116209);
   U86402 : OAI22_X1 port map( A1 => n98635, A2 => n120048, B1 => n114632, B2 
                           => n120042, ZN => n116181);
   U86403 : OAI22_X1 port map( A1 => n98634, A2 => n120048, B1 => n114631, B2 
                           => n120042, ZN => n116153);
   U86404 : OAI22_X1 port map( A1 => n98633, A2 => n120049, B1 => n114630, B2 
                           => n120043, ZN => n116125);
   U86405 : OAI22_X1 port map( A1 => n98632, A2 => n120049, B1 => n114629, B2 
                           => n120043, ZN => n116097);
   U86406 : OAI22_X1 port map( A1 => n98631, A2 => n120049, B1 => n114628, B2 
                           => n120043, ZN => n116069);
   U86407 : OAI22_X1 port map( A1 => n98630, A2 => n120049, B1 => n114627, B2 
                           => n120043, ZN => n116041);
   U86408 : OAI22_X1 port map( A1 => n98629, A2 => n120049, B1 => n114626, B2 
                           => n120043, ZN => n116013);
   U86409 : OAI22_X1 port map( A1 => n98628, A2 => n120049, B1 => n114625, B2 
                           => n120043, ZN => n115985);
   U86410 : OAI22_X1 port map( A1 => n98627, A2 => n120049, B1 => n114624, B2 
                           => n120043, ZN => n115957);
   U86411 : OAI22_X1 port map( A1 => n98626, A2 => n120049, B1 => n114623, B2 
                           => n120043, ZN => n115929);
   U86412 : OAI22_X1 port map( A1 => n98625, A2 => n120049, B1 => n114622, B2 
                           => n120043, ZN => n115901);
   U86413 : OAI22_X1 port map( A1 => n98624, A2 => n120049, B1 => n114621, B2 
                           => n120043, ZN => n115873);
   U86414 : OAI22_X1 port map( A1 => n98623, A2 => n120049, B1 => n114620, B2 
                           => n120043, ZN => n115845);
   U86415 : OAI22_X1 port map( A1 => n98622, A2 => n120049, B1 => n114619, B2 
                           => n120043, ZN => n115817);
   U86416 : OAI22_X1 port map( A1 => n98621, A2 => n120050, B1 => n114618, B2 
                           => n120044, ZN => n115789);
   U86417 : OAI22_X1 port map( A1 => n98620, A2 => n120050, B1 => n114617, B2 
                           => n120044, ZN => n115761);
   U86418 : OAI22_X1 port map( A1 => n98619, A2 => n120050, B1 => n114616, B2 
                           => n120044, ZN => n115733);
   U86419 : OAI22_X1 port map( A1 => n98618, A2 => n120050, B1 => n114615, B2 
                           => n120044, ZN => n115705);
   U86420 : OAI22_X1 port map( A1 => n98617, A2 => n120050, B1 => n114614, B2 
                           => n120044, ZN => n115677);
   U86421 : OAI22_X1 port map( A1 => n98616, A2 => n120050, B1 => n114613, B2 
                           => n120044, ZN => n115649);
   U86422 : OAI22_X1 port map( A1 => n98615, A2 => n120050, B1 => n114612, B2 
                           => n120044, ZN => n115621);
   U86423 : OAI22_X1 port map( A1 => n98614, A2 => n120050, B1 => n114611, B2 
                           => n120044, ZN => n115593);
   U86424 : OAI22_X1 port map( A1 => n98613, A2 => n120050, B1 => n114610, B2 
                           => n120044, ZN => n115565);
   U86425 : OAI22_X1 port map( A1 => n98612, A2 => n120050, B1 => n114609, B2 
                           => n120044, ZN => n115537);
   U86426 : OAI22_X1 port map( A1 => n98611, A2 => n120050, B1 => n114608, B2 
                           => n120044, ZN => n115509);
   U86427 : OAI22_X1 port map( A1 => n98610, A2 => n120050, B1 => n114607, B2 
                           => n120044, ZN => n115481);
   U86428 : OAI22_X1 port map( A1 => n98609, A2 => n120051, B1 => n114606, B2 
                           => n120045, ZN => n115453);
   U86429 : OAI22_X1 port map( A1 => n98608, A2 => n120051, B1 => n114605, B2 
                           => n120045, ZN => n115425);
   U86430 : OAI22_X1 port map( A1 => n98607, A2 => n120051, B1 => n114604, B2 
                           => n120045, ZN => n115397);
   U86431 : OAI22_X1 port map( A1 => n98606, A2 => n120051, B1 => n114603, B2 
                           => n120045, ZN => n115369);
   U86432 : OAI22_X1 port map( A1 => n98605, A2 => n120051, B1 => n114602, B2 
                           => n120045, ZN => n115341);
   U86433 : OAI22_X1 port map( A1 => n98604, A2 => n120051, B1 => n114601, B2 
                           => n120045, ZN => n115313);
   U86434 : OAI22_X1 port map( A1 => n98603, A2 => n120051, B1 => n114600, B2 
                           => n120045, ZN => n115285);
   U86435 : OAI22_X1 port map( A1 => n98602, A2 => n120051, B1 => n114599, B2 
                           => n120045, ZN => n115257);
   U86436 : OAI22_X1 port map( A1 => n98601, A2 => n120051, B1 => n114598, B2 
                           => n120045, ZN => n115229);
   U86437 : OAI22_X1 port map( A1 => n98600, A2 => n120051, B1 => n114597, B2 
                           => n120045, ZN => n115201);
   U86438 : OAI22_X1 port map( A1 => n89500, A2 => n120829, B1 => n120826, B2 
                           => n120809, ZN => n7483);
   U86439 : OAI22_X1 port map( A1 => n89498, A2 => n120829, B1 => n120826, B2 
                           => n120812, ZN => n7484);
   U86440 : OAI22_X1 port map( A1 => n89496, A2 => n120829, B1 => n120826, B2 
                           => n120815, ZN => n7485);
   U86441 : OAI22_X1 port map( A1 => n89493, A2 => n120829, B1 => n120826, B2 
                           => n120818, ZN => n7486);
   U86442 : OAI22_X1 port map( A1 => n120622, A2 => n113900, B1 => n120809, B2 
                           => n120616, ZN => n7419);
   U86443 : OAI22_X1 port map( A1 => n120622, A2 => n113899, B1 => n120812, B2 
                           => n120616, ZN => n7420);
   U86444 : OAI22_X1 port map( A1 => n120622, A2 => n113898, B1 => n120815, B2 
                           => n120616, ZN => n7421);
   U86445 : OAI22_X1 port map( A1 => n120622, A2 => n113896, B1 => n120818, B2 
                           => n120616, ZN => n7422);
   U86446 : OAI22_X1 port map( A1 => n99183, A2 => n120475, B1 => n120810, B2 
                           => n120469, ZN => n6651);
   U86447 : OAI22_X1 port map( A1 => n99182, A2 => n120475, B1 => n120813, B2 
                           => n120469, ZN => n6652);
   U86448 : OAI22_X1 port map( A1 => n99181, A2 => n120475, B1 => n120816, B2 
                           => n120469, ZN => n6653);
   U86449 : OAI22_X1 port map( A1 => n99179, A2 => n120475, B1 => n120819, B2 
                           => n120469, ZN => n6654);
   U86450 : OAI22_X1 port map( A1 => n99315, A2 => n120451, B1 => n120810, B2 
                           => n120445, ZN => n6523);
   U86451 : OAI22_X1 port map( A1 => n99314, A2 => n120451, B1 => n120813, B2 
                           => n120445, ZN => n6524);
   U86452 : OAI22_X1 port map( A1 => n99313, A2 => n120451, B1 => n120816, B2 
                           => n120445, ZN => n6525);
   U86453 : OAI22_X1 port map( A1 => n99311, A2 => n120451, B1 => n120819, B2 
                           => n120445, ZN => n6526);
   U86454 : OAI22_X1 port map( A1 => n120524, A2 => n114060, B1 => n120809, B2 
                           => n120517, ZN => n6907);
   U86455 : OAI22_X1 port map( A1 => n120524, A2 => n114059, B1 => n120812, B2 
                           => n120517, ZN => n6908);
   U86456 : OAI22_X1 port map( A1 => n120524, A2 => n114058, B1 => n120815, B2 
                           => n120517, ZN => n6909);
   U86457 : OAI22_X1 port map( A1 => n120524, A2 => n114056, B1 => n120818, B2 
                           => n120517, ZN => n6910);
   U86458 : OAI22_X1 port map( A1 => n99051, A2 => n120499, B1 => n120809, B2 
                           => n120493, ZN => n6779);
   U86459 : OAI22_X1 port map( A1 => n99050, A2 => n120499, B1 => n120812, B2 
                           => n120493, ZN => n6780);
   U86460 : OAI22_X1 port map( A1 => n99049, A2 => n120499, B1 => n120815, B2 
                           => n120493, ZN => n6781);
   U86461 : OAI22_X1 port map( A1 => n99047, A2 => n120499, B1 => n120818, B2 
                           => n120493, ZN => n6782);
   U86462 : OAI22_X1 port map( A1 => n99117, A2 => n120487, B1 => n120810, B2 
                           => n120481, ZN => n6715);
   U86463 : OAI22_X1 port map( A1 => n99116, A2 => n120487, B1 => n120813, B2 
                           => n120481, ZN => n6716);
   U86464 : OAI22_X1 port map( A1 => n99115, A2 => n120487, B1 => n120816, B2 
                           => n120481, ZN => n6717);
   U86465 : OAI22_X1 port map( A1 => n99113, A2 => n120487, B1 => n120819, B2 
                           => n120481, ZN => n6718);
   U86466 : OAI22_X1 port map( A1 => n99249, A2 => n120463, B1 => n120810, B2 
                           => n120457, ZN => n6587);
   U86467 : OAI22_X1 port map( A1 => n99248, A2 => n120463, B1 => n120813, B2 
                           => n120457, ZN => n6588);
   U86468 : OAI22_X1 port map( A1 => n99247, A2 => n120463, B1 => n120816, B2 
                           => n120457, ZN => n6589);
   U86469 : OAI22_X1 port map( A1 => n99245, A2 => n120463, B1 => n120819, B2 
                           => n120457, ZN => n6590);
   U86470 : OAI22_X1 port map( A1 => n98718, A2 => n120586, B1 => n120809, B2 
                           => n120580, ZN => n7227);
   U86471 : OAI22_X1 port map( A1 => n98717, A2 => n120586, B1 => n120812, B2 
                           => n120580, ZN => n7228);
   U86472 : OAI22_X1 port map( A1 => n98716, A2 => n120586, B1 => n120815, B2 
                           => n120580, ZN => n7229);
   U86473 : OAI22_X1 port map( A1 => n98714, A2 => n120586, B1 => n120818, B2 
                           => n120580, ZN => n7230);
   U86474 : OAI22_X1 port map( A1 => n98652, A2 => n120598, B1 => n120809, B2 
                           => n120592, ZN => n7291);
   U86475 : OAI22_X1 port map( A1 => n98651, A2 => n120598, B1 => n120812, B2 
                           => n120592, ZN => n7292);
   U86476 : OAI22_X1 port map( A1 => n98650, A2 => n120598, B1 => n120815, B2 
                           => n120592, ZN => n7293);
   U86477 : OAI22_X1 port map( A1 => n98648, A2 => n120598, B1 => n120818, B2 
                           => n120592, ZN => n7294);
   U86478 : OAI22_X1 port map( A1 => n99584, A2 => n120365, B1 => n120810, B2 
                           => n120359, ZN => n6075);
   U86479 : OAI22_X1 port map( A1 => n99583, A2 => n120365, B1 => n120813, B2 
                           => n120359, ZN => n6076);
   U86480 : OAI22_X1 port map( A1 => n99582, A2 => n120365, B1 => n120816, B2 
                           => n120359, ZN => n6077);
   U86481 : OAI22_X1 port map( A1 => n99580, A2 => n120365, B1 => n120819, B2 
                           => n120359, ZN => n6078);
   U86482 : OAI22_X1 port map( A1 => n120341, A2 => n114310, B1 => n120810, B2 
                           => n120334, ZN => n5947);
   U86483 : OAI22_X1 port map( A1 => n120341, A2 => n114309, B1 => n120813, B2 
                           => n120334, ZN => n5948);
   U86484 : OAI22_X1 port map( A1 => n120341, A2 => n114308, B1 => n120816, B2 
                           => n120334, ZN => n5949);
   U86485 : OAI22_X1 port map( A1 => n120341, A2 => n114306, B1 => n120819, B2 
                           => n120334, ZN => n5950);
   U86486 : OAI22_X1 port map( A1 => n99450, A2 => n120402, B1 => n120810, B2 
                           => n120396, ZN => n6267);
   U86487 : OAI22_X1 port map( A1 => n99449, A2 => n120402, B1 => n120813, B2 
                           => n120396, ZN => n6268);
   U86488 : OAI22_X1 port map( A1 => n99448, A2 => n120402, B1 => n120816, B2 
                           => n120396, ZN => n6269);
   U86489 : OAI22_X1 port map( A1 => n99446, A2 => n120402, B1 => n120819, B2 
                           => n120396, ZN => n6270);
   U86490 : OAI22_X1 port map( A1 => n99720, A2 => n120328, B1 => n120811, B2 
                           => n120322, ZN => n5883);
   U86491 : OAI22_X1 port map( A1 => n99719, A2 => n120328, B1 => n120814, B2 
                           => n120322, ZN => n5884);
   U86492 : OAI22_X1 port map( A1 => n99718, A2 => n120328, B1 => n120817, B2 
                           => n120322, ZN => n5885);
   U86493 : OAI22_X1 port map( A1 => n99716, A2 => n120328, B1 => n120820, B2 
                           => n120322, ZN => n5886);
   U86494 : OAI22_X1 port map( A1 => n99918, A2 => n120277, B1 => n120811, B2 
                           => n120271, ZN => n5627);
   U86495 : OAI22_X1 port map( A1 => n99917, A2 => n120277, B1 => n120814, B2 
                           => n120271, ZN => n5628);
   U86496 : OAI22_X1 port map( A1 => n99916, A2 => n120277, B1 => n120817, B2 
                           => n120271, ZN => n5629);
   U86497 : OAI22_X1 port map( A1 => n99914, A2 => n120277, B1 => n120820, B2 
                           => n120271, ZN => n5630);
   U86498 : OAI22_X1 port map( A1 => n90035, A2 => n120536, B1 => n120809, B2 
                           => n120530, ZN => n6971);
   U86499 : OAI22_X1 port map( A1 => n90034, A2 => n120536, B1 => n120812, B2 
                           => n120530, ZN => n6972);
   U86500 : OAI22_X1 port map( A1 => n90033, A2 => n120536, B1 => n120815, B2 
                           => n120530, ZN => n6973);
   U86501 : OAI22_X1 port map( A1 => n90031, A2 => n120536, B1 => n120818, B2 
                           => n120530, ZN => n6974);
   U86502 : OAI22_X1 port map( A1 => n89969, A2 => n120545, B1 => n120809, B2 
                           => n120542, ZN => n7035);
   U86503 : OAI22_X1 port map( A1 => n89968, A2 => n120545, B1 => n120812, B2 
                           => n120542, ZN => n7036);
   U86504 : OAI22_X1 port map( A1 => n89967, A2 => n120545, B1 => n120815, B2 
                           => n120542, ZN => n7037);
   U86505 : OAI22_X1 port map( A1 => n89965, A2 => n120545, B1 => n120818, B2 
                           => n120542, ZN => n7038);
   U86506 : OAI22_X1 port map( A1 => n90516, A2 => n120385, B1 => n120810, B2 
                           => n120384, ZN => n6203);
   U86507 : OAI22_X1 port map( A1 => n90515, A2 => n120385, B1 => n120813, B2 
                           => n120384, ZN => n6204);
   U86508 : OAI22_X1 port map( A1 => n90514, A2 => n120385, B1 => n120816, B2 
                           => n120384, ZN => n6205);
   U86509 : OAI22_X1 port map( A1 => n90512, A2 => n120387, B1 => n120819, B2 
                           => n120384, ZN => n6206);
   U86510 : OAI22_X1 port map( A1 => n90310, A2 => n120439, B1 => n120810, B2 
                           => n120433, ZN => n6459);
   U86511 : OAI22_X1 port map( A1 => n90309, A2 => n120439, B1 => n120813, B2 
                           => n120433, ZN => n6460);
   U86512 : OAI22_X1 port map( A1 => n90308, A2 => n120439, B1 => n120816, B2 
                           => n120433, ZN => n6461);
   U86513 : OAI22_X1 port map( A1 => n90306, A2 => n120439, B1 => n120819, B2 
                           => n120433, ZN => n6462);
   U86514 : OAI22_X1 port map( A1 => n90377, A2 => n120427, B1 => n120810, B2 
                           => n120421, ZN => n6395);
   U86515 : OAI22_X1 port map( A1 => n90376, A2 => n120427, B1 => n120813, B2 
                           => n120421, ZN => n6396);
   U86516 : OAI22_X1 port map( A1 => n90375, A2 => n120427, B1 => n120816, B2 
                           => n120421, ZN => n6397);
   U86517 : OAI22_X1 port map( A1 => n90373, A2 => n120427, B1 => n120819, B2 
                           => n120421, ZN => n6398);
   U86518 : OAI22_X1 port map( A1 => n90715, A2 => n120353, B1 => n120810, B2 
                           => n120347, ZN => n6011);
   U86519 : OAI22_X1 port map( A1 => n90714, A2 => n120353, B1 => n120813, B2 
                           => n120347, ZN => n6012);
   U86520 : OAI22_X1 port map( A1 => n90713, A2 => n120353, B1 => n120816, B2 
                           => n120347, ZN => n6013);
   U86521 : OAI22_X1 port map( A1 => n90711, A2 => n120353, B1 => n120819, B2 
                           => n120347, ZN => n6014);
   U86522 : AOI22_X1 port map( A1 => n119976, A2 => n118922, B1 => n119970, B2 
                           => n111007, ZN => n117706);
   U86523 : AOI22_X1 port map( A1 => n120024, A2 => n118862, B1 => n120022, B2 
                           => OUT2_11_port, ZN => n117701);
   U86524 : AOI22_X1 port map( A1 => n119952, A2 => n118336, B1 => n119946, B2 
                           => n118216, ZN => n117708);
   U86525 : AOI22_X1 port map( A1 => n119977, A2 => n118923, B1 => n119971, B2 
                           => n111008, ZN => n117684);
   U86526 : AOI22_X1 port map( A1 => n120025, A2 => n118863, B1 => n120022, B2 
                           => OUT2_12_port, ZN => n117679);
   U86527 : AOI22_X1 port map( A1 => n119953, A2 => n118337, B1 => n119947, B2 
                           => n118217, ZN => n117686);
   U86528 : AOI22_X1 port map( A1 => n119977, A2 => n118924, B1 => n119971, B2 
                           => n111009, ZN => n117662);
   U86529 : AOI22_X1 port map( A1 => n120025, A2 => n118864, B1 => n120022, B2 
                           => OUT2_13_port, ZN => n117657);
   U86530 : AOI22_X1 port map( A1 => n119953, A2 => n118338, B1 => n119947, B2 
                           => n118218, ZN => n117664);
   U86531 : AOI22_X1 port map( A1 => n119977, A2 => n118925, B1 => n119971, B2 
                           => n111010, ZN => n117640);
   U86532 : AOI22_X1 port map( A1 => n120025, A2 => n118865, B1 => n120022, B2 
                           => OUT2_14_port, ZN => n117635);
   U86533 : AOI22_X1 port map( A1 => n119953, A2 => n118339, B1 => n119947, B2 
                           => n118219, ZN => n117642);
   U86534 : AOI22_X1 port map( A1 => n119977, A2 => n118926, B1 => n119971, B2 
                           => n111011, ZN => n117618);
   U86535 : AOI22_X1 port map( A1 => n120025, A2 => n118866, B1 => n120022, B2 
                           => OUT2_15_port, ZN => n117613);
   U86536 : AOI22_X1 port map( A1 => n119953, A2 => n118340, B1 => n119947, B2 
                           => n118220, ZN => n117620);
   U86537 : AOI22_X1 port map( A1 => n119977, A2 => n118927, B1 => n119971, B2 
                           => n111012, ZN => n117596);
   U86538 : AOI22_X1 port map( A1 => n120025, A2 => n118867, B1 => n120022, B2 
                           => OUT2_16_port, ZN => n117591);
   U86539 : AOI22_X1 port map( A1 => n119953, A2 => n118341, B1 => n119947, B2 
                           => n118221, ZN => n117598);
   U86540 : AOI22_X1 port map( A1 => n119977, A2 => n118928, B1 => n119971, B2 
                           => n111013, ZN => n117574);
   U86541 : AOI22_X1 port map( A1 => n120025, A2 => n118868, B1 => n120021, B2 
                           => OUT2_17_port, ZN => n117569);
   U86542 : AOI22_X1 port map( A1 => n119953, A2 => n118342, B1 => n119947, B2 
                           => n118222, ZN => n117576);
   U86543 : AOI22_X1 port map( A1 => n119977, A2 => n118929, B1 => n119971, B2 
                           => n111014, ZN => n117552);
   U86544 : AOI22_X1 port map( A1 => n120025, A2 => n118869, B1 => n120021, B2 
                           => OUT2_18_port, ZN => n117547);
   U86545 : AOI22_X1 port map( A1 => n119953, A2 => n118343, B1 => n119947, B2 
                           => n118223, ZN => n117554);
   U86546 : AOI22_X1 port map( A1 => n119977, A2 => n118930, B1 => n119971, B2 
                           => n111015, ZN => n117529);
   U86547 : AOI22_X1 port map( A1 => n120025, A2 => n118870, B1 => n120021, B2 
                           => OUT2_19_port, ZN => n117524);
   U86548 : AOI22_X1 port map( A1 => n119953, A2 => n118344, B1 => n119947, B2 
                           => n118224, ZN => n117531);
   U86549 : AOI22_X1 port map( A1 => n119977, A2 => n118931, B1 => n119971, B2 
                           => n111016, ZN => n117506);
   U86550 : AOI22_X1 port map( A1 => n120025, A2 => n118871, B1 => n120021, B2 
                           => OUT2_20_port, ZN => n117501);
   U86551 : AOI22_X1 port map( A1 => n119953, A2 => n118345, B1 => n119947, B2 
                           => n118225, ZN => n117508);
   U86552 : AOI22_X1 port map( A1 => n119977, A2 => n118932, B1 => n119971, B2 
                           => n111017, ZN => n117483);
   U86553 : AOI22_X1 port map( A1 => n120025, A2 => n118872, B1 => n120021, B2 
                           => OUT2_21_port, ZN => n117478);
   U86554 : AOI22_X1 port map( A1 => n119953, A2 => n118346, B1 => n119947, B2 
                           => n118226, ZN => n117485);
   U86555 : AOI22_X1 port map( A1 => n119977, A2 => n118933, B1 => n119971, B2 
                           => n111018, ZN => n117460);
   U86556 : AOI22_X1 port map( A1 => n120025, A2 => n118873, B1 => n120021, B2 
                           => OUT2_22_port, ZN => n117455);
   U86557 : AOI22_X1 port map( A1 => n119953, A2 => n118347, B1 => n119947, B2 
                           => n118227, ZN => n117462);
   U86558 : AOI22_X1 port map( A1 => n119977, A2 => n118934, B1 => n119971, B2 
                           => n111019, ZN => n117437);
   U86559 : AOI22_X1 port map( A1 => n120025, A2 => n118874, B1 => n120021, B2 
                           => OUT2_23_port, ZN => n117432);
   U86560 : AOI22_X1 port map( A1 => n119953, A2 => n118348, B1 => n119947, B2 
                           => n118228, ZN => n117439);
   U86561 : AOI22_X1 port map( A1 => n119978, A2 => n118935, B1 => n119972, B2 
                           => n111020, ZN => n117414);
   U86562 : AOI22_X1 port map( A1 => n120026, A2 => n118875, B1 => n120021, B2 
                           => OUT2_24_port, ZN => n117409);
   U86563 : AOI22_X1 port map( A1 => n119954, A2 => n118349, B1 => n119948, B2 
                           => n118229, ZN => n117416);
   U86564 : AOI22_X1 port map( A1 => n119978, A2 => n118936, B1 => n119972, B2 
                           => n111021, ZN => n117391);
   U86565 : AOI22_X1 port map( A1 => n120026, A2 => n118876, B1 => n120021, B2 
                           => OUT2_25_port, ZN => n117386);
   U86566 : AOI22_X1 port map( A1 => n119954, A2 => n118350, B1 => n119948, B2 
                           => n118230, ZN => n117393);
   U86567 : AOI22_X1 port map( A1 => n119978, A2 => n118937, B1 => n119972, B2 
                           => n111022, ZN => n117368);
   U86568 : AOI22_X1 port map( A1 => n120026, A2 => n118877, B1 => n120021, B2 
                           => OUT2_26_port, ZN => n117363);
   U86569 : AOI22_X1 port map( A1 => n119954, A2 => n118351, B1 => n119948, B2 
                           => n118231, ZN => n117370);
   U86570 : AOI22_X1 port map( A1 => n119978, A2 => n118938, B1 => n119972, B2 
                           => n111023, ZN => n117345);
   U86571 : AOI22_X1 port map( A1 => n120026, A2 => n118878, B1 => n120021, B2 
                           => OUT2_27_port, ZN => n117340);
   U86572 : AOI22_X1 port map( A1 => n119954, A2 => n118352, B1 => n119948, B2 
                           => n118232, ZN => n117347);
   U86573 : AOI22_X1 port map( A1 => n119978, A2 => n118939, B1 => n119972, B2 
                           => n111024, ZN => n117322);
   U86574 : AOI22_X1 port map( A1 => n120026, A2 => n118879, B1 => n120021, B2 
                           => OUT2_28_port, ZN => n117317);
   U86575 : AOI22_X1 port map( A1 => n119954, A2 => n118353, B1 => n119948, B2 
                           => n118233, ZN => n117324);
   U86576 : AOI22_X1 port map( A1 => n119978, A2 => n118940, B1 => n119972, B2 
                           => n111025, ZN => n117299);
   U86577 : AOI22_X1 port map( A1 => n120026, A2 => n118880, B1 => n120021, B2 
                           => OUT2_29_port, ZN => n117294);
   U86578 : AOI22_X1 port map( A1 => n119954, A2 => n118354, B1 => n119948, B2 
                           => n118234, ZN => n117301);
   U86579 : AOI22_X1 port map( A1 => n119978, A2 => n118941, B1 => n119972, B2 
                           => n111026, ZN => n117276);
   U86580 : AOI22_X1 port map( A1 => n120026, A2 => n118881, B1 => n120020, B2 
                           => OUT2_30_port, ZN => n117271);
   U86581 : AOI22_X1 port map( A1 => n119954, A2 => n118355, B1 => n119948, B2 
                           => n118235, ZN => n117278);
   U86582 : AOI22_X1 port map( A1 => n119978, A2 => n118942, B1 => n119972, B2 
                           => n111027, ZN => n117253);
   U86583 : AOI22_X1 port map( A1 => n120026, A2 => n118882, B1 => n120020, B2 
                           => OUT2_31_port, ZN => n117248);
   U86584 : AOI22_X1 port map( A1 => n119954, A2 => n118356, B1 => n119948, B2 
                           => n118236, ZN => n117255);
   U86585 : AOI22_X1 port map( A1 => n119978, A2 => n118943, B1 => n119972, B2 
                           => n111028, ZN => n117230);
   U86586 : AOI22_X1 port map( A1 => n120026, A2 => n118883, B1 => n120020, B2 
                           => OUT2_32_port, ZN => n117225);
   U86587 : AOI22_X1 port map( A1 => n119954, A2 => n118357, B1 => n119948, B2 
                           => n118237, ZN => n117232);
   U86588 : AOI22_X1 port map( A1 => n119978, A2 => n118944, B1 => n119972, B2 
                           => n111029, ZN => n117207);
   U86589 : AOI22_X1 port map( A1 => n120026, A2 => n118884, B1 => n120020, B2 
                           => OUT2_33_port, ZN => n117202);
   U86590 : AOI22_X1 port map( A1 => n119954, A2 => n118358, B1 => n119948, B2 
                           => n118238, ZN => n117209);
   U86591 : AOI22_X1 port map( A1 => n119978, A2 => n118945, B1 => n119972, B2 
                           => n111030, ZN => n117184);
   U86592 : AOI22_X1 port map( A1 => n120026, A2 => n118885, B1 => n120020, B2 
                           => OUT2_34_port, ZN => n117179);
   U86593 : AOI22_X1 port map( A1 => n119954, A2 => n118359, B1 => n119948, B2 
                           => n118239, ZN => n117186);
   U86594 : AOI22_X1 port map( A1 => n119978, A2 => n118946, B1 => n119972, B2 
                           => n111031, ZN => n117161);
   U86595 : AOI22_X1 port map( A1 => n120026, A2 => n118886, B1 => n120020, B2 
                           => OUT2_35_port, ZN => n117156);
   U86596 : AOI22_X1 port map( A1 => n119954, A2 => n118360, B1 => n119948, B2 
                           => n118240, ZN => n117163);
   U86597 : AOI22_X1 port map( A1 => n119979, A2 => n118947, B1 => n119973, B2 
                           => n111032, ZN => n117138);
   U86598 : AOI22_X1 port map( A1 => n120027, A2 => n118887, B1 => n120020, B2 
                           => OUT2_36_port, ZN => n117133);
   U86599 : AOI22_X1 port map( A1 => n119955, A2 => n118361, B1 => n119949, B2 
                           => n118241, ZN => n117140);
   U86600 : AOI22_X1 port map( A1 => n119979, A2 => n118948, B1 => n119973, B2 
                           => n111033, ZN => n117115);
   U86601 : AOI22_X1 port map( A1 => n120027, A2 => n118888, B1 => n120020, B2 
                           => OUT2_37_port, ZN => n117110);
   U86602 : AOI22_X1 port map( A1 => n119955, A2 => n118362, B1 => n119949, B2 
                           => n118242, ZN => n117117);
   U86603 : AOI22_X1 port map( A1 => n119979, A2 => n118949, B1 => n119973, B2 
                           => n111034, ZN => n117092);
   U86604 : AOI22_X1 port map( A1 => n120027, A2 => n118889, B1 => n120020, B2 
                           => OUT2_38_port, ZN => n117087);
   U86605 : AOI22_X1 port map( A1 => n119955, A2 => n118363, B1 => n119949, B2 
                           => n118243, ZN => n117094);
   U86606 : AOI22_X1 port map( A1 => n119979, A2 => n118950, B1 => n119973, B2 
                           => n111035, ZN => n117069);
   U86607 : AOI22_X1 port map( A1 => n120027, A2 => n118890, B1 => n120020, B2 
                           => OUT2_39_port, ZN => n117064);
   U86608 : AOI22_X1 port map( A1 => n119955, A2 => n118364, B1 => n119949, B2 
                           => n118244, ZN => n117071);
   U86609 : AOI22_X1 port map( A1 => n119979, A2 => n118951, B1 => n119973, B2 
                           => n111036, ZN => n117046);
   U86610 : AOI22_X1 port map( A1 => n120027, A2 => n118891, B1 => n120020, B2 
                           => OUT2_40_port, ZN => n117041);
   U86611 : AOI22_X1 port map( A1 => n119955, A2 => n118365, B1 => n119949, B2 
                           => n118245, ZN => n117048);
   U86612 : AOI22_X1 port map( A1 => n119979, A2 => n118952, B1 => n119973, B2 
                           => n111037, ZN => n117023);
   U86613 : AOI22_X1 port map( A1 => n120027, A2 => n118892, B1 => n120020, B2 
                           => OUT2_41_port, ZN => n117018);
   U86614 : AOI22_X1 port map( A1 => n119955, A2 => n118366, B1 => n119949, B2 
                           => n118246, ZN => n117025);
   U86615 : AOI22_X1 port map( A1 => n119979, A2 => n118953, B1 => n119973, B2 
                           => n111038, ZN => n117000);
   U86616 : AOI22_X1 port map( A1 => n120027, A2 => n118893, B1 => n120019, B2 
                           => OUT2_42_port, ZN => n116995);
   U86617 : AOI22_X1 port map( A1 => n119955, A2 => n118367, B1 => n119949, B2 
                           => n118247, ZN => n117002);
   U86618 : AOI22_X1 port map( A1 => n119979, A2 => n118954, B1 => n119973, B2 
                           => n111039, ZN => n116977);
   U86619 : AOI22_X1 port map( A1 => n120027, A2 => n118894, B1 => n120019, B2 
                           => OUT2_43_port, ZN => n116972);
   U86620 : AOI22_X1 port map( A1 => n119955, A2 => n118368, B1 => n119949, B2 
                           => n118248, ZN => n116979);
   U86621 : AOI22_X1 port map( A1 => n119979, A2 => n118955, B1 => n119973, B2 
                           => n111040, ZN => n116954);
   U86622 : AOI22_X1 port map( A1 => n120027, A2 => n118895, B1 => n120019, B2 
                           => OUT2_44_port, ZN => n116949);
   U86623 : AOI22_X1 port map( A1 => n119955, A2 => n118369, B1 => n119949, B2 
                           => n118249, ZN => n116956);
   U86624 : AOI22_X1 port map( A1 => n119979, A2 => n118956, B1 => n119973, B2 
                           => n118070, ZN => n116931);
   U86625 : AOI22_X1 port map( A1 => n120027, A2 => n118896, B1 => n120019, B2 
                           => OUT2_45_port, ZN => n116926);
   U86626 : AOI22_X1 port map( A1 => n119955, A2 => n118370, B1 => n119949, B2 
                           => n118250, ZN => n116933);
   U86627 : AOI22_X1 port map( A1 => n119979, A2 => n118957, B1 => n119973, B2 
                           => n118071, ZN => n116908);
   U86628 : AOI22_X1 port map( A1 => n120027, A2 => n118897, B1 => n120019, B2 
                           => OUT2_46_port, ZN => n116903);
   U86629 : AOI22_X1 port map( A1 => n119955, A2 => n118371, B1 => n119949, B2 
                           => n118251, ZN => n116910);
   U86630 : AOI22_X1 port map( A1 => n119979, A2 => n118958, B1 => n119973, B2 
                           => n118072, ZN => n116885);
   U86631 : AOI22_X1 port map( A1 => n120027, A2 => n118898, B1 => n120019, B2 
                           => OUT2_47_port, ZN => n116880);
   U86632 : AOI22_X1 port map( A1 => n119955, A2 => n118372, B1 => n119949, B2 
                           => n118252, ZN => n116887);
   U86633 : AOI22_X1 port map( A1 => n119980, A2 => n118959, B1 => n119974, B2 
                           => n118073, ZN => n116862);
   U86634 : AOI22_X1 port map( A1 => n120028, A2 => n118899, B1 => n120019, B2 
                           => OUT2_48_port, ZN => n116857);
   U86635 : AOI22_X1 port map( A1 => n119956, A2 => n118373, B1 => n119950, B2 
                           => n118253, ZN => n116864);
   U86636 : AOI22_X1 port map( A1 => n119980, A2 => n118960, B1 => n119974, B2 
                           => n118074, ZN => n116839);
   U86637 : AOI22_X1 port map( A1 => n120028, A2 => n118900, B1 => n120019, B2 
                           => OUT2_49_port, ZN => n116834);
   U86638 : AOI22_X1 port map( A1 => n119956, A2 => n118374, B1 => n119950, B2 
                           => n118254, ZN => n116841);
   U86639 : AOI22_X1 port map( A1 => n119980, A2 => n118961, B1 => n119974, B2 
                           => n118075, ZN => n116816);
   U86640 : AOI22_X1 port map( A1 => n120028, A2 => n118901, B1 => n120019, B2 
                           => OUT2_50_port, ZN => n116811);
   U86641 : AOI22_X1 port map( A1 => n119956, A2 => n118375, B1 => n119950, B2 
                           => n118255, ZN => n116818);
   U86642 : AOI22_X1 port map( A1 => n119980, A2 => n118962, B1 => n119974, B2 
                           => n118076, ZN => n116793);
   U86643 : AOI22_X1 port map( A1 => n120028, A2 => n118902, B1 => n120019, B2 
                           => OUT2_51_port, ZN => n116788);
   U86644 : AOI22_X1 port map( A1 => n119956, A2 => n118376, B1 => n119950, B2 
                           => n118256, ZN => n116795);
   U86645 : AOI22_X1 port map( A1 => n119980, A2 => n118963, B1 => n119974, B2 
                           => n118077, ZN => n116770);
   U86646 : AOI22_X1 port map( A1 => n120028, A2 => n118903, B1 => n120019, B2 
                           => OUT2_52_port, ZN => n116765);
   U86647 : AOI22_X1 port map( A1 => n119956, A2 => n118377, B1 => n119950, B2 
                           => n118257, ZN => n116772);
   U86648 : AOI22_X1 port map( A1 => n119980, A2 => n118964, B1 => n119974, B2 
                           => n118078, ZN => n116747);
   U86649 : AOI22_X1 port map( A1 => n120028, A2 => n118904, B1 => n120019, B2 
                           => OUT2_53_port, ZN => n116742);
   U86650 : AOI22_X1 port map( A1 => n119956, A2 => n118378, B1 => n119950, B2 
                           => n118258, ZN => n116749);
   U86651 : AOI22_X1 port map( A1 => n119980, A2 => n118965, B1 => n119974, B2 
                           => n118079, ZN => n116724);
   U86652 : AOI22_X1 port map( A1 => n120028, A2 => n118905, B1 => n120019, B2 
                           => OUT2_54_port, ZN => n116719);
   U86653 : AOI22_X1 port map( A1 => n119956, A2 => n118379, B1 => n119950, B2 
                           => n118259, ZN => n116726);
   U86654 : AOI22_X1 port map( A1 => n119980, A2 => n118966, B1 => n119974, B2 
                           => n118080, ZN => n116701);
   U86655 : AOI22_X1 port map( A1 => n120028, A2 => n118906, B1 => n120018, B2 
                           => OUT2_55_port, ZN => n116696);
   U86656 : AOI22_X1 port map( A1 => n119956, A2 => n118380, B1 => n119950, B2 
                           => n118260, ZN => n116703);
   U86657 : AOI22_X1 port map( A1 => n119980, A2 => n118967, B1 => n119974, B2 
                           => n118081, ZN => n116678);
   U86658 : AOI22_X1 port map( A1 => n120028, A2 => n118907, B1 => n120018, B2 
                           => OUT2_56_port, ZN => n116673);
   U86659 : AOI22_X1 port map( A1 => n119956, A2 => n118381, B1 => n119950, B2 
                           => n118261, ZN => n116680);
   U86660 : AOI22_X1 port map( A1 => n119980, A2 => n118968, B1 => n119974, B2 
                           => n118082, ZN => n116655);
   U86661 : AOI22_X1 port map( A1 => n120028, A2 => n118908, B1 => n120018, B2 
                           => OUT2_57_port, ZN => n116650);
   U86662 : AOI22_X1 port map( A1 => n119956, A2 => n118382, B1 => n119950, B2 
                           => n118262, ZN => n116657);
   U86663 : AOI22_X1 port map( A1 => n119980, A2 => n118969, B1 => n119974, B2 
                           => n118083, ZN => n116632);
   U86664 : AOI22_X1 port map( A1 => n120028, A2 => n118909, B1 => n120018, B2 
                           => OUT2_58_port, ZN => n116627);
   U86665 : AOI22_X1 port map( A1 => n119956, A2 => n118383, B1 => n119950, B2 
                           => n118263, ZN => n116634);
   U86666 : AOI22_X1 port map( A1 => n119980, A2 => n118970, B1 => n119974, B2 
                           => n118084, ZN => n116609);
   U86667 : AOI22_X1 port map( A1 => n120028, A2 => n118910, B1 => n120018, B2 
                           => OUT2_59_port, ZN => n116604);
   U86668 : AOI22_X1 port map( A1 => n119956, A2 => n118384, B1 => n119950, B2 
                           => n118264, ZN => n116611);
   U86669 : AOI22_X1 port map( A1 => n120225, A2 => n118532, B1 => n120217, B2 
                           => OUT1_46_port, ZN => n115155);
   U86670 : AOI22_X1 port map( A1 => n120177, A2 => n118251, B1 => n120171, B2 
                           => n119114, ZN => n115160);
   U86671 : AOI22_X1 port map( A1 => n120153, A2 => n118738, B1 => n120147, B2 
                           => n119050, ZN => n115162);
   U86672 : AOI22_X1 port map( A1 => n120225, A2 => n118533, B1 => n120217, B2 
                           => OUT1_47_port, ZN => n115127);
   U86673 : AOI22_X1 port map( A1 => n120177, A2 => n118252, B1 => n120171, B2 
                           => n119115, ZN => n115132);
   U86674 : AOI22_X1 port map( A1 => n120153, A2 => n118739, B1 => n120147, B2 
                           => n119051, ZN => n115134);
   U86675 : AOI22_X1 port map( A1 => n120226, A2 => n118534, B1 => n120217, B2 
                           => OUT1_48_port, ZN => n115099);
   U86676 : AOI22_X1 port map( A1 => n120178, A2 => n118253, B1 => n120172, B2 
                           => n119116, ZN => n115104);
   U86677 : AOI22_X1 port map( A1 => n120154, A2 => n118740, B1 => n120148, B2 
                           => n119052, ZN => n115106);
   U86678 : AOI22_X1 port map( A1 => n120226, A2 => n118535, B1 => n120217, B2 
                           => OUT1_49_port, ZN => n115071);
   U86679 : AOI22_X1 port map( A1 => n120178, A2 => n118254, B1 => n120172, B2 
                           => n119117, ZN => n115076);
   U86680 : AOI22_X1 port map( A1 => n120154, A2 => n118741, B1 => n120148, B2 
                           => n119053, ZN => n115078);
   U86681 : AOI22_X1 port map( A1 => n120226, A2 => n118536, B1 => n120217, B2 
                           => OUT1_50_port, ZN => n115043);
   U86682 : AOI22_X1 port map( A1 => n120178, A2 => n118255, B1 => n120172, B2 
                           => n119118, ZN => n115048);
   U86683 : AOI22_X1 port map( A1 => n120154, A2 => n118742, B1 => n120148, B2 
                           => n119054, ZN => n115050);
   U86684 : AOI22_X1 port map( A1 => n120226, A2 => n118537, B1 => n120217, B2 
                           => OUT1_51_port, ZN => n115015);
   U86685 : AOI22_X1 port map( A1 => n120178, A2 => n118256, B1 => n120172, B2 
                           => n119119, ZN => n115020);
   U86686 : AOI22_X1 port map( A1 => n120154, A2 => n118743, B1 => n120148, B2 
                           => n119055, ZN => n115022);
   U86687 : AOI22_X1 port map( A1 => n120226, A2 => n118538, B1 => n120217, B2 
                           => OUT1_52_port, ZN => n114987);
   U86688 : AOI22_X1 port map( A1 => n120178, A2 => n118257, B1 => n120172, B2 
                           => n119120, ZN => n114992);
   U86689 : AOI22_X1 port map( A1 => n120154, A2 => n118744, B1 => n120148, B2 
                           => n119056, ZN => n114994);
   U86690 : AOI22_X1 port map( A1 => n120226, A2 => n118539, B1 => n120217, B2 
                           => OUT1_53_port, ZN => n114959);
   U86691 : AOI22_X1 port map( A1 => n120178, A2 => n118258, B1 => n120172, B2 
                           => n119121, ZN => n114964);
   U86692 : AOI22_X1 port map( A1 => n120154, A2 => n118745, B1 => n120148, B2 
                           => n119057, ZN => n114966);
   U86693 : AOI22_X1 port map( A1 => n120226, A2 => n118540, B1 => n120217, B2 
                           => OUT1_54_port, ZN => n114931);
   U86694 : AOI22_X1 port map( A1 => n120178, A2 => n118259, B1 => n120172, B2 
                           => n119122, ZN => n114936);
   U86695 : AOI22_X1 port map( A1 => n120154, A2 => n118746, B1 => n120148, B2 
                           => n119058, ZN => n114938);
   U86696 : AOI22_X1 port map( A1 => n120226, A2 => n118541, B1 => n120216, B2 
                           => OUT1_55_port, ZN => n114903);
   U86697 : AOI22_X1 port map( A1 => n120178, A2 => n118260, B1 => n120172, B2 
                           => n119123, ZN => n114908);
   U86698 : AOI22_X1 port map( A1 => n120154, A2 => n118747, B1 => n120148, B2 
                           => n119059, ZN => n114910);
   U86699 : AOI22_X1 port map( A1 => n120226, A2 => n118542, B1 => n120216, B2 
                           => OUT1_56_port, ZN => n114875);
   U86700 : AOI22_X1 port map( A1 => n120178, A2 => n118261, B1 => n120172, B2 
                           => n119124, ZN => n114880);
   U86701 : AOI22_X1 port map( A1 => n120154, A2 => n118748, B1 => n120148, B2 
                           => n119060, ZN => n114882);
   U86702 : AOI22_X1 port map( A1 => n120226, A2 => n118543, B1 => n120216, B2 
                           => OUT1_57_port, ZN => n114847);
   U86703 : AOI22_X1 port map( A1 => n120178, A2 => n118262, B1 => n120172, B2 
                           => n119125, ZN => n114852);
   U86704 : AOI22_X1 port map( A1 => n120154, A2 => n118749, B1 => n120148, B2 
                           => n119061, ZN => n114854);
   U86705 : AOI22_X1 port map( A1 => n120226, A2 => n118544, B1 => n120216, B2 
                           => OUT1_58_port, ZN => n114819);
   U86706 : AOI22_X1 port map( A1 => n120178, A2 => n118263, B1 => n120172, B2 
                           => n119126, ZN => n114824);
   U86707 : AOI22_X1 port map( A1 => n120154, A2 => n118750, B1 => n120148, B2 
                           => n119062, ZN => n114826);
   U86708 : AOI22_X1 port map( A1 => n120226, A2 => n118545, B1 => n120216, B2 
                           => OUT1_59_port, ZN => n114791);
   U86709 : AOI22_X1 port map( A1 => n120178, A2 => n118264, B1 => n120172, B2 
                           => n119127, ZN => n114796);
   U86710 : AOI22_X1 port map( A1 => n120154, A2 => n118751, B1 => n120148, B2 
                           => n119063, ZN => n114798);
   U86711 : AOI22_X1 port map( A1 => n120222, A2 => n118810, B1 => n120216, B2 
                           => OUT1_0_port, ZN => n116443);
   U86712 : AOI22_X1 port map( A1 => n120174, A2 => n118205, B1 => n120168, B2 
                           => n119128, ZN => n116455);
   U86713 : AOI22_X1 port map( A1 => n120150, A2 => n118752, B1 => n120144, B2 
                           => n119064, ZN => n116460);
   U86714 : AOI22_X1 port map( A1 => n120222, A2 => n118811, B1 => n120221, B2 
                           => OUT1_1_port, ZN => n116415);
   U86715 : AOI22_X1 port map( A1 => n120174, A2 => n118206, B1 => n120168, B2 
                           => n119129, ZN => n116420);
   U86716 : AOI22_X1 port map( A1 => n120150, A2 => n118753, B1 => n120144, B2 
                           => n119065, ZN => n116422);
   U86717 : AOI22_X1 port map( A1 => n120222, A2 => n118812, B1 => n120221, B2 
                           => OUT1_2_port, ZN => n116387);
   U86718 : AOI22_X1 port map( A1 => n120174, A2 => n118207, B1 => n120168, B2 
                           => n119130, ZN => n116392);
   U86719 : AOI22_X1 port map( A1 => n120150, A2 => n118754, B1 => n120144, B2 
                           => n119066, ZN => n116394);
   U86720 : AOI22_X1 port map( A1 => n120222, A2 => n118813, B1 => n120221, B2 
                           => OUT1_3_port, ZN => n116359);
   U86721 : AOI22_X1 port map( A1 => n120174, A2 => n118208, B1 => n120168, B2 
                           => n119131, ZN => n116364);
   U86722 : AOI22_X1 port map( A1 => n120150, A2 => n118755, B1 => n120144, B2 
                           => n119067, ZN => n116366);
   U86723 : AOI22_X1 port map( A1 => n119976, A2 => n118971, B1 => n119970, B2 
                           => n111003, ZN => n117794);
   U86724 : AOI22_X1 port map( A1 => n120024, A2 => n118911, B1 => n120022, B2 
                           => OUT2_7_port, ZN => n117789);
   U86725 : AOI22_X1 port map( A1 => n119952, A2 => n118332, B1 => n119946, B2 
                           => n118212, ZN => n117796);
   U86726 : AOI22_X1 port map( A1 => n119976, A2 => n118972, B1 => n119970, B2 
                           => n111004, ZN => n117772);
   U86727 : AOI22_X1 port map( A1 => n120024, A2 => n118912, B1 => n120022, B2 
                           => OUT2_8_port, ZN => n117767);
   U86728 : AOI22_X1 port map( A1 => n119952, A2 => n118333, B1 => n119946, B2 
                           => n118213, ZN => n117774);
   U86729 : AOI22_X1 port map( A1 => n119976, A2 => n118973, B1 => n119970, B2 
                           => n111005, ZN => n117750);
   U86730 : AOI22_X1 port map( A1 => n120024, A2 => n118913, B1 => n120022, B2 
                           => OUT2_9_port, ZN => n117745);
   U86731 : AOI22_X1 port map( A1 => n119952, A2 => n118334, B1 => n119946, B2 
                           => n118214, ZN => n117752);
   U86732 : AOI22_X1 port map( A1 => n119976, A2 => n118974, B1 => n119970, B2 
                           => n111006, ZN => n117728);
   U86733 : AOI22_X1 port map( A1 => n120024, A2 => n118914, B1 => n120022, B2 
                           => OUT2_10_port, ZN => n117723);
   U86734 : AOI22_X1 port map( A1 => n119952, A2 => n118335, B1 => n119946, B2 
                           => n118215, ZN => n117730);
   U86735 : AOI22_X1 port map( A1 => n119976, A2 => n118975, B1 => n119970, B2 
                           => n110996, ZN => n117956);
   U86736 : AOI22_X1 port map( A1 => n120024, A2 => n118915, B1 => n120018, B2 
                           => OUT2_0_port, ZN => n117943);
   U86737 : AOI22_X1 port map( A1 => n119952, A2 => n118325, B1 => n119946, B2 
                           => n118205, ZN => n117960);
   U86738 : AOI22_X1 port map( A1 => n119976, A2 => n118976, B1 => n119970, B2 
                           => n110997, ZN => n117926);
   U86739 : AOI22_X1 port map( A1 => n120024, A2 => n118916, B1 => n120023, B2 
                           => OUT2_1_port, ZN => n117921);
   U86740 : AOI22_X1 port map( A1 => n119952, A2 => n118326, B1 => n119946, B2 
                           => n118206, ZN => n117928);
   U86741 : AOI22_X1 port map( A1 => n119976, A2 => n118977, B1 => n119970, B2 
                           => n110998, ZN => n117904);
   U86742 : AOI22_X1 port map( A1 => n120024, A2 => n118917, B1 => n120023, B2 
                           => OUT2_2_port, ZN => n117899);
   U86743 : AOI22_X1 port map( A1 => n119952, A2 => n118327, B1 => n119946, B2 
                           => n118207, ZN => n117906);
   U86744 : AOI22_X1 port map( A1 => n119976, A2 => n118978, B1 => n119970, B2 
                           => n110999, ZN => n117882);
   U86745 : AOI22_X1 port map( A1 => n120024, A2 => n118918, B1 => n120023, B2 
                           => OUT2_3_port, ZN => n117877);
   U86746 : AOI22_X1 port map( A1 => n119952, A2 => n118328, B1 => n119946, B2 
                           => n118208, ZN => n117884);
   U86747 : AOI22_X1 port map( A1 => n119976, A2 => n118979, B1 => n119970, B2 
                           => n111000, ZN => n117860);
   U86748 : AOI22_X1 port map( A1 => n120024, A2 => n118919, B1 => n120022, B2 
                           => OUT2_4_port, ZN => n117855);
   U86749 : AOI22_X1 port map( A1 => n119952, A2 => n118329, B1 => n119946, B2 
                           => n118209, ZN => n117862);
   U86750 : AOI22_X1 port map( A1 => n119976, A2 => n118980, B1 => n119970, B2 
                           => n111001, ZN => n117838);
   U86751 : AOI22_X1 port map( A1 => n120024, A2 => n118920, B1 => n120022, B2 
                           => OUT2_5_port, ZN => n117833);
   U86752 : AOI22_X1 port map( A1 => n119952, A2 => n118330, B1 => n119946, B2 
                           => n118210, ZN => n117840);
   U86753 : AOI22_X1 port map( A1 => n119976, A2 => n118981, B1 => n119970, B2 
                           => n111002, ZN => n117816);
   U86754 : AOI22_X1 port map( A1 => n120024, A2 => n118921, B1 => n120022, B2 
                           => OUT2_6_port, ZN => n117811);
   U86755 : AOI22_X1 port map( A1 => n119952, A2 => n118331, B1 => n119946, B2 
                           => n118211, ZN => n117818);
   U86756 : AOI22_X1 port map( A1 => n120222, A2 => n118814, B1 => n120220, B2 
                           => OUT1_4_port, ZN => n116331);
   U86757 : AOI22_X1 port map( A1 => n120174, A2 => n118209, B1 => n120168, B2 
                           => n119132, ZN => n116336);
   U86758 : AOI22_X1 port map( A1 => n120150, A2 => n118756, B1 => n120144, B2 
                           => n119068, ZN => n116338);
   U86759 : AOI22_X1 port map( A1 => n120222, A2 => n118815, B1 => n120220, B2 
                           => OUT1_5_port, ZN => n116303);
   U86760 : AOI22_X1 port map( A1 => n120174, A2 => n118210, B1 => n120168, B2 
                           => n119133, ZN => n116308);
   U86761 : AOI22_X1 port map( A1 => n120150, A2 => n118757, B1 => n120144, B2 
                           => n119069, ZN => n116310);
   U86762 : AOI22_X1 port map( A1 => n120222, A2 => n118816, B1 => n120220, B2 
                           => OUT1_6_port, ZN => n116275);
   U86763 : AOI22_X1 port map( A1 => n120174, A2 => n118211, B1 => n120168, B2 
                           => n119134, ZN => n116280);
   U86764 : AOI22_X1 port map( A1 => n120150, A2 => n118758, B1 => n120144, B2 
                           => n119070, ZN => n116282);
   U86765 : AOI22_X1 port map( A1 => n120222, A2 => n118806, B1 => n120220, B2 
                           => OUT1_7_port, ZN => n116247);
   U86766 : AOI22_X1 port map( A1 => n120174, A2 => n118212, B1 => n120168, B2 
                           => n119135, ZN => n116252);
   U86767 : AOI22_X1 port map( A1 => n120150, A2 => n118759, B1 => n120144, B2 
                           => n119071, ZN => n116254);
   U86768 : AOI22_X1 port map( A1 => n120222, A2 => n118807, B1 => n120220, B2 
                           => OUT1_8_port, ZN => n116219);
   U86769 : AOI22_X1 port map( A1 => n120174, A2 => n118213, B1 => n120168, B2 
                           => n119136, ZN => n116224);
   U86770 : AOI22_X1 port map( A1 => n120150, A2 => n118760, B1 => n120144, B2 
                           => n119072, ZN => n116226);
   U86771 : AOI22_X1 port map( A1 => n120222, A2 => n118808, B1 => n120220, B2 
                           => OUT1_9_port, ZN => n116191);
   U86772 : AOI22_X1 port map( A1 => n120174, A2 => n118214, B1 => n120168, B2 
                           => n119137, ZN => n116196);
   U86773 : AOI22_X1 port map( A1 => n120150, A2 => n118761, B1 => n120144, B2 
                           => n119073, ZN => n116198);
   U86774 : AOI22_X1 port map( A1 => n120222, A2 => n118809, B1 => n120220, B2 
                           => OUT1_10_port, ZN => n116163);
   U86775 : AOI22_X1 port map( A1 => n120174, A2 => n118215, B1 => n120168, B2 
                           => n119138, ZN => n116168);
   U86776 : AOI22_X1 port map( A1 => n120150, A2 => n118762, B1 => n120144, B2 
                           => n119074, ZN => n116170);
   U86777 : AOI22_X1 port map( A1 => n120222, A2 => n118798, B1 => n120220, B2 
                           => OUT1_11_port, ZN => n116135);
   U86778 : AOI22_X1 port map( A1 => n120174, A2 => n118216, B1 => n120168, B2 
                           => n119139, ZN => n116140);
   U86779 : AOI22_X1 port map( A1 => n120150, A2 => n118763, B1 => n120144, B2 
                           => n119075, ZN => n116142);
   U86780 : AOI22_X1 port map( A1 => n120223, A2 => n118799, B1 => n120220, B2 
                           => OUT1_12_port, ZN => n116107);
   U86781 : AOI22_X1 port map( A1 => n120175, A2 => n118217, B1 => n120169, B2 
                           => n119140, ZN => n116112);
   U86782 : AOI22_X1 port map( A1 => n120151, A2 => n118764, B1 => n120145, B2 
                           => n119076, ZN => n116114);
   U86783 : AOI22_X1 port map( A1 => n120223, A2 => n118800, B1 => n120220, B2 
                           => OUT1_13_port, ZN => n116079);
   U86784 : AOI22_X1 port map( A1 => n120175, A2 => n118218, B1 => n120169, B2 
                           => n119141, ZN => n116084);
   U86785 : AOI22_X1 port map( A1 => n120151, A2 => n118765, B1 => n120145, B2 
                           => n119077, ZN => n116086);
   U86786 : AOI22_X1 port map( A1 => n120223, A2 => n118801, B1 => n120220, B2 
                           => OUT1_14_port, ZN => n116051);
   U86787 : AOI22_X1 port map( A1 => n120175, A2 => n118219, B1 => n120169, B2 
                           => n119142, ZN => n116056);
   U86788 : AOI22_X1 port map( A1 => n120151, A2 => n118766, B1 => n120145, B2 
                           => n119078, ZN => n116058);
   U86789 : AOI22_X1 port map( A1 => n120223, A2 => n118802, B1 => n120220, B2 
                           => OUT1_15_port, ZN => n116023);
   U86790 : AOI22_X1 port map( A1 => n120175, A2 => n118220, B1 => n120169, B2 
                           => n119143, ZN => n116028);
   U86791 : AOI22_X1 port map( A1 => n120151, A2 => n118767, B1 => n120145, B2 
                           => n119079, ZN => n116030);
   U86792 : AOI22_X1 port map( A1 => n120223, A2 => n118803, B1 => n120220, B2 
                           => OUT1_16_port, ZN => n115995);
   U86793 : AOI22_X1 port map( A1 => n120175, A2 => n118221, B1 => n120169, B2 
                           => n119144, ZN => n116000);
   U86794 : AOI22_X1 port map( A1 => n120151, A2 => n118768, B1 => n120145, B2 
                           => n119080, ZN => n116002);
   U86795 : AOI22_X1 port map( A1 => n120223, A2 => n118804, B1 => n120219, B2 
                           => OUT1_17_port, ZN => n115967);
   U86796 : AOI22_X1 port map( A1 => n120175, A2 => n118222, B1 => n120169, B2 
                           => n119145, ZN => n115972);
   U86797 : AOI22_X1 port map( A1 => n120151, A2 => n118769, B1 => n120145, B2 
                           => n119081, ZN => n115974);
   U86798 : AOI22_X1 port map( A1 => n120223, A2 => n118805, B1 => n120219, B2 
                           => OUT1_18_port, ZN => n115939);
   U86799 : AOI22_X1 port map( A1 => n120175, A2 => n118223, B1 => n120169, B2 
                           => n119146, ZN => n115944);
   U86800 : AOI22_X1 port map( A1 => n120151, A2 => n118770, B1 => n120145, B2 
                           => n119082, ZN => n115946);
   U86801 : AOI22_X1 port map( A1 => n120223, A2 => n118505, B1 => n120219, B2 
                           => OUT1_19_port, ZN => n115911);
   U86802 : AOI22_X1 port map( A1 => n120175, A2 => n118224, B1 => n120169, B2 
                           => n119147, ZN => n115916);
   U86803 : AOI22_X1 port map( A1 => n120151, A2 => n118771, B1 => n120145, B2 
                           => n119083, ZN => n115918);
   U86804 : AOI22_X1 port map( A1 => n120223, A2 => n118506, B1 => n120219, B2 
                           => OUT1_20_port, ZN => n115883);
   U86805 : AOI22_X1 port map( A1 => n120175, A2 => n118225, B1 => n120169, B2 
                           => n119148, ZN => n115888);
   U86806 : AOI22_X1 port map( A1 => n120151, A2 => n118772, B1 => n120145, B2 
                           => n119084, ZN => n115890);
   U86807 : AOI22_X1 port map( A1 => n120223, A2 => n118507, B1 => n120219, B2 
                           => OUT1_21_port, ZN => n115855);
   U86808 : AOI22_X1 port map( A1 => n120175, A2 => n118226, B1 => n120169, B2 
                           => n119149, ZN => n115860);
   U86809 : AOI22_X1 port map( A1 => n120151, A2 => n118773, B1 => n120145, B2 
                           => n119085, ZN => n115862);
   U86810 : AOI22_X1 port map( A1 => n120223, A2 => n118508, B1 => n120219, B2 
                           => OUT1_22_port, ZN => n115827);
   U86811 : AOI22_X1 port map( A1 => n120175, A2 => n118227, B1 => n120169, B2 
                           => n119150, ZN => n115832);
   U86812 : AOI22_X1 port map( A1 => n120151, A2 => n118774, B1 => n120145, B2 
                           => n119086, ZN => n115834);
   U86813 : AOI22_X1 port map( A1 => n120223, A2 => n118509, B1 => n120219, B2 
                           => OUT1_23_port, ZN => n115799);
   U86814 : AOI22_X1 port map( A1 => n120175, A2 => n118228, B1 => n120169, B2 
                           => n119151, ZN => n115804);
   U86815 : AOI22_X1 port map( A1 => n120151, A2 => n118775, B1 => n120145, B2 
                           => n119087, ZN => n115806);
   U86816 : AOI22_X1 port map( A1 => n120224, A2 => n118510, B1 => n120219, B2 
                           => OUT1_24_port, ZN => n115771);
   U86817 : AOI22_X1 port map( A1 => n120176, A2 => n118229, B1 => n120170, B2 
                           => n119152, ZN => n115776);
   U86818 : AOI22_X1 port map( A1 => n120152, A2 => n118776, B1 => n120146, B2 
                           => n119088, ZN => n115778);
   U86819 : AOI22_X1 port map( A1 => n120224, A2 => n118511, B1 => n120219, B2 
                           => OUT1_25_port, ZN => n115743);
   U86820 : AOI22_X1 port map( A1 => n120176, A2 => n118230, B1 => n120170, B2 
                           => n119153, ZN => n115748);
   U86821 : AOI22_X1 port map( A1 => n120152, A2 => n118777, B1 => n120146, B2 
                           => n119089, ZN => n115750);
   U86822 : AOI22_X1 port map( A1 => n120224, A2 => n118512, B1 => n120219, B2 
                           => OUT1_26_port, ZN => n115715);
   U86823 : AOI22_X1 port map( A1 => n120176, A2 => n118231, B1 => n120170, B2 
                           => n119154, ZN => n115720);
   U86824 : AOI22_X1 port map( A1 => n120152, A2 => n118778, B1 => n120146, B2 
                           => n119090, ZN => n115722);
   U86825 : AOI22_X1 port map( A1 => n120224, A2 => n118513, B1 => n120219, B2 
                           => OUT1_27_port, ZN => n115687);
   U86826 : AOI22_X1 port map( A1 => n120176, A2 => n118232, B1 => n120170, B2 
                           => n119155, ZN => n115692);
   U86827 : AOI22_X1 port map( A1 => n120152, A2 => n118779, B1 => n120146, B2 
                           => n119091, ZN => n115694);
   U86828 : AOI22_X1 port map( A1 => n120224, A2 => n118514, B1 => n120219, B2 
                           => OUT1_28_port, ZN => n115659);
   U86829 : AOI22_X1 port map( A1 => n120176, A2 => n118233, B1 => n120170, B2 
                           => n119156, ZN => n115664);
   U86830 : AOI22_X1 port map( A1 => n120152, A2 => n118780, B1 => n120146, B2 
                           => n119092, ZN => n115666);
   U86831 : AOI22_X1 port map( A1 => n120224, A2 => n118515, B1 => n120219, B2 
                           => OUT1_29_port, ZN => n115631);
   U86832 : AOI22_X1 port map( A1 => n120176, A2 => n118234, B1 => n120170, B2 
                           => n119157, ZN => n115636);
   U86833 : AOI22_X1 port map( A1 => n120152, A2 => n118781, B1 => n120146, B2 
                           => n119093, ZN => n115638);
   U86834 : AOI22_X1 port map( A1 => n120224, A2 => n118516, B1 => n120218, B2 
                           => OUT1_30_port, ZN => n115603);
   U86835 : AOI22_X1 port map( A1 => n120176, A2 => n118235, B1 => n120170, B2 
                           => n119158, ZN => n115608);
   U86836 : AOI22_X1 port map( A1 => n120152, A2 => n118782, B1 => n120146, B2 
                           => n119094, ZN => n115610);
   U86837 : AOI22_X1 port map( A1 => n120224, A2 => n118517, B1 => n120218, B2 
                           => OUT1_31_port, ZN => n115575);
   U86838 : AOI22_X1 port map( A1 => n120176, A2 => n118236, B1 => n120170, B2 
                           => n119159, ZN => n115580);
   U86839 : AOI22_X1 port map( A1 => n120152, A2 => n118783, B1 => n120146, B2 
                           => n119095, ZN => n115582);
   U86840 : AOI22_X1 port map( A1 => n120224, A2 => n118518, B1 => n120218, B2 
                           => OUT1_32_port, ZN => n115547);
   U86841 : AOI22_X1 port map( A1 => n120176, A2 => n118237, B1 => n120170, B2 
                           => n119160, ZN => n115552);
   U86842 : AOI22_X1 port map( A1 => n120152, A2 => n118784, B1 => n120146, B2 
                           => n119096, ZN => n115554);
   U86843 : AOI22_X1 port map( A1 => n120224, A2 => n118519, B1 => n120218, B2 
                           => OUT1_33_port, ZN => n115519);
   U86844 : AOI22_X1 port map( A1 => n120176, A2 => n118238, B1 => n120170, B2 
                           => n119161, ZN => n115524);
   U86845 : AOI22_X1 port map( A1 => n120152, A2 => n118785, B1 => n120146, B2 
                           => n119097, ZN => n115526);
   U86846 : AOI22_X1 port map( A1 => n120224, A2 => n118520, B1 => n120218, B2 
                           => OUT1_34_port, ZN => n115491);
   U86847 : AOI22_X1 port map( A1 => n120176, A2 => n118239, B1 => n120170, B2 
                           => n119162, ZN => n115496);
   U86848 : AOI22_X1 port map( A1 => n120152, A2 => n118786, B1 => n120146, B2 
                           => n119098, ZN => n115498);
   U86849 : AOI22_X1 port map( A1 => n120224, A2 => n118521, B1 => n120218, B2 
                           => OUT1_35_port, ZN => n115463);
   U86850 : AOI22_X1 port map( A1 => n120176, A2 => n118240, B1 => n120170, B2 
                           => n119163, ZN => n115468);
   U86851 : AOI22_X1 port map( A1 => n120152, A2 => n118787, B1 => n120146, B2 
                           => n119099, ZN => n115470);
   U86852 : AOI22_X1 port map( A1 => n120225, A2 => n118522, B1 => n120218, B2 
                           => OUT1_36_port, ZN => n115435);
   U86853 : AOI22_X1 port map( A1 => n120177, A2 => n118241, B1 => n120171, B2 
                           => n119164, ZN => n115440);
   U86854 : AOI22_X1 port map( A1 => n120153, A2 => n118788, B1 => n120147, B2 
                           => n119100, ZN => n115442);
   U86855 : AOI22_X1 port map( A1 => n120225, A2 => n118523, B1 => n120218, B2 
                           => OUT1_37_port, ZN => n115407);
   U86856 : AOI22_X1 port map( A1 => n120177, A2 => n118242, B1 => n120171, B2 
                           => n119165, ZN => n115412);
   U86857 : AOI22_X1 port map( A1 => n120153, A2 => n118789, B1 => n120147, B2 
                           => n119101, ZN => n115414);
   U86858 : AOI22_X1 port map( A1 => n120225, A2 => n118524, B1 => n120218, B2 
                           => OUT1_38_port, ZN => n115379);
   U86859 : AOI22_X1 port map( A1 => n120177, A2 => n118243, B1 => n120171, B2 
                           => n119166, ZN => n115384);
   U86860 : AOI22_X1 port map( A1 => n120153, A2 => n118790, B1 => n120147, B2 
                           => n119102, ZN => n115386);
   U86861 : AOI22_X1 port map( A1 => n120225, A2 => n118525, B1 => n120218, B2 
                           => OUT1_39_port, ZN => n115351);
   U86862 : AOI22_X1 port map( A1 => n120177, A2 => n118244, B1 => n120171, B2 
                           => n119167, ZN => n115356);
   U86863 : AOI22_X1 port map( A1 => n120153, A2 => n118791, B1 => n120147, B2 
                           => n119103, ZN => n115358);
   U86864 : AOI22_X1 port map( A1 => n120225, A2 => n118526, B1 => n120218, B2 
                           => OUT1_40_port, ZN => n115323);
   U86865 : AOI22_X1 port map( A1 => n120177, A2 => n118245, B1 => n120171, B2 
                           => n119168, ZN => n115328);
   U86866 : AOI22_X1 port map( A1 => n120153, A2 => n118792, B1 => n120147, B2 
                           => n119104, ZN => n115330);
   U86867 : AOI22_X1 port map( A1 => n120225, A2 => n118527, B1 => n120218, B2 
                           => OUT1_41_port, ZN => n115295);
   U86868 : AOI22_X1 port map( A1 => n120177, A2 => n118246, B1 => n120171, B2 
                           => n119169, ZN => n115300);
   U86869 : AOI22_X1 port map( A1 => n120153, A2 => n118793, B1 => n120147, B2 
                           => n119105, ZN => n115302);
   U86870 : AOI22_X1 port map( A1 => n120225, A2 => n118528, B1 => n120217, B2 
                           => OUT1_42_port, ZN => n115267);
   U86871 : AOI22_X1 port map( A1 => n120177, A2 => n118247, B1 => n120171, B2 
                           => n119170, ZN => n115272);
   U86872 : AOI22_X1 port map( A1 => n120153, A2 => n118794, B1 => n120147, B2 
                           => n119106, ZN => n115274);
   U86873 : AOI22_X1 port map( A1 => n120225, A2 => n118529, B1 => n120217, B2 
                           => OUT1_43_port, ZN => n115239);
   U86874 : AOI22_X1 port map( A1 => n120177, A2 => n118248, B1 => n120171, B2 
                           => n119171, ZN => n115244);
   U86875 : AOI22_X1 port map( A1 => n120153, A2 => n118795, B1 => n120147, B2 
                           => n119107, ZN => n115246);
   U86876 : AOI22_X1 port map( A1 => n120225, A2 => n118530, B1 => n120217, B2 
                           => OUT1_44_port, ZN => n115211);
   U86877 : AOI22_X1 port map( A1 => n120177, A2 => n118249, B1 => n120171, B2 
                           => n119172, ZN => n115216);
   U86878 : AOI22_X1 port map( A1 => n120153, A2 => n118796, B1 => n120147, B2 
                           => n119108, ZN => n115218);
   U86879 : AOI22_X1 port map( A1 => n120225, A2 => n118531, B1 => n120217, B2 
                           => OUT1_45_port, ZN => n115183);
   U86880 : AOI22_X1 port map( A1 => n120177, A2 => n118250, B1 => n120171, B2 
                           => n119173, ZN => n115188);
   U86881 : AOI22_X1 port map( A1 => n120153, A2 => n118797, B1 => n120147, B2 
                           => n119109, ZN => n115190);
   U86882 : OAI221_X1 port map( B1 => n99967, B2 => n120012, C1 => n114431, C2 
                           => n120006, A => n117703, ZN => n117699);
   U86883 : AOI22_X1 port map( A1 => n120000, A2 => n118670, B1 => n119994, B2 
                           => n119302, ZN => n117703);
   U86884 : OAI221_X1 port map( B1 => n99966, B2 => n120013, C1 => n114430, C2 
                           => n120007, A => n117681, ZN => n117677);
   U86885 : AOI22_X1 port map( A1 => n120001, A2 => n118671, B1 => n119995, B2 
                           => n119303, ZN => n117681);
   U86886 : OAI221_X1 port map( B1 => n99965, B2 => n120013, C1 => n114429, C2 
                           => n120007, A => n117659, ZN => n117655);
   U86887 : AOI22_X1 port map( A1 => n120001, A2 => n118672, B1 => n119995, B2 
                           => n119304, ZN => n117659);
   U86888 : OAI221_X1 port map( B1 => n99964, B2 => n120013, C1 => n114428, C2 
                           => n120007, A => n117637, ZN => n117633);
   U86889 : AOI22_X1 port map( A1 => n120001, A2 => n118673, B1 => n119995, B2 
                           => n119305, ZN => n117637);
   U86890 : OAI221_X1 port map( B1 => n99963, B2 => n120013, C1 => n114427, C2 
                           => n120007, A => n117615, ZN => n117611);
   U86891 : AOI22_X1 port map( A1 => n120001, A2 => n118674, B1 => n119995, B2 
                           => n119306, ZN => n117615);
   U86892 : OAI221_X1 port map( B1 => n99962, B2 => n120013, C1 => n114426, C2 
                           => n120007, A => n117593, ZN => n117589);
   U86893 : AOI22_X1 port map( A1 => n120001, A2 => n118675, B1 => n119995, B2 
                           => n119307, ZN => n117593);
   U86894 : OAI221_X1 port map( B1 => n99961, B2 => n120013, C1 => n114425, C2 
                           => n120007, A => n117571, ZN => n117567);
   U86895 : AOI22_X1 port map( A1 => n120001, A2 => n118676, B1 => n119995, B2 
                           => n119308, ZN => n117571);
   U86896 : OAI221_X1 port map( B1 => n99960, B2 => n120013, C1 => n114424, C2 
                           => n120007, A => n117549, ZN => n117545);
   U86897 : AOI22_X1 port map( A1 => n120001, A2 => n118677, B1 => n119995, B2 
                           => n119309, ZN => n117549);
   U86898 : OAI221_X1 port map( B1 => n99959, B2 => n120013, C1 => n114423, C2 
                           => n120007, A => n117526, ZN => n117522);
   U86899 : AOI22_X1 port map( A1 => n120001, A2 => n118678, B1 => n119995, B2 
                           => n119310, ZN => n117526);
   U86900 : OAI221_X1 port map( B1 => n99958, B2 => n120013, C1 => n114422, C2 
                           => n120007, A => n117503, ZN => n117499);
   U86901 : AOI22_X1 port map( A1 => n120001, A2 => n118679, B1 => n119995, B2 
                           => n119311, ZN => n117503);
   U86902 : OAI221_X1 port map( B1 => n99957, B2 => n120013, C1 => n114421, C2 
                           => n120007, A => n117480, ZN => n117476);
   U86903 : AOI22_X1 port map( A1 => n120001, A2 => n118680, B1 => n119995, B2 
                           => n119312, ZN => n117480);
   U86904 : OAI221_X1 port map( B1 => n99956, B2 => n120013, C1 => n114420, C2 
                           => n120007, A => n117457, ZN => n117453);
   U86905 : AOI22_X1 port map( A1 => n120001, A2 => n118681, B1 => n119995, B2 
                           => n119313, ZN => n117457);
   U86906 : OAI221_X1 port map( B1 => n99955, B2 => n120013, C1 => n114419, C2 
                           => n120007, A => n117434, ZN => n117430);
   U86907 : AOI22_X1 port map( A1 => n120001, A2 => n118682, B1 => n119995, B2 
                           => n119314, ZN => n117434);
   U86908 : OAI221_X1 port map( B1 => n99954, B2 => n120014, C1 => n114418, C2 
                           => n120008, A => n117411, ZN => n117407);
   U86909 : AOI22_X1 port map( A1 => n120002, A2 => n118683, B1 => n119996, B2 
                           => n119315, ZN => n117411);
   U86910 : OAI221_X1 port map( B1 => n99953, B2 => n120014, C1 => n114417, C2 
                           => n120008, A => n117388, ZN => n117384);
   U86911 : AOI22_X1 port map( A1 => n120002, A2 => n118684, B1 => n119996, B2 
                           => n119316, ZN => n117388);
   U86912 : OAI221_X1 port map( B1 => n99952, B2 => n120014, C1 => n114416, C2 
                           => n120008, A => n117365, ZN => n117361);
   U86913 : AOI22_X1 port map( A1 => n120002, A2 => n118685, B1 => n119996, B2 
                           => n119317, ZN => n117365);
   U86914 : OAI221_X1 port map( B1 => n99951, B2 => n120014, C1 => n114415, C2 
                           => n120008, A => n117342, ZN => n117338);
   U86915 : AOI22_X1 port map( A1 => n120002, A2 => n118686, B1 => n119996, B2 
                           => n119318, ZN => n117342);
   U86916 : OAI221_X1 port map( B1 => n99950, B2 => n120014, C1 => n114414, C2 
                           => n120008, A => n117319, ZN => n117315);
   U86917 : AOI22_X1 port map( A1 => n120002, A2 => n118687, B1 => n119996, B2 
                           => n119319, ZN => n117319);
   U86918 : OAI221_X1 port map( B1 => n99949, B2 => n120014, C1 => n114413, C2 
                           => n120008, A => n117296, ZN => n117292);
   U86919 : AOI22_X1 port map( A1 => n120002, A2 => n118688, B1 => n119996, B2 
                           => n119320, ZN => n117296);
   U86920 : OAI221_X1 port map( B1 => n99948, B2 => n120014, C1 => n114412, C2 
                           => n120008, A => n117273, ZN => n117269);
   U86921 : AOI22_X1 port map( A1 => n120002, A2 => n118689, B1 => n119996, B2 
                           => n119321, ZN => n117273);
   U86922 : OAI221_X1 port map( B1 => n99947, B2 => n120014, C1 => n114411, C2 
                           => n120008, A => n117250, ZN => n117246);
   U86923 : AOI22_X1 port map( A1 => n120002, A2 => n118690, B1 => n119996, B2 
                           => n119322, ZN => n117250);
   U86924 : OAI221_X1 port map( B1 => n99946, B2 => n120014, C1 => n114410, C2 
                           => n120008, A => n117227, ZN => n117223);
   U86925 : AOI22_X1 port map( A1 => n120002, A2 => n118691, B1 => n119996, B2 
                           => n119323, ZN => n117227);
   U86926 : OAI221_X1 port map( B1 => n99945, B2 => n120014, C1 => n114409, C2 
                           => n120008, A => n117204, ZN => n117200);
   U86927 : AOI22_X1 port map( A1 => n120002, A2 => n118692, B1 => n119996, B2 
                           => n119324, ZN => n117204);
   U86928 : OAI221_X1 port map( B1 => n99944, B2 => n120014, C1 => n114408, C2 
                           => n120008, A => n117181, ZN => n117177);
   U86929 : AOI22_X1 port map( A1 => n120002, A2 => n118693, B1 => n119996, B2 
                           => n119325, ZN => n117181);
   U86930 : OAI221_X1 port map( B1 => n99943, B2 => n120014, C1 => n114407, C2 
                           => n120008, A => n117158, ZN => n117154);
   U86931 : AOI22_X1 port map( A1 => n120002, A2 => n118694, B1 => n119996, B2 
                           => n119326, ZN => n117158);
   U86932 : OAI221_X1 port map( B1 => n99942, B2 => n120015, C1 => n114406, C2 
                           => n120009, A => n117135, ZN => n117131);
   U86933 : AOI22_X1 port map( A1 => n120003, A2 => n118695, B1 => n119997, B2 
                           => n119327, ZN => n117135);
   U86934 : OAI221_X1 port map( B1 => n99941, B2 => n120015, C1 => n114405, C2 
                           => n120009, A => n117112, ZN => n117108);
   U86935 : AOI22_X1 port map( A1 => n120003, A2 => n118696, B1 => n119997, B2 
                           => n119328, ZN => n117112);
   U86936 : OAI221_X1 port map( B1 => n99940, B2 => n120015, C1 => n114404, C2 
                           => n120009, A => n117089, ZN => n117085);
   U86937 : AOI22_X1 port map( A1 => n120003, A2 => n118697, B1 => n119997, B2 
                           => n119329, ZN => n117089);
   U86938 : OAI221_X1 port map( B1 => n99939, B2 => n120015, C1 => n114403, C2 
                           => n120009, A => n117066, ZN => n117062);
   U86939 : AOI22_X1 port map( A1 => n120003, A2 => n118698, B1 => n119997, B2 
                           => n119330, ZN => n117066);
   U86940 : OAI221_X1 port map( B1 => n99938, B2 => n120015, C1 => n114402, C2 
                           => n120009, A => n117043, ZN => n117039);
   U86941 : AOI22_X1 port map( A1 => n120003, A2 => n118699, B1 => n119997, B2 
                           => n119331, ZN => n117043);
   U86942 : OAI221_X1 port map( B1 => n99937, B2 => n120015, C1 => n114401, C2 
                           => n120009, A => n117020, ZN => n117016);
   U86943 : AOI22_X1 port map( A1 => n120003, A2 => n118700, B1 => n119997, B2 
                           => n119332, ZN => n117020);
   U86944 : OAI221_X1 port map( B1 => n99936, B2 => n120015, C1 => n114400, C2 
                           => n120009, A => n116997, ZN => n116993);
   U86945 : AOI22_X1 port map( A1 => n120003, A2 => n118701, B1 => n119997, B2 
                           => n119333, ZN => n116997);
   U86946 : OAI221_X1 port map( B1 => n99935, B2 => n120015, C1 => n114399, C2 
                           => n120009, A => n116974, ZN => n116970);
   U86947 : AOI22_X1 port map( A1 => n120003, A2 => n118702, B1 => n119997, B2 
                           => n119334, ZN => n116974);
   U86948 : OAI221_X1 port map( B1 => n99934, B2 => n120015, C1 => n114398, C2 
                           => n120009, A => n116951, ZN => n116947);
   U86949 : AOI22_X1 port map( A1 => n120003, A2 => n118703, B1 => n119997, B2 
                           => n119335, ZN => n116951);
   U86950 : OAI221_X1 port map( B1 => n99933, B2 => n120015, C1 => n114397, C2 
                           => n120009, A => n116928, ZN => n116924);
   U86951 : AOI22_X1 port map( A1 => n120003, A2 => n118704, B1 => n119997, B2 
                           => n119336, ZN => n116928);
   U86952 : OAI221_X1 port map( B1 => n99932, B2 => n120015, C1 => n114396, C2 
                           => n120009, A => n116905, ZN => n116901);
   U86953 : AOI22_X1 port map( A1 => n120003, A2 => n118705, B1 => n119997, B2 
                           => n119337, ZN => n116905);
   U86954 : OAI221_X1 port map( B1 => n99931, B2 => n120015, C1 => n114395, C2 
                           => n120009, A => n116882, ZN => n116878);
   U86955 : AOI22_X1 port map( A1 => n120003, A2 => n118706, B1 => n119997, B2 
                           => n119338, ZN => n116882);
   U86956 : OAI221_X1 port map( B1 => n99930, B2 => n120016, C1 => n114394, C2 
                           => n120010, A => n116859, ZN => n116855);
   U86957 : AOI22_X1 port map( A1 => n120004, A2 => n118707, B1 => n119998, B2 
                           => n119339, ZN => n116859);
   U86958 : OAI221_X1 port map( B1 => n99929, B2 => n120016, C1 => n114393, C2 
                           => n120010, A => n116836, ZN => n116832);
   U86959 : AOI22_X1 port map( A1 => n120004, A2 => n118708, B1 => n119998, B2 
                           => n119340, ZN => n116836);
   U86960 : OAI221_X1 port map( B1 => n99928, B2 => n120016, C1 => n114392, C2 
                           => n120010, A => n116813, ZN => n116809);
   U86961 : AOI22_X1 port map( A1 => n120004, A2 => n118709, B1 => n119998, B2 
                           => n119341, ZN => n116813);
   U86962 : OAI221_X1 port map( B1 => n99927, B2 => n120016, C1 => n114391, C2 
                           => n120010, A => n116790, ZN => n116786);
   U86963 : AOI22_X1 port map( A1 => n120004, A2 => n118710, B1 => n119998, B2 
                           => n119342, ZN => n116790);
   U86964 : OAI221_X1 port map( B1 => n99926, B2 => n120016, C1 => n114390, C2 
                           => n120010, A => n116767, ZN => n116763);
   U86965 : AOI22_X1 port map( A1 => n120004, A2 => n118711, B1 => n119998, B2 
                           => n119343, ZN => n116767);
   U86966 : OAI221_X1 port map( B1 => n99925, B2 => n120016, C1 => n114389, C2 
                           => n120010, A => n116744, ZN => n116740);
   U86967 : AOI22_X1 port map( A1 => n120004, A2 => n118712, B1 => n119998, B2 
                           => n119344, ZN => n116744);
   U86968 : OAI221_X1 port map( B1 => n99924, B2 => n120016, C1 => n114388, C2 
                           => n120010, A => n116721, ZN => n116717);
   U86969 : AOI22_X1 port map( A1 => n120004, A2 => n118713, B1 => n119998, B2 
                           => n119345, ZN => n116721);
   U86970 : OAI221_X1 port map( B1 => n99923, B2 => n120016, C1 => n114387, C2 
                           => n120010, A => n116698, ZN => n116694);
   U86971 : AOI22_X1 port map( A1 => n120004, A2 => n118714, B1 => n119998, B2 
                           => n119346, ZN => n116698);
   U86972 : OAI221_X1 port map( B1 => n99922, B2 => n120016, C1 => n114386, C2 
                           => n120010, A => n116675, ZN => n116671);
   U86973 : AOI22_X1 port map( A1 => n120004, A2 => n118715, B1 => n119998, B2 
                           => n119347, ZN => n116675);
   U86974 : OAI221_X1 port map( B1 => n99921, B2 => n120016, C1 => n114385, C2 
                           => n120010, A => n116652, ZN => n116648);
   U86975 : AOI22_X1 port map( A1 => n120004, A2 => n118716, B1 => n119998, B2 
                           => n119348, ZN => n116652);
   U86976 : OAI221_X1 port map( B1 => n99920, B2 => n120016, C1 => n114384, C2 
                           => n120010, A => n116629, ZN => n116625);
   U86977 : AOI22_X1 port map( A1 => n120004, A2 => n118717, B1 => n119998, B2 
                           => n119349, ZN => n116629);
   U86978 : OAI221_X1 port map( B1 => n99919, B2 => n120016, C1 => n114383, C2 
                           => n120010, A => n116606, ZN => n116602);
   U86979 : AOI22_X1 port map( A1 => n120004, A2 => n118718, B1 => n119998, B2 
                           => n119350, ZN => n116606);
   U86980 : OAI221_X1 port map( B1 => n114150, B2 => n120215, C1 => n98652, C2 
                           => n120209, A => n114766, ZN => n114763);
   U86981 : AOI22_X1 port map( A1 => n120203, A2 => n118719, B1 => n120197, B2 
                           => n119298, ZN => n114766);
   U86982 : OAI221_X1 port map( B1 => n114149, B2 => n120215, C1 => n98651, C2 
                           => n120209, A => n114740, ZN => n114737);
   U86983 : AOI22_X1 port map( A1 => n120203, A2 => n118720, B1 => n120197, B2 
                           => n119299, ZN => n114740);
   U86984 : OAI221_X1 port map( B1 => n114148, B2 => n120215, C1 => n98650, C2 
                           => n120209, A => n114714, ZN => n114711);
   U86985 : AOI22_X1 port map( A1 => n120203, A2 => n118721, B1 => n120197, B2 
                           => n119300, ZN => n114714);
   U86986 : OAI221_X1 port map( B1 => n114146, B2 => n120215, C1 => n98648, C2 
                           => n120209, A => n114661, ZN => n114652);
   U86987 : AOI22_X1 port map( A1 => n120203, A2 => n118722, B1 => n120197, B2 
                           => n119301, ZN => n114661);
   U86988 : OAI221_X1 port map( B1 => n99918, B2 => n120017, C1 => n114382, C2 
                           => n120011, A => n116584, ZN => n116581);
   U86989 : AOI22_X1 port map( A1 => n120005, A2 => n118723, B1 => n119999, B2 
                           => n119351, ZN => n116584);
   U86990 : OAI221_X1 port map( B1 => n99917, B2 => n120017, C1 => n114381, C2 
                           => n120011, A => n116563, ZN => n116560);
   U86991 : AOI22_X1 port map( A1 => n120005, A2 => n118724, B1 => n119999, B2 
                           => n119352, ZN => n116563);
   U86992 : OAI221_X1 port map( B1 => n99916, B2 => n120017, C1 => n114380, C2 
                           => n120011, A => n116542, ZN => n116539);
   U86993 : AOI22_X1 port map( A1 => n120005, A2 => n118725, B1 => n119999, B2 
                           => n119353, ZN => n116542);
   U86994 : OAI221_X1 port map( B1 => n99914, B2 => n120017, C1 => n114378, C2 
                           => n120011, A => n116494, ZN => n116485);
   U86995 : AOI22_X1 port map( A1 => n120005, A2 => n118726, B1 => n119999, B2 
                           => n119354, ZN => n116494);
   U86996 : OAI221_X1 port map( B1 => n99971, B2 => n120012, C1 => n114435, C2 
                           => n120006, A => n117791, ZN => n117787);
   U86997 : AOI22_X1 port map( A1 => n120000, A2 => n118727, B1 => n119994, B2 
                           => n119355, ZN => n117791);
   U86998 : OAI221_X1 port map( B1 => n99970, B2 => n120012, C1 => n114434, C2 
                           => n120006, A => n117769, ZN => n117765);
   U86999 : AOI22_X1 port map( A1 => n120000, A2 => n118728, B1 => n119994, B2 
                           => n119356, ZN => n117769);
   U87000 : OAI221_X1 port map( B1 => n99969, B2 => n120012, C1 => n114433, C2 
                           => n120006, A => n117747, ZN => n117743);
   U87001 : AOI22_X1 port map( A1 => n120000, A2 => n118729, B1 => n119994, B2 
                           => n119357, ZN => n117747);
   U87002 : OAI221_X1 port map( B1 => n99968, B2 => n120012, C1 => n114432, C2 
                           => n120006, A => n117725, ZN => n117721);
   U87003 : AOI22_X1 port map( A1 => n120000, A2 => n118730, B1 => n119994, B2 
                           => n119358, ZN => n117725);
   U87004 : OAI221_X1 port map( B1 => n99978, B2 => n120012, C1 => n114442, C2 
                           => n120006, A => n117950, ZN => n117941);
   U87005 : AOI22_X1 port map( A1 => n120000, A2 => n118731, B1 => n119994, B2 
                           => n119359, ZN => n117950);
   U87006 : OAI221_X1 port map( B1 => n99977, B2 => n120012, C1 => n114441, C2 
                           => n120006, A => n117923, ZN => n117919);
   U87007 : AOI22_X1 port map( A1 => n120000, A2 => n118732, B1 => n119994, B2 
                           => n119360, ZN => n117923);
   U87008 : OAI221_X1 port map( B1 => n99976, B2 => n120012, C1 => n114440, C2 
                           => n120006, A => n117901, ZN => n117897);
   U87009 : AOI22_X1 port map( A1 => n120000, A2 => n118733, B1 => n119994, B2 
                           => n119361, ZN => n117901);
   U87010 : OAI221_X1 port map( B1 => n99975, B2 => n120012, C1 => n114439, C2 
                           => n120006, A => n117879, ZN => n117875);
   U87011 : AOI22_X1 port map( A1 => n120000, A2 => n118734, B1 => n119994, B2 
                           => n119362, ZN => n117879);
   U87012 : OAI221_X1 port map( B1 => n99974, B2 => n120012, C1 => n114438, C2 
                           => n120006, A => n117857, ZN => n117853);
   U87013 : AOI22_X1 port map( A1 => n120000, A2 => n118735, B1 => n119994, B2 
                           => n119363, ZN => n117857);
   U87014 : OAI221_X1 port map( B1 => n99973, B2 => n120012, C1 => n114437, C2 
                           => n120006, A => n117835, ZN => n117831);
   U87015 : AOI22_X1 port map( A1 => n120000, A2 => n118736, B1 => n119994, B2 
                           => n119364, ZN => n117835);
   U87016 : OAI221_X1 port map( B1 => n99972, B2 => n120012, C1 => n114436, C2 
                           => n120006, A => n117813, ZN => n117809);
   U87017 : AOI22_X1 port map( A1 => n120000, A2 => n118737, B1 => n119994, B2 
                           => n119365, ZN => n117813);
   U87018 : OAI22_X1 port map( A1 => n99780, A2 => n120323, B1 => n120631, B2 
                           => n120317, ZN => n5823);
   U87019 : OAI22_X1 port map( A1 => n99779, A2 => n120323, B1 => n120634, B2 
                           => n120317, ZN => n5824);
   U87020 : OAI22_X1 port map( A1 => n99778, A2 => n120323, B1 => n120637, B2 
                           => n120317, ZN => n5825);
   U87021 : OAI22_X1 port map( A1 => n99777, A2 => n120323, B1 => n120640, B2 
                           => n120317, ZN => n5826);
   U87022 : OAI22_X1 port map( A1 => n99776, A2 => n120323, B1 => n120643, B2 
                           => n120317, ZN => n5827);
   U87023 : OAI22_X1 port map( A1 => n99775, A2 => n120323, B1 => n120646, B2 
                           => n120317, ZN => n5828);
   U87024 : OAI22_X1 port map( A1 => n99774, A2 => n120323, B1 => n120649, B2 
                           => n120317, ZN => n5829);
   U87025 : OAI22_X1 port map( A1 => n99773, A2 => n120323, B1 => n120652, B2 
                           => n120317, ZN => n5830);
   U87026 : OAI22_X1 port map( A1 => n99772, A2 => n120323, B1 => n120655, B2 
                           => n120317, ZN => n5831);
   U87027 : OAI22_X1 port map( A1 => n99771, A2 => n120323, B1 => n120658, B2 
                           => n120317, ZN => n5832);
   U87028 : OAI22_X1 port map( A1 => n99770, A2 => n120323, B1 => n120661, B2 
                           => n120317, ZN => n5833);
   U87029 : OAI22_X1 port map( A1 => n99769, A2 => n120324, B1 => n120664, B2 
                           => n120317, ZN => n5834);
   U87030 : OAI22_X1 port map( A1 => n99768, A2 => n120324, B1 => n120667, B2 
                           => n120318, ZN => n5835);
   U87031 : OAI22_X1 port map( A1 => n99767, A2 => n120324, B1 => n120670, B2 
                           => n120318, ZN => n5836);
   U87032 : OAI22_X1 port map( A1 => n99766, A2 => n120324, B1 => n120673, B2 
                           => n120318, ZN => n5837);
   U87033 : OAI22_X1 port map( A1 => n99765, A2 => n120324, B1 => n120676, B2 
                           => n120318, ZN => n5838);
   U87034 : OAI22_X1 port map( A1 => n99764, A2 => n120324, B1 => n120679, B2 
                           => n120318, ZN => n5839);
   U87035 : OAI22_X1 port map( A1 => n99763, A2 => n120324, B1 => n120682, B2 
                           => n120318, ZN => n5840);
   U87036 : OAI22_X1 port map( A1 => n99762, A2 => n120324, B1 => n120685, B2 
                           => n120318, ZN => n5841);
   U87037 : OAI22_X1 port map( A1 => n99761, A2 => n120324, B1 => n120688, B2 
                           => n120318, ZN => n5842);
   U87038 : OAI22_X1 port map( A1 => n99760, A2 => n120324, B1 => n120691, B2 
                           => n120318, ZN => n5843);
   U87039 : OAI22_X1 port map( A1 => n99759, A2 => n120324, B1 => n120694, B2 
                           => n120318, ZN => n5844);
   U87040 : OAI22_X1 port map( A1 => n99758, A2 => n120324, B1 => n120697, B2 
                           => n120318, ZN => n5845);
   U87041 : OAI22_X1 port map( A1 => n99757, A2 => n120325, B1 => n120700, B2 
                           => n120318, ZN => n5846);
   U87042 : OAI22_X1 port map( A1 => n99756, A2 => n120325, B1 => n120703, B2 
                           => n120319, ZN => n5847);
   U87043 : OAI22_X1 port map( A1 => n99755, A2 => n120325, B1 => n120706, B2 
                           => n120319, ZN => n5848);
   U87044 : OAI22_X1 port map( A1 => n99754, A2 => n120325, B1 => n120709, B2 
                           => n120319, ZN => n5849);
   U87045 : OAI22_X1 port map( A1 => n99753, A2 => n120325, B1 => n120712, B2 
                           => n120319, ZN => n5850);
   U87046 : OAI22_X1 port map( A1 => n99752, A2 => n120325, B1 => n120715, B2 
                           => n120319, ZN => n5851);
   U87047 : OAI22_X1 port map( A1 => n99751, A2 => n120325, B1 => n120718, B2 
                           => n120319, ZN => n5852);
   U87048 : OAI22_X1 port map( A1 => n99750, A2 => n120325, B1 => n120721, B2 
                           => n120319, ZN => n5853);
   U87049 : OAI22_X1 port map( A1 => n99749, A2 => n120325, B1 => n120724, B2 
                           => n120319, ZN => n5854);
   U87050 : OAI22_X1 port map( A1 => n99748, A2 => n120325, B1 => n120727, B2 
                           => n120319, ZN => n5855);
   U87051 : OAI22_X1 port map( A1 => n99747, A2 => n120325, B1 => n120730, B2 
                           => n120319, ZN => n5856);
   U87052 : OAI22_X1 port map( A1 => n99746, A2 => n120325, B1 => n120733, B2 
                           => n120319, ZN => n5857);
   U87053 : OAI22_X1 port map( A1 => n99745, A2 => n120326, B1 => n120736, B2 
                           => n120319, ZN => n5858);
   U87054 : OAI22_X1 port map( A1 => n99744, A2 => n120326, B1 => n120739, B2 
                           => n120320, ZN => n5859);
   U87055 : OAI22_X1 port map( A1 => n99743, A2 => n120326, B1 => n120742, B2 
                           => n120320, ZN => n5860);
   U87056 : OAI22_X1 port map( A1 => n99742, A2 => n120326, B1 => n120745, B2 
                           => n120320, ZN => n5861);
   U87057 : OAI22_X1 port map( A1 => n99741, A2 => n120326, B1 => n120748, B2 
                           => n120320, ZN => n5862);
   U87058 : OAI22_X1 port map( A1 => n99740, A2 => n120326, B1 => n120751, B2 
                           => n120320, ZN => n5863);
   U87059 : OAI22_X1 port map( A1 => n99739, A2 => n120326, B1 => n120754, B2 
                           => n120320, ZN => n5864);
   U87060 : OAI22_X1 port map( A1 => n99738, A2 => n120326, B1 => n120757, B2 
                           => n120320, ZN => n5865);
   U87061 : OAI22_X1 port map( A1 => n99737, A2 => n120326, B1 => n120760, B2 
                           => n120320, ZN => n5866);
   U87062 : OAI22_X1 port map( A1 => n99736, A2 => n120326, B1 => n120763, B2 
                           => n120320, ZN => n5867);
   U87063 : OAI22_X1 port map( A1 => n99735, A2 => n120326, B1 => n120766, B2 
                           => n120320, ZN => n5868);
   U87064 : OAI22_X1 port map( A1 => n99734, A2 => n120326, B1 => n120769, B2 
                           => n120320, ZN => n5869);
   U87065 : OAI22_X1 port map( A1 => n99733, A2 => n120327, B1 => n120772, B2 
                           => n120320, ZN => n5870);
   U87066 : OAI22_X1 port map( A1 => n99732, A2 => n120327, B1 => n120775, B2 
                           => n120321, ZN => n5871);
   U87067 : OAI22_X1 port map( A1 => n99731, A2 => n120327, B1 => n120778, B2 
                           => n120321, ZN => n5872);
   U87068 : OAI22_X1 port map( A1 => n99730, A2 => n120327, B1 => n120781, B2 
                           => n120321, ZN => n5873);
   U87069 : OAI22_X1 port map( A1 => n99729, A2 => n120327, B1 => n120784, B2 
                           => n120321, ZN => n5874);
   U87070 : OAI22_X1 port map( A1 => n99728, A2 => n120327, B1 => n120787, B2 
                           => n120321, ZN => n5875);
   U87071 : OAI22_X1 port map( A1 => n99727, A2 => n120327, B1 => n120790, B2 
                           => n120321, ZN => n5876);
   U87072 : OAI22_X1 port map( A1 => n99726, A2 => n120327, B1 => n120793, B2 
                           => n120321, ZN => n5877);
   U87073 : OAI22_X1 port map( A1 => n99725, A2 => n120327, B1 => n120796, B2 
                           => n120321, ZN => n5878);
   U87074 : OAI22_X1 port map( A1 => n99724, A2 => n120327, B1 => n120799, B2 
                           => n120321, ZN => n5879);
   U87075 : OAI22_X1 port map( A1 => n99723, A2 => n120327, B1 => n120802, B2 
                           => n120321, ZN => n5880);
   U87076 : OAI22_X1 port map( A1 => n99722, A2 => n120327, B1 => n120805, B2 
                           => n120321, ZN => n5881);
   U87077 : OAI22_X1 port map( A1 => n99721, A2 => n120328, B1 => n120808, B2 
                           => n120321, ZN => n5882);
   U87078 : OAI22_X1 port map( A1 => n99978, A2 => n120272, B1 => n120631, B2 
                           => n120266, ZN => n5567);
   U87079 : OAI22_X1 port map( A1 => n99977, A2 => n120272, B1 => n120634, B2 
                           => n120266, ZN => n5568);
   U87080 : OAI22_X1 port map( A1 => n99976, A2 => n120272, B1 => n120637, B2 
                           => n120266, ZN => n5569);
   U87081 : OAI22_X1 port map( A1 => n99975, A2 => n120272, B1 => n120640, B2 
                           => n120266, ZN => n5570);
   U87082 : OAI22_X1 port map( A1 => n99974, A2 => n120272, B1 => n120643, B2 
                           => n120266, ZN => n5571);
   U87083 : OAI22_X1 port map( A1 => n99973, A2 => n120272, B1 => n120646, B2 
                           => n120266, ZN => n5572);
   U87084 : OAI22_X1 port map( A1 => n99972, A2 => n120272, B1 => n120649, B2 
                           => n120266, ZN => n5573);
   U87085 : OAI22_X1 port map( A1 => n99971, A2 => n120272, B1 => n120652, B2 
                           => n120266, ZN => n5574);
   U87086 : OAI22_X1 port map( A1 => n99970, A2 => n120272, B1 => n120655, B2 
                           => n120266, ZN => n5575);
   U87087 : OAI22_X1 port map( A1 => n99969, A2 => n120272, B1 => n120658, B2 
                           => n120266, ZN => n5576);
   U87088 : OAI22_X1 port map( A1 => n99968, A2 => n120272, B1 => n120661, B2 
                           => n120266, ZN => n5577);
   U87089 : OAI22_X1 port map( A1 => n99967, A2 => n120273, B1 => n120664, B2 
                           => n120266, ZN => n5578);
   U87090 : OAI22_X1 port map( A1 => n99966, A2 => n120273, B1 => n120667, B2 
                           => n120267, ZN => n5579);
   U87091 : OAI22_X1 port map( A1 => n99965, A2 => n120273, B1 => n120670, B2 
                           => n120267, ZN => n5580);
   U87092 : OAI22_X1 port map( A1 => n99964, A2 => n120273, B1 => n120673, B2 
                           => n120267, ZN => n5581);
   U87093 : OAI22_X1 port map( A1 => n99963, A2 => n120273, B1 => n120676, B2 
                           => n120267, ZN => n5582);
   U87094 : OAI22_X1 port map( A1 => n99962, A2 => n120273, B1 => n120679, B2 
                           => n120267, ZN => n5583);
   U87095 : OAI22_X1 port map( A1 => n99961, A2 => n120273, B1 => n120682, B2 
                           => n120267, ZN => n5584);
   U87096 : OAI22_X1 port map( A1 => n99960, A2 => n120273, B1 => n120685, B2 
                           => n120267, ZN => n5585);
   U87097 : OAI22_X1 port map( A1 => n99959, A2 => n120273, B1 => n120688, B2 
                           => n120267, ZN => n5586);
   U87098 : OAI22_X1 port map( A1 => n99958, A2 => n120273, B1 => n120691, B2 
                           => n120267, ZN => n5587);
   U87099 : OAI22_X1 port map( A1 => n99957, A2 => n120273, B1 => n120694, B2 
                           => n120267, ZN => n5588);
   U87100 : OAI22_X1 port map( A1 => n99956, A2 => n120273, B1 => n120697, B2 
                           => n120267, ZN => n5589);
   U87101 : OAI22_X1 port map( A1 => n99955, A2 => n120274, B1 => n120700, B2 
                           => n120267, ZN => n5590);
   U87102 : OAI22_X1 port map( A1 => n99954, A2 => n120274, B1 => n120703, B2 
                           => n120268, ZN => n5591);
   U87103 : OAI22_X1 port map( A1 => n99953, A2 => n120274, B1 => n120706, B2 
                           => n120268, ZN => n5592);
   U87104 : OAI22_X1 port map( A1 => n99952, A2 => n120274, B1 => n120709, B2 
                           => n120268, ZN => n5593);
   U87105 : OAI22_X1 port map( A1 => n99951, A2 => n120274, B1 => n120712, B2 
                           => n120268, ZN => n5594);
   U87106 : OAI22_X1 port map( A1 => n99950, A2 => n120274, B1 => n120715, B2 
                           => n120268, ZN => n5595);
   U87107 : OAI22_X1 port map( A1 => n99949, A2 => n120274, B1 => n120718, B2 
                           => n120268, ZN => n5596);
   U87108 : OAI22_X1 port map( A1 => n99948, A2 => n120274, B1 => n120721, B2 
                           => n120268, ZN => n5597);
   U87109 : OAI22_X1 port map( A1 => n99947, A2 => n120274, B1 => n120724, B2 
                           => n120268, ZN => n5598);
   U87110 : OAI22_X1 port map( A1 => n99946, A2 => n120274, B1 => n120727, B2 
                           => n120268, ZN => n5599);
   U87111 : OAI22_X1 port map( A1 => n99945, A2 => n120274, B1 => n120730, B2 
                           => n120268, ZN => n5600);
   U87112 : OAI22_X1 port map( A1 => n99944, A2 => n120274, B1 => n120733, B2 
                           => n120268, ZN => n5601);
   U87113 : OAI22_X1 port map( A1 => n99943, A2 => n120275, B1 => n120736, B2 
                           => n120268, ZN => n5602);
   U87114 : OAI22_X1 port map( A1 => n99942, A2 => n120275, B1 => n120739, B2 
                           => n120269, ZN => n5603);
   U87115 : OAI22_X1 port map( A1 => n99941, A2 => n120275, B1 => n120742, B2 
                           => n120269, ZN => n5604);
   U87116 : OAI22_X1 port map( A1 => n99940, A2 => n120275, B1 => n120745, B2 
                           => n120269, ZN => n5605);
   U87117 : OAI22_X1 port map( A1 => n99939, A2 => n120275, B1 => n120748, B2 
                           => n120269, ZN => n5606);
   U87118 : OAI22_X1 port map( A1 => n99938, A2 => n120275, B1 => n120751, B2 
                           => n120269, ZN => n5607);
   U87119 : OAI22_X1 port map( A1 => n99937, A2 => n120275, B1 => n120754, B2 
                           => n120269, ZN => n5608);
   U87120 : OAI22_X1 port map( A1 => n99936, A2 => n120275, B1 => n120757, B2 
                           => n120269, ZN => n5609);
   U87121 : OAI22_X1 port map( A1 => n99935, A2 => n120275, B1 => n120760, B2 
                           => n120269, ZN => n5610);
   U87122 : OAI22_X1 port map( A1 => n99934, A2 => n120275, B1 => n120763, B2 
                           => n120269, ZN => n5611);
   U87123 : OAI22_X1 port map( A1 => n99933, A2 => n120275, B1 => n120766, B2 
                           => n120269, ZN => n5612);
   U87124 : OAI22_X1 port map( A1 => n99932, A2 => n120275, B1 => n120769, B2 
                           => n120269, ZN => n5613);
   U87125 : OAI22_X1 port map( A1 => n99931, A2 => n120276, B1 => n120772, B2 
                           => n120269, ZN => n5614);
   U87126 : OAI22_X1 port map( A1 => n99930, A2 => n120276, B1 => n120775, B2 
                           => n120270, ZN => n5615);
   U87127 : OAI22_X1 port map( A1 => n99929, A2 => n120276, B1 => n120778, B2 
                           => n120270, ZN => n5616);
   U87128 : OAI22_X1 port map( A1 => n99928, A2 => n120276, B1 => n120781, B2 
                           => n120270, ZN => n5617);
   U87129 : OAI22_X1 port map( A1 => n99927, A2 => n120276, B1 => n120784, B2 
                           => n120270, ZN => n5618);
   U87130 : OAI22_X1 port map( A1 => n99926, A2 => n120276, B1 => n120787, B2 
                           => n120270, ZN => n5619);
   U87131 : OAI22_X1 port map( A1 => n99925, A2 => n120276, B1 => n120790, B2 
                           => n120270, ZN => n5620);
   U87132 : OAI22_X1 port map( A1 => n99924, A2 => n120276, B1 => n120793, B2 
                           => n120270, ZN => n5621);
   U87133 : OAI22_X1 port map( A1 => n99923, A2 => n120276, B1 => n120796, B2 
                           => n120270, ZN => n5622);
   U87134 : OAI22_X1 port map( A1 => n99922, A2 => n120276, B1 => n120799, B2 
                           => n120270, ZN => n5623);
   U87135 : OAI22_X1 port map( A1 => n99921, A2 => n120276, B1 => n120802, B2 
                           => n120270, ZN => n5624);
   U87136 : OAI22_X1 port map( A1 => n99920, A2 => n120276, B1 => n120805, B2 
                           => n120270, ZN => n5625);
   U87137 : OAI22_X1 port map( A1 => n99919, A2 => n120277, B1 => n120808, B2 
                           => n120270, ZN => n5626);
   U87138 : OAI22_X1 port map( A1 => n99243, A2 => n120470, B1 => n120630, B2 
                           => n120464, ZN => n6591);
   U87139 : OAI22_X1 port map( A1 => n99242, A2 => n120470, B1 => n120633, B2 
                           => n120464, ZN => n6592);
   U87140 : OAI22_X1 port map( A1 => n99241, A2 => n120470, B1 => n120636, B2 
                           => n120464, ZN => n6593);
   U87141 : OAI22_X1 port map( A1 => n99240, A2 => n120470, B1 => n120639, B2 
                           => n120464, ZN => n6594);
   U87142 : OAI22_X1 port map( A1 => n99239, A2 => n120470, B1 => n120642, B2 
                           => n120464, ZN => n6595);
   U87143 : OAI22_X1 port map( A1 => n99238, A2 => n120470, B1 => n120645, B2 
                           => n120464, ZN => n6596);
   U87144 : OAI22_X1 port map( A1 => n99237, A2 => n120470, B1 => n120648, B2 
                           => n120464, ZN => n6597);
   U87145 : OAI22_X1 port map( A1 => n99236, A2 => n120470, B1 => n120651, B2 
                           => n120464, ZN => n6598);
   U87146 : OAI22_X1 port map( A1 => n99235, A2 => n120470, B1 => n120654, B2 
                           => n120464, ZN => n6599);
   U87147 : OAI22_X1 port map( A1 => n99234, A2 => n120470, B1 => n120657, B2 
                           => n120464, ZN => n6600);
   U87148 : OAI22_X1 port map( A1 => n99233, A2 => n120470, B1 => n120660, B2 
                           => n120464, ZN => n6601);
   U87149 : OAI22_X1 port map( A1 => n99232, A2 => n120471, B1 => n120663, B2 
                           => n120464, ZN => n6602);
   U87150 : OAI22_X1 port map( A1 => n99231, A2 => n120471, B1 => n120666, B2 
                           => n120465, ZN => n6603);
   U87151 : OAI22_X1 port map( A1 => n99230, A2 => n120471, B1 => n120669, B2 
                           => n120465, ZN => n6604);
   U87152 : OAI22_X1 port map( A1 => n99229, A2 => n120471, B1 => n120672, B2 
                           => n120465, ZN => n6605);
   U87153 : OAI22_X1 port map( A1 => n99228, A2 => n120471, B1 => n120675, B2 
                           => n120465, ZN => n6606);
   U87154 : OAI22_X1 port map( A1 => n99227, A2 => n120471, B1 => n120678, B2 
                           => n120465, ZN => n6607);
   U87155 : OAI22_X1 port map( A1 => n99226, A2 => n120471, B1 => n120681, B2 
                           => n120465, ZN => n6608);
   U87156 : OAI22_X1 port map( A1 => n99225, A2 => n120471, B1 => n120684, B2 
                           => n120465, ZN => n6609);
   U87157 : OAI22_X1 port map( A1 => n99224, A2 => n120471, B1 => n120687, B2 
                           => n120465, ZN => n6610);
   U87158 : OAI22_X1 port map( A1 => n99223, A2 => n120471, B1 => n120690, B2 
                           => n120465, ZN => n6611);
   U87159 : OAI22_X1 port map( A1 => n99222, A2 => n120471, B1 => n120693, B2 
                           => n120465, ZN => n6612);
   U87160 : OAI22_X1 port map( A1 => n99221, A2 => n120471, B1 => n120696, B2 
                           => n120465, ZN => n6613);
   U87161 : OAI22_X1 port map( A1 => n99220, A2 => n120472, B1 => n120699, B2 
                           => n120465, ZN => n6614);
   U87162 : OAI22_X1 port map( A1 => n99219, A2 => n120472, B1 => n120702, B2 
                           => n120466, ZN => n6615);
   U87163 : OAI22_X1 port map( A1 => n99218, A2 => n120472, B1 => n120705, B2 
                           => n120466, ZN => n6616);
   U87164 : OAI22_X1 port map( A1 => n99217, A2 => n120472, B1 => n120708, B2 
                           => n120466, ZN => n6617);
   U87165 : OAI22_X1 port map( A1 => n99216, A2 => n120472, B1 => n120711, B2 
                           => n120466, ZN => n6618);
   U87166 : OAI22_X1 port map( A1 => n99215, A2 => n120472, B1 => n120714, B2 
                           => n120466, ZN => n6619);
   U87167 : OAI22_X1 port map( A1 => n99214, A2 => n120472, B1 => n120717, B2 
                           => n120466, ZN => n6620);
   U87168 : OAI22_X1 port map( A1 => n99213, A2 => n120472, B1 => n120720, B2 
                           => n120466, ZN => n6621);
   U87169 : OAI22_X1 port map( A1 => n99212, A2 => n120472, B1 => n120723, B2 
                           => n120466, ZN => n6622);
   U87170 : OAI22_X1 port map( A1 => n99211, A2 => n120472, B1 => n120726, B2 
                           => n120466, ZN => n6623);
   U87171 : OAI22_X1 port map( A1 => n99210, A2 => n120472, B1 => n120729, B2 
                           => n120466, ZN => n6624);
   U87172 : OAI22_X1 port map( A1 => n99209, A2 => n120472, B1 => n120732, B2 
                           => n120466, ZN => n6625);
   U87173 : OAI22_X1 port map( A1 => n99208, A2 => n120473, B1 => n120735, B2 
                           => n120466, ZN => n6626);
   U87174 : OAI22_X1 port map( A1 => n99207, A2 => n120473, B1 => n120738, B2 
                           => n120467, ZN => n6627);
   U87175 : OAI22_X1 port map( A1 => n99206, A2 => n120473, B1 => n120741, B2 
                           => n120467, ZN => n6628);
   U87176 : OAI22_X1 port map( A1 => n99205, A2 => n120473, B1 => n120744, B2 
                           => n120467, ZN => n6629);
   U87177 : OAI22_X1 port map( A1 => n99204, A2 => n120473, B1 => n120747, B2 
                           => n120467, ZN => n6630);
   U87178 : OAI22_X1 port map( A1 => n99203, A2 => n120473, B1 => n120750, B2 
                           => n120467, ZN => n6631);
   U87179 : OAI22_X1 port map( A1 => n99202, A2 => n120473, B1 => n120753, B2 
                           => n120467, ZN => n6632);
   U87180 : OAI22_X1 port map( A1 => n99201, A2 => n120473, B1 => n120756, B2 
                           => n120467, ZN => n6633);
   U87181 : OAI22_X1 port map( A1 => n99200, A2 => n120473, B1 => n120759, B2 
                           => n120467, ZN => n6634);
   U87182 : OAI22_X1 port map( A1 => n99199, A2 => n120473, B1 => n120762, B2 
                           => n120467, ZN => n6635);
   U87183 : OAI22_X1 port map( A1 => n99198, A2 => n120473, B1 => n120765, B2 
                           => n120467, ZN => n6636);
   U87184 : OAI22_X1 port map( A1 => n99197, A2 => n120473, B1 => n120768, B2 
                           => n120467, ZN => n6637);
   U87185 : OAI22_X1 port map( A1 => n99196, A2 => n120474, B1 => n120771, B2 
                           => n120467, ZN => n6638);
   U87186 : OAI22_X1 port map( A1 => n99195, A2 => n120474, B1 => n120774, B2 
                           => n120468, ZN => n6639);
   U87187 : OAI22_X1 port map( A1 => n99194, A2 => n120474, B1 => n120777, B2 
                           => n120468, ZN => n6640);
   U87188 : OAI22_X1 port map( A1 => n99193, A2 => n120474, B1 => n120780, B2 
                           => n120468, ZN => n6641);
   U87189 : OAI22_X1 port map( A1 => n99192, A2 => n120474, B1 => n120783, B2 
                           => n120468, ZN => n6642);
   U87190 : OAI22_X1 port map( A1 => n99191, A2 => n120474, B1 => n120786, B2 
                           => n120468, ZN => n6643);
   U87191 : OAI22_X1 port map( A1 => n99190, A2 => n120474, B1 => n120789, B2 
                           => n120468, ZN => n6644);
   U87192 : OAI22_X1 port map( A1 => n99189, A2 => n120474, B1 => n120792, B2 
                           => n120468, ZN => n6645);
   U87193 : OAI22_X1 port map( A1 => n99188, A2 => n120474, B1 => n120795, B2 
                           => n120468, ZN => n6646);
   U87194 : OAI22_X1 port map( A1 => n99187, A2 => n120474, B1 => n120798, B2 
                           => n120468, ZN => n6647);
   U87195 : OAI22_X1 port map( A1 => n99186, A2 => n120474, B1 => n120801, B2 
                           => n120468, ZN => n6648);
   U87196 : OAI22_X1 port map( A1 => n99185, A2 => n120474, B1 => n120804, B2 
                           => n120468, ZN => n6649);
   U87197 : OAI22_X1 port map( A1 => n99184, A2 => n120475, B1 => n120807, B2 
                           => n120468, ZN => n6650);
   U87198 : OAI22_X1 port map( A1 => n99375, A2 => n120446, B1 => n120630, B2 
                           => n120440, ZN => n6463);
   U87199 : OAI22_X1 port map( A1 => n99374, A2 => n120446, B1 => n120633, B2 
                           => n120440, ZN => n6464);
   U87200 : OAI22_X1 port map( A1 => n99373, A2 => n120446, B1 => n120636, B2 
                           => n120440, ZN => n6465);
   U87201 : OAI22_X1 port map( A1 => n99372, A2 => n120446, B1 => n120639, B2 
                           => n120440, ZN => n6466);
   U87202 : OAI22_X1 port map( A1 => n99371, A2 => n120446, B1 => n120642, B2 
                           => n120440, ZN => n6467);
   U87203 : OAI22_X1 port map( A1 => n99370, A2 => n120446, B1 => n120645, B2 
                           => n120440, ZN => n6468);
   U87204 : OAI22_X1 port map( A1 => n99369, A2 => n120446, B1 => n120648, B2 
                           => n120440, ZN => n6469);
   U87205 : OAI22_X1 port map( A1 => n99368, A2 => n120446, B1 => n120651, B2 
                           => n120440, ZN => n6470);
   U87206 : OAI22_X1 port map( A1 => n99367, A2 => n120446, B1 => n120654, B2 
                           => n120440, ZN => n6471);
   U87207 : OAI22_X1 port map( A1 => n99366, A2 => n120446, B1 => n120657, B2 
                           => n120440, ZN => n6472);
   U87208 : OAI22_X1 port map( A1 => n99365, A2 => n120446, B1 => n120660, B2 
                           => n120440, ZN => n6473);
   U87209 : OAI22_X1 port map( A1 => n99364, A2 => n120447, B1 => n120663, B2 
                           => n120440, ZN => n6474);
   U87210 : OAI22_X1 port map( A1 => n99363, A2 => n120447, B1 => n120666, B2 
                           => n120441, ZN => n6475);
   U87211 : OAI22_X1 port map( A1 => n99362, A2 => n120447, B1 => n120669, B2 
                           => n120441, ZN => n6476);
   U87212 : OAI22_X1 port map( A1 => n99361, A2 => n120447, B1 => n120672, B2 
                           => n120441, ZN => n6477);
   U87213 : OAI22_X1 port map( A1 => n99360, A2 => n120447, B1 => n120675, B2 
                           => n120441, ZN => n6478);
   U87214 : OAI22_X1 port map( A1 => n99359, A2 => n120447, B1 => n120678, B2 
                           => n120441, ZN => n6479);
   U87215 : OAI22_X1 port map( A1 => n99358, A2 => n120447, B1 => n120681, B2 
                           => n120441, ZN => n6480);
   U87216 : OAI22_X1 port map( A1 => n99357, A2 => n120447, B1 => n120684, B2 
                           => n120441, ZN => n6481);
   U87217 : OAI22_X1 port map( A1 => n99356, A2 => n120447, B1 => n120687, B2 
                           => n120441, ZN => n6482);
   U87218 : OAI22_X1 port map( A1 => n99355, A2 => n120447, B1 => n120690, B2 
                           => n120441, ZN => n6483);
   U87219 : OAI22_X1 port map( A1 => n99354, A2 => n120447, B1 => n120693, B2 
                           => n120441, ZN => n6484);
   U87220 : OAI22_X1 port map( A1 => n99353, A2 => n120447, B1 => n120696, B2 
                           => n120441, ZN => n6485);
   U87221 : OAI22_X1 port map( A1 => n99352, A2 => n120448, B1 => n120699, B2 
                           => n120441, ZN => n6486);
   U87222 : OAI22_X1 port map( A1 => n99351, A2 => n120448, B1 => n120702, B2 
                           => n120442, ZN => n6487);
   U87223 : OAI22_X1 port map( A1 => n99350, A2 => n120448, B1 => n120705, B2 
                           => n120442, ZN => n6488);
   U87224 : OAI22_X1 port map( A1 => n99349, A2 => n120448, B1 => n120708, B2 
                           => n120442, ZN => n6489);
   U87225 : OAI22_X1 port map( A1 => n99348, A2 => n120448, B1 => n120711, B2 
                           => n120442, ZN => n6490);
   U87226 : OAI22_X1 port map( A1 => n99347, A2 => n120448, B1 => n120714, B2 
                           => n120442, ZN => n6491);
   U87227 : OAI22_X1 port map( A1 => n99346, A2 => n120448, B1 => n120717, B2 
                           => n120442, ZN => n6492);
   U87228 : OAI22_X1 port map( A1 => n99345, A2 => n120448, B1 => n120720, B2 
                           => n120442, ZN => n6493);
   U87229 : OAI22_X1 port map( A1 => n99344, A2 => n120448, B1 => n120723, B2 
                           => n120442, ZN => n6494);
   U87230 : OAI22_X1 port map( A1 => n99343, A2 => n120448, B1 => n120726, B2 
                           => n120442, ZN => n6495);
   U87231 : OAI22_X1 port map( A1 => n99342, A2 => n120448, B1 => n120729, B2 
                           => n120442, ZN => n6496);
   U87232 : OAI22_X1 port map( A1 => n99341, A2 => n120448, B1 => n120732, B2 
                           => n120442, ZN => n6497);
   U87233 : OAI22_X1 port map( A1 => n99340, A2 => n120449, B1 => n120735, B2 
                           => n120442, ZN => n6498);
   U87234 : OAI22_X1 port map( A1 => n99339, A2 => n120449, B1 => n120738, B2 
                           => n120443, ZN => n6499);
   U87235 : OAI22_X1 port map( A1 => n99338, A2 => n120449, B1 => n120741, B2 
                           => n120443, ZN => n6500);
   U87236 : OAI22_X1 port map( A1 => n99337, A2 => n120449, B1 => n120744, B2 
                           => n120443, ZN => n6501);
   U87237 : OAI22_X1 port map( A1 => n99336, A2 => n120449, B1 => n120747, B2 
                           => n120443, ZN => n6502);
   U87238 : OAI22_X1 port map( A1 => n99335, A2 => n120449, B1 => n120750, B2 
                           => n120443, ZN => n6503);
   U87239 : OAI22_X1 port map( A1 => n99334, A2 => n120449, B1 => n120753, B2 
                           => n120443, ZN => n6504);
   U87240 : OAI22_X1 port map( A1 => n99333, A2 => n120449, B1 => n120756, B2 
                           => n120443, ZN => n6505);
   U87241 : OAI22_X1 port map( A1 => n99332, A2 => n120449, B1 => n120759, B2 
                           => n120443, ZN => n6506);
   U87242 : OAI22_X1 port map( A1 => n99331, A2 => n120449, B1 => n120762, B2 
                           => n120443, ZN => n6507);
   U87243 : OAI22_X1 port map( A1 => n99330, A2 => n120449, B1 => n120765, B2 
                           => n120443, ZN => n6508);
   U87244 : OAI22_X1 port map( A1 => n99329, A2 => n120449, B1 => n120768, B2 
                           => n120443, ZN => n6509);
   U87245 : OAI22_X1 port map( A1 => n99328, A2 => n120450, B1 => n120771, B2 
                           => n120443, ZN => n6510);
   U87246 : OAI22_X1 port map( A1 => n99327, A2 => n120450, B1 => n120774, B2 
                           => n120444, ZN => n6511);
   U87247 : OAI22_X1 port map( A1 => n99326, A2 => n120450, B1 => n120777, B2 
                           => n120444, ZN => n6512);
   U87248 : OAI22_X1 port map( A1 => n99325, A2 => n120450, B1 => n120780, B2 
                           => n120444, ZN => n6513);
   U87249 : OAI22_X1 port map( A1 => n99324, A2 => n120450, B1 => n120783, B2 
                           => n120444, ZN => n6514);
   U87250 : OAI22_X1 port map( A1 => n99323, A2 => n120450, B1 => n120786, B2 
                           => n120444, ZN => n6515);
   U87251 : OAI22_X1 port map( A1 => n99322, A2 => n120450, B1 => n120789, B2 
                           => n120444, ZN => n6516);
   U87252 : OAI22_X1 port map( A1 => n99321, A2 => n120450, B1 => n120792, B2 
                           => n120444, ZN => n6517);
   U87253 : OAI22_X1 port map( A1 => n99320, A2 => n120450, B1 => n120795, B2 
                           => n120444, ZN => n6518);
   U87254 : OAI22_X1 port map( A1 => n99319, A2 => n120450, B1 => n120798, B2 
                           => n120444, ZN => n6519);
   U87255 : OAI22_X1 port map( A1 => n99318, A2 => n120450, B1 => n120801, B2 
                           => n120444, ZN => n6520);
   U87256 : OAI22_X1 port map( A1 => n99317, A2 => n120450, B1 => n120804, B2 
                           => n120444, ZN => n6521);
   U87257 : OAI22_X1 port map( A1 => n99316, A2 => n120451, B1 => n120807, B2 
                           => n120444, ZN => n6522);
   U87258 : OAI22_X1 port map( A1 => n120520, A2 => n114120, B1 => n120629, B2 
                           => n120512, ZN => n6847);
   U87259 : OAI22_X1 port map( A1 => n120520, A2 => n114119, B1 => n120632, B2 
                           => n120512, ZN => n6848);
   U87260 : OAI22_X1 port map( A1 => n120520, A2 => n114118, B1 => n120635, B2 
                           => n120512, ZN => n6849);
   U87261 : OAI22_X1 port map( A1 => n120520, A2 => n114117, B1 => n120638, B2 
                           => n120512, ZN => n6850);
   U87262 : OAI22_X1 port map( A1 => n120520, A2 => n114116, B1 => n120641, B2 
                           => n120512, ZN => n6851);
   U87263 : OAI22_X1 port map( A1 => n120520, A2 => n114115, B1 => n120644, B2 
                           => n120512, ZN => n6852);
   U87264 : OAI22_X1 port map( A1 => n120520, A2 => n114114, B1 => n120647, B2 
                           => n120512, ZN => n6853);
   U87265 : OAI22_X1 port map( A1 => n120520, A2 => n114113, B1 => n120650, B2 
                           => n120512, ZN => n6854);
   U87266 : OAI22_X1 port map( A1 => n120520, A2 => n114112, B1 => n120653, B2 
                           => n120512, ZN => n6855);
   U87267 : OAI22_X1 port map( A1 => n120520, A2 => n114111, B1 => n120656, B2 
                           => n120512, ZN => n6856);
   U87268 : OAI22_X1 port map( A1 => n120520, A2 => n114110, B1 => n120659, B2 
                           => n120512, ZN => n6857);
   U87269 : OAI22_X1 port map( A1 => n120520, A2 => n114109, B1 => n120662, B2 
                           => n120512, ZN => n6858);
   U87270 : OAI22_X1 port map( A1 => n120521, A2 => n114108, B1 => n120665, B2 
                           => n120513, ZN => n6859);
   U87271 : OAI22_X1 port map( A1 => n120521, A2 => n114107, B1 => n120668, B2 
                           => n120513, ZN => n6860);
   U87272 : OAI22_X1 port map( A1 => n120521, A2 => n114106, B1 => n120671, B2 
                           => n120513, ZN => n6861);
   U87273 : OAI22_X1 port map( A1 => n120521, A2 => n114105, B1 => n120674, B2 
                           => n120513, ZN => n6862);
   U87274 : OAI22_X1 port map( A1 => n120521, A2 => n114104, B1 => n120677, B2 
                           => n120513, ZN => n6863);
   U87275 : OAI22_X1 port map( A1 => n120521, A2 => n114103, B1 => n120680, B2 
                           => n120513, ZN => n6864);
   U87276 : OAI22_X1 port map( A1 => n120521, A2 => n114102, B1 => n120683, B2 
                           => n120513, ZN => n6865);
   U87277 : OAI22_X1 port map( A1 => n120521, A2 => n114101, B1 => n120686, B2 
                           => n120513, ZN => n6866);
   U87278 : OAI22_X1 port map( A1 => n120521, A2 => n114100, B1 => n120689, B2 
                           => n120513, ZN => n6867);
   U87279 : OAI22_X1 port map( A1 => n120521, A2 => n114099, B1 => n120692, B2 
                           => n120513, ZN => n6868);
   U87280 : OAI22_X1 port map( A1 => n120521, A2 => n114098, B1 => n120695, B2 
                           => n120513, ZN => n6869);
   U87281 : OAI22_X1 port map( A1 => n120521, A2 => n114097, B1 => n120698, B2 
                           => n120513, ZN => n6870);
   U87282 : OAI22_X1 port map( A1 => n120521, A2 => n114096, B1 => n120701, B2 
                           => n120514, ZN => n6871);
   U87283 : OAI22_X1 port map( A1 => n120522, A2 => n114095, B1 => n120704, B2 
                           => n120514, ZN => n6872);
   U87284 : OAI22_X1 port map( A1 => n120522, A2 => n114094, B1 => n120707, B2 
                           => n120514, ZN => n6873);
   U87285 : OAI22_X1 port map( A1 => n120522, A2 => n114093, B1 => n120710, B2 
                           => n120514, ZN => n6874);
   U87286 : OAI22_X1 port map( A1 => n120522, A2 => n114092, B1 => n120713, B2 
                           => n120514, ZN => n6875);
   U87287 : OAI22_X1 port map( A1 => n120522, A2 => n114091, B1 => n120716, B2 
                           => n120514, ZN => n6876);
   U87288 : OAI22_X1 port map( A1 => n120522, A2 => n114090, B1 => n120719, B2 
                           => n120514, ZN => n6877);
   U87289 : OAI22_X1 port map( A1 => n120522, A2 => n114089, B1 => n120722, B2 
                           => n120514, ZN => n6878);
   U87290 : OAI22_X1 port map( A1 => n120522, A2 => n114088, B1 => n120725, B2 
                           => n120514, ZN => n6879);
   U87291 : OAI22_X1 port map( A1 => n120522, A2 => n114087, B1 => n120728, B2 
                           => n120514, ZN => n6880);
   U87292 : OAI22_X1 port map( A1 => n120522, A2 => n114086, B1 => n120731, B2 
                           => n120514, ZN => n6881);
   U87293 : OAI22_X1 port map( A1 => n120522, A2 => n114085, B1 => n120734, B2 
                           => n120514, ZN => n6882);
   U87294 : OAI22_X1 port map( A1 => n120522, A2 => n114084, B1 => n120737, B2 
                           => n120515, ZN => n6883);
   U87295 : OAI22_X1 port map( A1 => n120522, A2 => n114083, B1 => n120740, B2 
                           => n120515, ZN => n6884);
   U87296 : OAI22_X1 port map( A1 => n120523, A2 => n114082, B1 => n120743, B2 
                           => n120515, ZN => n6885);
   U87297 : OAI22_X1 port map( A1 => n120523, A2 => n114081, B1 => n120746, B2 
                           => n120515, ZN => n6886);
   U87298 : OAI22_X1 port map( A1 => n120523, A2 => n114080, B1 => n120749, B2 
                           => n120515, ZN => n6887);
   U87299 : OAI22_X1 port map( A1 => n120523, A2 => n114079, B1 => n120752, B2 
                           => n120515, ZN => n6888);
   U87300 : OAI22_X1 port map( A1 => n120523, A2 => n114078, B1 => n120755, B2 
                           => n120515, ZN => n6889);
   U87301 : OAI22_X1 port map( A1 => n120523, A2 => n114077, B1 => n120758, B2 
                           => n120515, ZN => n6890);
   U87302 : OAI22_X1 port map( A1 => n120523, A2 => n114076, B1 => n120761, B2 
                           => n120515, ZN => n6891);
   U87303 : OAI22_X1 port map( A1 => n120523, A2 => n114075, B1 => n120764, B2 
                           => n120515, ZN => n6892);
   U87304 : OAI22_X1 port map( A1 => n120523, A2 => n114074, B1 => n120767, B2 
                           => n120515, ZN => n6893);
   U87305 : OAI22_X1 port map( A1 => n120523, A2 => n114073, B1 => n120770, B2 
                           => n120515, ZN => n6894);
   U87306 : OAI22_X1 port map( A1 => n120523, A2 => n114072, B1 => n120773, B2 
                           => n120516, ZN => n6895);
   U87307 : OAI22_X1 port map( A1 => n120523, A2 => n114071, B1 => n120776, B2 
                           => n120516, ZN => n6896);
   U87308 : OAI22_X1 port map( A1 => n120523, A2 => n114070, B1 => n120779, B2 
                           => n120516, ZN => n6897);
   U87309 : OAI22_X1 port map( A1 => n120524, A2 => n114069, B1 => n120782, B2 
                           => n120516, ZN => n6898);
   U87310 : OAI22_X1 port map( A1 => n120524, A2 => n114068, B1 => n120785, B2 
                           => n120516, ZN => n6899);
   U87311 : OAI22_X1 port map( A1 => n120524, A2 => n114067, B1 => n120788, B2 
                           => n120516, ZN => n6900);
   U87312 : OAI22_X1 port map( A1 => n120524, A2 => n114066, B1 => n120791, B2 
                           => n120516, ZN => n6901);
   U87313 : OAI22_X1 port map( A1 => n120524, A2 => n114065, B1 => n120794, B2 
                           => n120516, ZN => n6902);
   U87314 : OAI22_X1 port map( A1 => n120524, A2 => n114064, B1 => n120797, B2 
                           => n120516, ZN => n6903);
   U87315 : OAI22_X1 port map( A1 => n120524, A2 => n114063, B1 => n120800, B2 
                           => n120516, ZN => n6904);
   U87316 : OAI22_X1 port map( A1 => n120524, A2 => n114062, B1 => n120803, B2 
                           => n120516, ZN => n6905);
   U87317 : OAI22_X1 port map( A1 => n120524, A2 => n114061, B1 => n120806, B2 
                           => n120516, ZN => n6906);
   U87318 : OAI22_X1 port map( A1 => n99111, A2 => n120494, B1 => n120629, B2 
                           => n120488, ZN => n6719);
   U87319 : OAI22_X1 port map( A1 => n99110, A2 => n120494, B1 => n120632, B2 
                           => n120488, ZN => n6720);
   U87320 : OAI22_X1 port map( A1 => n99109, A2 => n120494, B1 => n120635, B2 
                           => n120488, ZN => n6721);
   U87321 : OAI22_X1 port map( A1 => n99108, A2 => n120494, B1 => n120638, B2 
                           => n120488, ZN => n6722);
   U87322 : OAI22_X1 port map( A1 => n99107, A2 => n120494, B1 => n120641, B2 
                           => n120488, ZN => n6723);
   U87323 : OAI22_X1 port map( A1 => n99106, A2 => n120494, B1 => n120644, B2 
                           => n120488, ZN => n6724);
   U87324 : OAI22_X1 port map( A1 => n99105, A2 => n120494, B1 => n120647, B2 
                           => n120488, ZN => n6725);
   U87325 : OAI22_X1 port map( A1 => n99104, A2 => n120494, B1 => n120650, B2 
                           => n120488, ZN => n6726);
   U87326 : OAI22_X1 port map( A1 => n99103, A2 => n120494, B1 => n120653, B2 
                           => n120488, ZN => n6727);
   U87327 : OAI22_X1 port map( A1 => n99102, A2 => n120494, B1 => n120656, B2 
                           => n120488, ZN => n6728);
   U87328 : OAI22_X1 port map( A1 => n99101, A2 => n120494, B1 => n120659, B2 
                           => n120488, ZN => n6729);
   U87329 : OAI22_X1 port map( A1 => n99100, A2 => n120495, B1 => n120662, B2 
                           => n120488, ZN => n6730);
   U87330 : OAI22_X1 port map( A1 => n99099, A2 => n120495, B1 => n120665, B2 
                           => n120489, ZN => n6731);
   U87331 : OAI22_X1 port map( A1 => n99098, A2 => n120495, B1 => n120668, B2 
                           => n120489, ZN => n6732);
   U87332 : OAI22_X1 port map( A1 => n99097, A2 => n120495, B1 => n120671, B2 
                           => n120489, ZN => n6733);
   U87333 : OAI22_X1 port map( A1 => n99096, A2 => n120495, B1 => n120674, B2 
                           => n120489, ZN => n6734);
   U87334 : OAI22_X1 port map( A1 => n99095, A2 => n120495, B1 => n120677, B2 
                           => n120489, ZN => n6735);
   U87335 : OAI22_X1 port map( A1 => n99094, A2 => n120495, B1 => n120680, B2 
                           => n120489, ZN => n6736);
   U87336 : OAI22_X1 port map( A1 => n99093, A2 => n120495, B1 => n120683, B2 
                           => n120489, ZN => n6737);
   U87337 : OAI22_X1 port map( A1 => n99092, A2 => n120495, B1 => n120686, B2 
                           => n120489, ZN => n6738);
   U87338 : OAI22_X1 port map( A1 => n99091, A2 => n120495, B1 => n120689, B2 
                           => n120489, ZN => n6739);
   U87339 : OAI22_X1 port map( A1 => n99090, A2 => n120495, B1 => n120692, B2 
                           => n120489, ZN => n6740);
   U87340 : OAI22_X1 port map( A1 => n99089, A2 => n120495, B1 => n120695, B2 
                           => n120489, ZN => n6741);
   U87341 : OAI22_X1 port map( A1 => n99088, A2 => n120496, B1 => n120698, B2 
                           => n120489, ZN => n6742);
   U87342 : OAI22_X1 port map( A1 => n99087, A2 => n120496, B1 => n120701, B2 
                           => n120490, ZN => n6743);
   U87343 : OAI22_X1 port map( A1 => n99086, A2 => n120496, B1 => n120704, B2 
                           => n120490, ZN => n6744);
   U87344 : OAI22_X1 port map( A1 => n99085, A2 => n120496, B1 => n120707, B2 
                           => n120490, ZN => n6745);
   U87345 : OAI22_X1 port map( A1 => n99084, A2 => n120496, B1 => n120710, B2 
                           => n120490, ZN => n6746);
   U87346 : OAI22_X1 port map( A1 => n99083, A2 => n120496, B1 => n120713, B2 
                           => n120490, ZN => n6747);
   U87347 : OAI22_X1 port map( A1 => n99082, A2 => n120496, B1 => n120716, B2 
                           => n120490, ZN => n6748);
   U87348 : OAI22_X1 port map( A1 => n99081, A2 => n120496, B1 => n120719, B2 
                           => n120490, ZN => n6749);
   U87349 : OAI22_X1 port map( A1 => n99080, A2 => n120496, B1 => n120722, B2 
                           => n120490, ZN => n6750);
   U87350 : OAI22_X1 port map( A1 => n99079, A2 => n120496, B1 => n120725, B2 
                           => n120490, ZN => n6751);
   U87351 : OAI22_X1 port map( A1 => n99078, A2 => n120496, B1 => n120728, B2 
                           => n120490, ZN => n6752);
   U87352 : OAI22_X1 port map( A1 => n99077, A2 => n120496, B1 => n120731, B2 
                           => n120490, ZN => n6753);
   U87353 : OAI22_X1 port map( A1 => n99076, A2 => n120497, B1 => n120734, B2 
                           => n120490, ZN => n6754);
   U87354 : OAI22_X1 port map( A1 => n99075, A2 => n120497, B1 => n120737, B2 
                           => n120491, ZN => n6755);
   U87355 : OAI22_X1 port map( A1 => n99074, A2 => n120497, B1 => n120740, B2 
                           => n120491, ZN => n6756);
   U87356 : OAI22_X1 port map( A1 => n99073, A2 => n120497, B1 => n120743, B2 
                           => n120491, ZN => n6757);
   U87357 : OAI22_X1 port map( A1 => n99072, A2 => n120497, B1 => n120746, B2 
                           => n120491, ZN => n6758);
   U87358 : OAI22_X1 port map( A1 => n99071, A2 => n120497, B1 => n120749, B2 
                           => n120491, ZN => n6759);
   U87359 : OAI22_X1 port map( A1 => n99070, A2 => n120497, B1 => n120752, B2 
                           => n120491, ZN => n6760);
   U87360 : OAI22_X1 port map( A1 => n99069, A2 => n120497, B1 => n120755, B2 
                           => n120491, ZN => n6761);
   U87361 : OAI22_X1 port map( A1 => n99068, A2 => n120497, B1 => n120758, B2 
                           => n120491, ZN => n6762);
   U87362 : OAI22_X1 port map( A1 => n99067, A2 => n120497, B1 => n120761, B2 
                           => n120491, ZN => n6763);
   U87363 : OAI22_X1 port map( A1 => n99066, A2 => n120497, B1 => n120764, B2 
                           => n120491, ZN => n6764);
   U87364 : OAI22_X1 port map( A1 => n99065, A2 => n120497, B1 => n120767, B2 
                           => n120491, ZN => n6765);
   U87365 : OAI22_X1 port map( A1 => n99064, A2 => n120498, B1 => n120770, B2 
                           => n120491, ZN => n6766);
   U87366 : OAI22_X1 port map( A1 => n99063, A2 => n120498, B1 => n120773, B2 
                           => n120492, ZN => n6767);
   U87367 : OAI22_X1 port map( A1 => n99062, A2 => n120498, B1 => n120776, B2 
                           => n120492, ZN => n6768);
   U87368 : OAI22_X1 port map( A1 => n99061, A2 => n120498, B1 => n120779, B2 
                           => n120492, ZN => n6769);
   U87369 : OAI22_X1 port map( A1 => n99060, A2 => n120498, B1 => n120782, B2 
                           => n120492, ZN => n6770);
   U87370 : OAI22_X1 port map( A1 => n99059, A2 => n120498, B1 => n120785, B2 
                           => n120492, ZN => n6771);
   U87371 : OAI22_X1 port map( A1 => n99058, A2 => n120498, B1 => n120788, B2 
                           => n120492, ZN => n6772);
   U87372 : OAI22_X1 port map( A1 => n99057, A2 => n120498, B1 => n120791, B2 
                           => n120492, ZN => n6773);
   U87373 : OAI22_X1 port map( A1 => n99056, A2 => n120498, B1 => n120794, B2 
                           => n120492, ZN => n6774);
   U87374 : OAI22_X1 port map( A1 => n99055, A2 => n120498, B1 => n120797, B2 
                           => n120492, ZN => n6775);
   U87375 : OAI22_X1 port map( A1 => n99054, A2 => n120498, B1 => n120800, B2 
                           => n120492, ZN => n6776);
   U87376 : OAI22_X1 port map( A1 => n99053, A2 => n120498, B1 => n120803, B2 
                           => n120492, ZN => n6777);
   U87377 : OAI22_X1 port map( A1 => n99052, A2 => n120499, B1 => n120806, B2 
                           => n120492, ZN => n6778);
   U87378 : OAI22_X1 port map( A1 => n99177, A2 => n120482, B1 => n120630, B2 
                           => n120476, ZN => n6655);
   U87379 : OAI22_X1 port map( A1 => n99176, A2 => n120482, B1 => n120633, B2 
                           => n120476, ZN => n6656);
   U87380 : OAI22_X1 port map( A1 => n99175, A2 => n120482, B1 => n120636, B2 
                           => n120476, ZN => n6657);
   U87381 : OAI22_X1 port map( A1 => n99174, A2 => n120482, B1 => n120639, B2 
                           => n120476, ZN => n6658);
   U87382 : OAI22_X1 port map( A1 => n99173, A2 => n120482, B1 => n120642, B2 
                           => n120476, ZN => n6659);
   U87383 : OAI22_X1 port map( A1 => n99172, A2 => n120482, B1 => n120645, B2 
                           => n120476, ZN => n6660);
   U87384 : OAI22_X1 port map( A1 => n99171, A2 => n120482, B1 => n120648, B2 
                           => n120476, ZN => n6661);
   U87385 : OAI22_X1 port map( A1 => n99170, A2 => n120482, B1 => n120651, B2 
                           => n120476, ZN => n6662);
   U87386 : OAI22_X1 port map( A1 => n99169, A2 => n120482, B1 => n120654, B2 
                           => n120476, ZN => n6663);
   U87387 : OAI22_X1 port map( A1 => n99168, A2 => n120482, B1 => n120657, B2 
                           => n120476, ZN => n6664);
   U87388 : OAI22_X1 port map( A1 => n99167, A2 => n120482, B1 => n120660, B2 
                           => n120476, ZN => n6665);
   U87389 : OAI22_X1 port map( A1 => n99166, A2 => n120483, B1 => n120663, B2 
                           => n120476, ZN => n6666);
   U87390 : OAI22_X1 port map( A1 => n99165, A2 => n120483, B1 => n120666, B2 
                           => n120477, ZN => n6667);
   U87391 : OAI22_X1 port map( A1 => n99164, A2 => n120483, B1 => n120669, B2 
                           => n120477, ZN => n6668);
   U87392 : OAI22_X1 port map( A1 => n99163, A2 => n120483, B1 => n120672, B2 
                           => n120477, ZN => n6669);
   U87393 : OAI22_X1 port map( A1 => n99162, A2 => n120483, B1 => n120675, B2 
                           => n120477, ZN => n6670);
   U87394 : OAI22_X1 port map( A1 => n99161, A2 => n120483, B1 => n120678, B2 
                           => n120477, ZN => n6671);
   U87395 : OAI22_X1 port map( A1 => n99160, A2 => n120483, B1 => n120681, B2 
                           => n120477, ZN => n6672);
   U87396 : OAI22_X1 port map( A1 => n99159, A2 => n120483, B1 => n120684, B2 
                           => n120477, ZN => n6673);
   U87397 : OAI22_X1 port map( A1 => n99158, A2 => n120483, B1 => n120687, B2 
                           => n120477, ZN => n6674);
   U87398 : OAI22_X1 port map( A1 => n99157, A2 => n120483, B1 => n120690, B2 
                           => n120477, ZN => n6675);
   U87399 : OAI22_X1 port map( A1 => n99156, A2 => n120483, B1 => n120693, B2 
                           => n120477, ZN => n6676);
   U87400 : OAI22_X1 port map( A1 => n99155, A2 => n120483, B1 => n120696, B2 
                           => n120477, ZN => n6677);
   U87401 : OAI22_X1 port map( A1 => n99154, A2 => n120484, B1 => n120699, B2 
                           => n120477, ZN => n6678);
   U87402 : OAI22_X1 port map( A1 => n99153, A2 => n120484, B1 => n120702, B2 
                           => n120478, ZN => n6679);
   U87403 : OAI22_X1 port map( A1 => n99152, A2 => n120484, B1 => n120705, B2 
                           => n120478, ZN => n6680);
   U87404 : OAI22_X1 port map( A1 => n99151, A2 => n120484, B1 => n120708, B2 
                           => n120478, ZN => n6681);
   U87405 : OAI22_X1 port map( A1 => n99150, A2 => n120484, B1 => n120711, B2 
                           => n120478, ZN => n6682);
   U87406 : OAI22_X1 port map( A1 => n99149, A2 => n120484, B1 => n120714, B2 
                           => n120478, ZN => n6683);
   U87407 : OAI22_X1 port map( A1 => n99148, A2 => n120484, B1 => n120717, B2 
                           => n120478, ZN => n6684);
   U87408 : OAI22_X1 port map( A1 => n99147, A2 => n120484, B1 => n120720, B2 
                           => n120478, ZN => n6685);
   U87409 : OAI22_X1 port map( A1 => n99146, A2 => n120484, B1 => n120723, B2 
                           => n120478, ZN => n6686);
   U87410 : OAI22_X1 port map( A1 => n99145, A2 => n120484, B1 => n120726, B2 
                           => n120478, ZN => n6687);
   U87411 : OAI22_X1 port map( A1 => n99144, A2 => n120484, B1 => n120729, B2 
                           => n120478, ZN => n6688);
   U87412 : OAI22_X1 port map( A1 => n99143, A2 => n120484, B1 => n120732, B2 
                           => n120478, ZN => n6689);
   U87413 : OAI22_X1 port map( A1 => n99142, A2 => n120485, B1 => n120735, B2 
                           => n120478, ZN => n6690);
   U87414 : OAI22_X1 port map( A1 => n99141, A2 => n120485, B1 => n120738, B2 
                           => n120479, ZN => n6691);
   U87415 : OAI22_X1 port map( A1 => n99140, A2 => n120485, B1 => n120741, B2 
                           => n120479, ZN => n6692);
   U87416 : OAI22_X1 port map( A1 => n99139, A2 => n120485, B1 => n120744, B2 
                           => n120479, ZN => n6693);
   U87417 : OAI22_X1 port map( A1 => n99138, A2 => n120485, B1 => n120747, B2 
                           => n120479, ZN => n6694);
   U87418 : OAI22_X1 port map( A1 => n99137, A2 => n120485, B1 => n120750, B2 
                           => n120479, ZN => n6695);
   U87419 : OAI22_X1 port map( A1 => n99136, A2 => n120485, B1 => n120753, B2 
                           => n120479, ZN => n6696);
   U87420 : OAI22_X1 port map( A1 => n99135, A2 => n120485, B1 => n120756, B2 
                           => n120479, ZN => n6697);
   U87421 : OAI22_X1 port map( A1 => n99134, A2 => n120485, B1 => n120759, B2 
                           => n120479, ZN => n6698);
   U87422 : OAI22_X1 port map( A1 => n99133, A2 => n120485, B1 => n120762, B2 
                           => n120479, ZN => n6699);
   U87423 : OAI22_X1 port map( A1 => n99132, A2 => n120485, B1 => n120765, B2 
                           => n120479, ZN => n6700);
   U87424 : OAI22_X1 port map( A1 => n99131, A2 => n120485, B1 => n120768, B2 
                           => n120479, ZN => n6701);
   U87425 : OAI22_X1 port map( A1 => n99130, A2 => n120486, B1 => n120771, B2 
                           => n120479, ZN => n6702);
   U87426 : OAI22_X1 port map( A1 => n99129, A2 => n120486, B1 => n120774, B2 
                           => n120480, ZN => n6703);
   U87427 : OAI22_X1 port map( A1 => n99128, A2 => n120486, B1 => n120777, B2 
                           => n120480, ZN => n6704);
   U87428 : OAI22_X1 port map( A1 => n99127, A2 => n120486, B1 => n120780, B2 
                           => n120480, ZN => n6705);
   U87429 : OAI22_X1 port map( A1 => n99126, A2 => n120486, B1 => n120783, B2 
                           => n120480, ZN => n6706);
   U87430 : OAI22_X1 port map( A1 => n99125, A2 => n120486, B1 => n120786, B2 
                           => n120480, ZN => n6707);
   U87431 : OAI22_X1 port map( A1 => n99124, A2 => n120486, B1 => n120789, B2 
                           => n120480, ZN => n6708);
   U87432 : OAI22_X1 port map( A1 => n99123, A2 => n120486, B1 => n120792, B2 
                           => n120480, ZN => n6709);
   U87433 : OAI22_X1 port map( A1 => n99122, A2 => n120486, B1 => n120795, B2 
                           => n120480, ZN => n6710);
   U87434 : OAI22_X1 port map( A1 => n99121, A2 => n120486, B1 => n120798, B2 
                           => n120480, ZN => n6711);
   U87435 : OAI22_X1 port map( A1 => n99120, A2 => n120486, B1 => n120801, B2 
                           => n120480, ZN => n6712);
   U87436 : OAI22_X1 port map( A1 => n99119, A2 => n120486, B1 => n120804, B2 
                           => n120480, ZN => n6713);
   U87437 : OAI22_X1 port map( A1 => n99118, A2 => n120487, B1 => n120807, B2 
                           => n120480, ZN => n6714);
   U87438 : OAI22_X1 port map( A1 => n99309, A2 => n120458, B1 => n120630, B2 
                           => n120452, ZN => n6527);
   U87439 : OAI22_X1 port map( A1 => n99308, A2 => n120458, B1 => n120633, B2 
                           => n120452, ZN => n6528);
   U87440 : OAI22_X1 port map( A1 => n99307, A2 => n120458, B1 => n120636, B2 
                           => n120452, ZN => n6529);
   U87441 : OAI22_X1 port map( A1 => n99306, A2 => n120458, B1 => n120639, B2 
                           => n120452, ZN => n6530);
   U87442 : OAI22_X1 port map( A1 => n99305, A2 => n120458, B1 => n120642, B2 
                           => n120452, ZN => n6531);
   U87443 : OAI22_X1 port map( A1 => n99304, A2 => n120458, B1 => n120645, B2 
                           => n120452, ZN => n6532);
   U87444 : OAI22_X1 port map( A1 => n99303, A2 => n120458, B1 => n120648, B2 
                           => n120452, ZN => n6533);
   U87445 : OAI22_X1 port map( A1 => n99302, A2 => n120458, B1 => n120651, B2 
                           => n120452, ZN => n6534);
   U87446 : OAI22_X1 port map( A1 => n99301, A2 => n120458, B1 => n120654, B2 
                           => n120452, ZN => n6535);
   U87447 : OAI22_X1 port map( A1 => n99300, A2 => n120458, B1 => n120657, B2 
                           => n120452, ZN => n6536);
   U87448 : OAI22_X1 port map( A1 => n99299, A2 => n120458, B1 => n120660, B2 
                           => n120452, ZN => n6537);
   U87449 : OAI22_X1 port map( A1 => n99298, A2 => n120459, B1 => n120663, B2 
                           => n120452, ZN => n6538);
   U87450 : OAI22_X1 port map( A1 => n99297, A2 => n120459, B1 => n120666, B2 
                           => n120453, ZN => n6539);
   U87451 : OAI22_X1 port map( A1 => n99296, A2 => n120459, B1 => n120669, B2 
                           => n120453, ZN => n6540);
   U87452 : OAI22_X1 port map( A1 => n99295, A2 => n120459, B1 => n120672, B2 
                           => n120453, ZN => n6541);
   U87453 : OAI22_X1 port map( A1 => n99294, A2 => n120459, B1 => n120675, B2 
                           => n120453, ZN => n6542);
   U87454 : OAI22_X1 port map( A1 => n99293, A2 => n120459, B1 => n120678, B2 
                           => n120453, ZN => n6543);
   U87455 : OAI22_X1 port map( A1 => n99292, A2 => n120459, B1 => n120681, B2 
                           => n120453, ZN => n6544);
   U87456 : OAI22_X1 port map( A1 => n99291, A2 => n120459, B1 => n120684, B2 
                           => n120453, ZN => n6545);
   U87457 : OAI22_X1 port map( A1 => n99290, A2 => n120459, B1 => n120687, B2 
                           => n120453, ZN => n6546);
   U87458 : OAI22_X1 port map( A1 => n99289, A2 => n120459, B1 => n120690, B2 
                           => n120453, ZN => n6547);
   U87459 : OAI22_X1 port map( A1 => n99288, A2 => n120459, B1 => n120693, B2 
                           => n120453, ZN => n6548);
   U87460 : OAI22_X1 port map( A1 => n99287, A2 => n120459, B1 => n120696, B2 
                           => n120453, ZN => n6549);
   U87461 : OAI22_X1 port map( A1 => n99286, A2 => n120460, B1 => n120699, B2 
                           => n120453, ZN => n6550);
   U87462 : OAI22_X1 port map( A1 => n99285, A2 => n120460, B1 => n120702, B2 
                           => n120454, ZN => n6551);
   U87463 : OAI22_X1 port map( A1 => n99284, A2 => n120460, B1 => n120705, B2 
                           => n120454, ZN => n6552);
   U87464 : OAI22_X1 port map( A1 => n99283, A2 => n120460, B1 => n120708, B2 
                           => n120454, ZN => n6553);
   U87465 : OAI22_X1 port map( A1 => n99282, A2 => n120460, B1 => n120711, B2 
                           => n120454, ZN => n6554);
   U87466 : OAI22_X1 port map( A1 => n99281, A2 => n120460, B1 => n120714, B2 
                           => n120454, ZN => n6555);
   U87467 : OAI22_X1 port map( A1 => n99280, A2 => n120460, B1 => n120717, B2 
                           => n120454, ZN => n6556);
   U87468 : OAI22_X1 port map( A1 => n99279, A2 => n120460, B1 => n120720, B2 
                           => n120454, ZN => n6557);
   U87469 : OAI22_X1 port map( A1 => n99278, A2 => n120460, B1 => n120723, B2 
                           => n120454, ZN => n6558);
   U87470 : OAI22_X1 port map( A1 => n99277, A2 => n120460, B1 => n120726, B2 
                           => n120454, ZN => n6559);
   U87471 : OAI22_X1 port map( A1 => n99276, A2 => n120460, B1 => n120729, B2 
                           => n120454, ZN => n6560);
   U87472 : OAI22_X1 port map( A1 => n99275, A2 => n120460, B1 => n120732, B2 
                           => n120454, ZN => n6561);
   U87473 : OAI22_X1 port map( A1 => n99274, A2 => n120461, B1 => n120735, B2 
                           => n120454, ZN => n6562);
   U87474 : OAI22_X1 port map( A1 => n99273, A2 => n120461, B1 => n120738, B2 
                           => n120455, ZN => n6563);
   U87475 : OAI22_X1 port map( A1 => n99272, A2 => n120461, B1 => n120741, B2 
                           => n120455, ZN => n6564);
   U87476 : OAI22_X1 port map( A1 => n99271, A2 => n120461, B1 => n120744, B2 
                           => n120455, ZN => n6565);
   U87477 : OAI22_X1 port map( A1 => n99270, A2 => n120461, B1 => n120747, B2 
                           => n120455, ZN => n6566);
   U87478 : OAI22_X1 port map( A1 => n99269, A2 => n120461, B1 => n120750, B2 
                           => n120455, ZN => n6567);
   U87479 : OAI22_X1 port map( A1 => n99268, A2 => n120461, B1 => n120753, B2 
                           => n120455, ZN => n6568);
   U87480 : OAI22_X1 port map( A1 => n99267, A2 => n120461, B1 => n120756, B2 
                           => n120455, ZN => n6569);
   U87481 : OAI22_X1 port map( A1 => n99266, A2 => n120461, B1 => n120759, B2 
                           => n120455, ZN => n6570);
   U87482 : OAI22_X1 port map( A1 => n99265, A2 => n120461, B1 => n120762, B2 
                           => n120455, ZN => n6571);
   U87483 : OAI22_X1 port map( A1 => n99264, A2 => n120461, B1 => n120765, B2 
                           => n120455, ZN => n6572);
   U87484 : OAI22_X1 port map( A1 => n99263, A2 => n120461, B1 => n120768, B2 
                           => n120455, ZN => n6573);
   U87485 : OAI22_X1 port map( A1 => n99262, A2 => n120462, B1 => n120771, B2 
                           => n120455, ZN => n6574);
   U87486 : OAI22_X1 port map( A1 => n99261, A2 => n120462, B1 => n120774, B2 
                           => n120456, ZN => n6575);
   U87487 : OAI22_X1 port map( A1 => n99260, A2 => n120462, B1 => n120777, B2 
                           => n120456, ZN => n6576);
   U87488 : OAI22_X1 port map( A1 => n99259, A2 => n120462, B1 => n120780, B2 
                           => n120456, ZN => n6577);
   U87489 : OAI22_X1 port map( A1 => n99258, A2 => n120462, B1 => n120783, B2 
                           => n120456, ZN => n6578);
   U87490 : OAI22_X1 port map( A1 => n99257, A2 => n120462, B1 => n120786, B2 
                           => n120456, ZN => n6579);
   U87491 : OAI22_X1 port map( A1 => n99256, A2 => n120462, B1 => n120789, B2 
                           => n120456, ZN => n6580);
   U87492 : OAI22_X1 port map( A1 => n99255, A2 => n120462, B1 => n120792, B2 
                           => n120456, ZN => n6581);
   U87493 : OAI22_X1 port map( A1 => n99254, A2 => n120462, B1 => n120795, B2 
                           => n120456, ZN => n6582);
   U87494 : OAI22_X1 port map( A1 => n99253, A2 => n120462, B1 => n120798, B2 
                           => n120456, ZN => n6583);
   U87495 : OAI22_X1 port map( A1 => n99252, A2 => n120462, B1 => n120801, B2 
                           => n120456, ZN => n6584);
   U87496 : OAI22_X1 port map( A1 => n99251, A2 => n120462, B1 => n120804, B2 
                           => n120456, ZN => n6585);
   U87497 : OAI22_X1 port map( A1 => n99250, A2 => n120463, B1 => n120807, B2 
                           => n120456, ZN => n6586);
   U87498 : OAI22_X1 port map( A1 => n98778, A2 => n120581, B1 => n120629, B2 
                           => n120575, ZN => n7167);
   U87499 : OAI22_X1 port map( A1 => n98777, A2 => n120581, B1 => n120632, B2 
                           => n120575, ZN => n7168);
   U87500 : OAI22_X1 port map( A1 => n98776, A2 => n120581, B1 => n120635, B2 
                           => n120575, ZN => n7169);
   U87501 : OAI22_X1 port map( A1 => n98775, A2 => n120581, B1 => n120638, B2 
                           => n120575, ZN => n7170);
   U87502 : OAI22_X1 port map( A1 => n98774, A2 => n120581, B1 => n120641, B2 
                           => n120575, ZN => n7171);
   U87503 : OAI22_X1 port map( A1 => n98773, A2 => n120581, B1 => n120644, B2 
                           => n120575, ZN => n7172);
   U87504 : OAI22_X1 port map( A1 => n98772, A2 => n120581, B1 => n120647, B2 
                           => n120575, ZN => n7173);
   U87505 : OAI22_X1 port map( A1 => n98771, A2 => n120581, B1 => n120650, B2 
                           => n120575, ZN => n7174);
   U87506 : OAI22_X1 port map( A1 => n98770, A2 => n120581, B1 => n120653, B2 
                           => n120575, ZN => n7175);
   U87507 : OAI22_X1 port map( A1 => n98769, A2 => n120581, B1 => n120656, B2 
                           => n120575, ZN => n7176);
   U87508 : OAI22_X1 port map( A1 => n98768, A2 => n120581, B1 => n120659, B2 
                           => n120575, ZN => n7177);
   U87509 : OAI22_X1 port map( A1 => n98767, A2 => n120582, B1 => n120662, B2 
                           => n120575, ZN => n7178);
   U87510 : OAI22_X1 port map( A1 => n98766, A2 => n120582, B1 => n120665, B2 
                           => n120576, ZN => n7179);
   U87511 : OAI22_X1 port map( A1 => n98765, A2 => n120582, B1 => n120668, B2 
                           => n120576, ZN => n7180);
   U87512 : OAI22_X1 port map( A1 => n98764, A2 => n120582, B1 => n120671, B2 
                           => n120576, ZN => n7181);
   U87513 : OAI22_X1 port map( A1 => n98763, A2 => n120582, B1 => n120674, B2 
                           => n120576, ZN => n7182);
   U87514 : OAI22_X1 port map( A1 => n98762, A2 => n120582, B1 => n120677, B2 
                           => n120576, ZN => n7183);
   U87515 : OAI22_X1 port map( A1 => n98761, A2 => n120582, B1 => n120680, B2 
                           => n120576, ZN => n7184);
   U87516 : OAI22_X1 port map( A1 => n98760, A2 => n120582, B1 => n120683, B2 
                           => n120576, ZN => n7185);
   U87517 : OAI22_X1 port map( A1 => n98759, A2 => n120582, B1 => n120686, B2 
                           => n120576, ZN => n7186);
   U87518 : OAI22_X1 port map( A1 => n98758, A2 => n120582, B1 => n120689, B2 
                           => n120576, ZN => n7187);
   U87519 : OAI22_X1 port map( A1 => n98757, A2 => n120582, B1 => n120692, B2 
                           => n120576, ZN => n7188);
   U87520 : OAI22_X1 port map( A1 => n98756, A2 => n120582, B1 => n120695, B2 
                           => n120576, ZN => n7189);
   U87521 : OAI22_X1 port map( A1 => n98755, A2 => n120583, B1 => n120698, B2 
                           => n120576, ZN => n7190);
   U87522 : OAI22_X1 port map( A1 => n98754, A2 => n120583, B1 => n120701, B2 
                           => n120577, ZN => n7191);
   U87523 : OAI22_X1 port map( A1 => n98753, A2 => n120583, B1 => n120704, B2 
                           => n120577, ZN => n7192);
   U87524 : OAI22_X1 port map( A1 => n98752, A2 => n120583, B1 => n120707, B2 
                           => n120577, ZN => n7193);
   U87525 : OAI22_X1 port map( A1 => n98751, A2 => n120583, B1 => n120710, B2 
                           => n120577, ZN => n7194);
   U87526 : OAI22_X1 port map( A1 => n98750, A2 => n120583, B1 => n120713, B2 
                           => n120577, ZN => n7195);
   U87527 : OAI22_X1 port map( A1 => n98749, A2 => n120583, B1 => n120716, B2 
                           => n120577, ZN => n7196);
   U87528 : OAI22_X1 port map( A1 => n98748, A2 => n120583, B1 => n120719, B2 
                           => n120577, ZN => n7197);
   U87529 : OAI22_X1 port map( A1 => n98747, A2 => n120583, B1 => n120722, B2 
                           => n120577, ZN => n7198);
   U87530 : OAI22_X1 port map( A1 => n98746, A2 => n120583, B1 => n120725, B2 
                           => n120577, ZN => n7199);
   U87531 : OAI22_X1 port map( A1 => n98745, A2 => n120583, B1 => n120728, B2 
                           => n120577, ZN => n7200);
   U87532 : OAI22_X1 port map( A1 => n98744, A2 => n120583, B1 => n120731, B2 
                           => n120577, ZN => n7201);
   U87533 : OAI22_X1 port map( A1 => n98743, A2 => n120584, B1 => n120734, B2 
                           => n120577, ZN => n7202);
   U87534 : OAI22_X1 port map( A1 => n98742, A2 => n120584, B1 => n120737, B2 
                           => n120578, ZN => n7203);
   U87535 : OAI22_X1 port map( A1 => n98741, A2 => n120584, B1 => n120740, B2 
                           => n120578, ZN => n7204);
   U87536 : OAI22_X1 port map( A1 => n98740, A2 => n120584, B1 => n120743, B2 
                           => n120578, ZN => n7205);
   U87537 : OAI22_X1 port map( A1 => n98739, A2 => n120584, B1 => n120746, B2 
                           => n120578, ZN => n7206);
   U87538 : OAI22_X1 port map( A1 => n98738, A2 => n120584, B1 => n120749, B2 
                           => n120578, ZN => n7207);
   U87539 : OAI22_X1 port map( A1 => n98737, A2 => n120584, B1 => n120752, B2 
                           => n120578, ZN => n7208);
   U87540 : OAI22_X1 port map( A1 => n98736, A2 => n120584, B1 => n120755, B2 
                           => n120578, ZN => n7209);
   U87541 : OAI22_X1 port map( A1 => n98735, A2 => n120584, B1 => n120758, B2 
                           => n120578, ZN => n7210);
   U87542 : OAI22_X1 port map( A1 => n98734, A2 => n120584, B1 => n120761, B2 
                           => n120578, ZN => n7211);
   U87543 : OAI22_X1 port map( A1 => n98733, A2 => n120584, B1 => n120764, B2 
                           => n120578, ZN => n7212);
   U87544 : OAI22_X1 port map( A1 => n98732, A2 => n120584, B1 => n120767, B2 
                           => n120578, ZN => n7213);
   U87545 : OAI22_X1 port map( A1 => n98731, A2 => n120585, B1 => n120770, B2 
                           => n120578, ZN => n7214);
   U87546 : OAI22_X1 port map( A1 => n98730, A2 => n120585, B1 => n120773, B2 
                           => n120579, ZN => n7215);
   U87547 : OAI22_X1 port map( A1 => n98729, A2 => n120585, B1 => n120776, B2 
                           => n120579, ZN => n7216);
   U87548 : OAI22_X1 port map( A1 => n98728, A2 => n120585, B1 => n120779, B2 
                           => n120579, ZN => n7217);
   U87549 : OAI22_X1 port map( A1 => n98727, A2 => n120585, B1 => n120782, B2 
                           => n120579, ZN => n7218);
   U87550 : OAI22_X1 port map( A1 => n98726, A2 => n120585, B1 => n120785, B2 
                           => n120579, ZN => n7219);
   U87551 : OAI22_X1 port map( A1 => n98725, A2 => n120585, B1 => n120788, B2 
                           => n120579, ZN => n7220);
   U87552 : OAI22_X1 port map( A1 => n98724, A2 => n120585, B1 => n120791, B2 
                           => n120579, ZN => n7221);
   U87553 : OAI22_X1 port map( A1 => n98723, A2 => n120585, B1 => n120794, B2 
                           => n120579, ZN => n7222);
   U87554 : OAI22_X1 port map( A1 => n98722, A2 => n120585, B1 => n120797, B2 
                           => n120579, ZN => n7223);
   U87555 : OAI22_X1 port map( A1 => n98721, A2 => n120585, B1 => n120800, B2 
                           => n120579, ZN => n7224);
   U87556 : OAI22_X1 port map( A1 => n98720, A2 => n120585, B1 => n120803, B2 
                           => n120579, ZN => n7225);
   U87557 : OAI22_X1 port map( A1 => n98719, A2 => n120586, B1 => n120806, B2 
                           => n120579, ZN => n7226);
   U87558 : OAI22_X1 port map( A1 => n99045, A2 => n120506, B1 => n120629, B2 
                           => n120500, ZN => n6783);
   U87559 : OAI22_X1 port map( A1 => n99044, A2 => n120506, B1 => n120632, B2 
                           => n120500, ZN => n6784);
   U87560 : OAI22_X1 port map( A1 => n99043, A2 => n120506, B1 => n120635, B2 
                           => n120500, ZN => n6785);
   U87561 : OAI22_X1 port map( A1 => n99042, A2 => n120506, B1 => n120638, B2 
                           => n120500, ZN => n6786);
   U87562 : OAI22_X1 port map( A1 => n99041, A2 => n120506, B1 => n120641, B2 
                           => n120500, ZN => n6787);
   U87563 : OAI22_X1 port map( A1 => n99040, A2 => n120506, B1 => n120644, B2 
                           => n120500, ZN => n6788);
   U87564 : OAI22_X1 port map( A1 => n99039, A2 => n120506, B1 => n120647, B2 
                           => n120500, ZN => n6789);
   U87565 : OAI22_X1 port map( A1 => n99038, A2 => n120506, B1 => n120650, B2 
                           => n120500, ZN => n6790);
   U87566 : OAI22_X1 port map( A1 => n99037, A2 => n120506, B1 => n120653, B2 
                           => n120500, ZN => n6791);
   U87567 : OAI22_X1 port map( A1 => n99036, A2 => n120506, B1 => n120656, B2 
                           => n120500, ZN => n6792);
   U87568 : OAI22_X1 port map( A1 => n99035, A2 => n120506, B1 => n120659, B2 
                           => n120500, ZN => n6793);
   U87569 : OAI22_X1 port map( A1 => n99034, A2 => n120507, B1 => n120662, B2 
                           => n120500, ZN => n6794);
   U87570 : OAI22_X1 port map( A1 => n99033, A2 => n120507, B1 => n120665, B2 
                           => n120501, ZN => n6795);
   U87571 : OAI22_X1 port map( A1 => n99032, A2 => n120507, B1 => n120668, B2 
                           => n120501, ZN => n6796);
   U87572 : OAI22_X1 port map( A1 => n99031, A2 => n120507, B1 => n120671, B2 
                           => n120501, ZN => n6797);
   U87573 : OAI22_X1 port map( A1 => n99030, A2 => n120507, B1 => n120674, B2 
                           => n120501, ZN => n6798);
   U87574 : OAI22_X1 port map( A1 => n99029, A2 => n120507, B1 => n120677, B2 
                           => n120501, ZN => n6799);
   U87575 : OAI22_X1 port map( A1 => n99028, A2 => n120507, B1 => n120680, B2 
                           => n120501, ZN => n6800);
   U87576 : OAI22_X1 port map( A1 => n99027, A2 => n120507, B1 => n120683, B2 
                           => n120501, ZN => n6801);
   U87577 : OAI22_X1 port map( A1 => n99026, A2 => n120507, B1 => n120686, B2 
                           => n120501, ZN => n6802);
   U87578 : OAI22_X1 port map( A1 => n99025, A2 => n120507, B1 => n120689, B2 
                           => n120501, ZN => n6803);
   U87579 : OAI22_X1 port map( A1 => n99024, A2 => n120507, B1 => n120692, B2 
                           => n120501, ZN => n6804);
   U87580 : OAI22_X1 port map( A1 => n99023, A2 => n120507, B1 => n120695, B2 
                           => n120501, ZN => n6805);
   U87581 : OAI22_X1 port map( A1 => n99022, A2 => n120508, B1 => n120698, B2 
                           => n120501, ZN => n6806);
   U87582 : OAI22_X1 port map( A1 => n99021, A2 => n120508, B1 => n120701, B2 
                           => n120502, ZN => n6807);
   U87583 : OAI22_X1 port map( A1 => n99020, A2 => n120508, B1 => n120704, B2 
                           => n120502, ZN => n6808);
   U87584 : OAI22_X1 port map( A1 => n99019, A2 => n120508, B1 => n120707, B2 
                           => n120502, ZN => n6809);
   U87585 : OAI22_X1 port map( A1 => n99018, A2 => n120508, B1 => n120710, B2 
                           => n120502, ZN => n6810);
   U87586 : OAI22_X1 port map( A1 => n99017, A2 => n120508, B1 => n120713, B2 
                           => n120502, ZN => n6811);
   U87587 : OAI22_X1 port map( A1 => n99016, A2 => n120508, B1 => n120716, B2 
                           => n120502, ZN => n6812);
   U87588 : OAI22_X1 port map( A1 => n99015, A2 => n120508, B1 => n120719, B2 
                           => n120502, ZN => n6813);
   U87589 : OAI22_X1 port map( A1 => n99014, A2 => n120508, B1 => n120722, B2 
                           => n120502, ZN => n6814);
   U87590 : OAI22_X1 port map( A1 => n99013, A2 => n120508, B1 => n120725, B2 
                           => n120502, ZN => n6815);
   U87591 : OAI22_X1 port map( A1 => n99012, A2 => n120508, B1 => n120728, B2 
                           => n120502, ZN => n6816);
   U87592 : OAI22_X1 port map( A1 => n99011, A2 => n120508, B1 => n120731, B2 
                           => n120502, ZN => n6817);
   U87593 : OAI22_X1 port map( A1 => n99010, A2 => n120509, B1 => n120734, B2 
                           => n120502, ZN => n6818);
   U87594 : OAI22_X1 port map( A1 => n99009, A2 => n120509, B1 => n120737, B2 
                           => n120503, ZN => n6819);
   U87595 : OAI22_X1 port map( A1 => n99008, A2 => n120509, B1 => n120740, B2 
                           => n120503, ZN => n6820);
   U87596 : OAI22_X1 port map( A1 => n99007, A2 => n120509, B1 => n120743, B2 
                           => n120503, ZN => n6821);
   U87597 : OAI22_X1 port map( A1 => n99006, A2 => n120509, B1 => n120746, B2 
                           => n120503, ZN => n6822);
   U87598 : OAI22_X1 port map( A1 => n99005, A2 => n120509, B1 => n120749, B2 
                           => n120503, ZN => n6823);
   U87599 : OAI22_X1 port map( A1 => n99004, A2 => n120509, B1 => n120752, B2 
                           => n120503, ZN => n6824);
   U87600 : OAI22_X1 port map( A1 => n99003, A2 => n120509, B1 => n120755, B2 
                           => n120503, ZN => n6825);
   U87601 : OAI22_X1 port map( A1 => n99002, A2 => n120509, B1 => n120758, B2 
                           => n120503, ZN => n6826);
   U87602 : OAI22_X1 port map( A1 => n99001, A2 => n120509, B1 => n120761, B2 
                           => n120503, ZN => n6827);
   U87603 : OAI22_X1 port map( A1 => n99000, A2 => n120509, B1 => n120764, B2 
                           => n120503, ZN => n6828);
   U87604 : OAI22_X1 port map( A1 => n98999, A2 => n120509, B1 => n120767, B2 
                           => n120503, ZN => n6829);
   U87605 : OAI22_X1 port map( A1 => n98998, A2 => n120510, B1 => n120770, B2 
                           => n120503, ZN => n6830);
   U87606 : OAI22_X1 port map( A1 => n98997, A2 => n120510, B1 => n120773, B2 
                           => n120504, ZN => n6831);
   U87607 : OAI22_X1 port map( A1 => n98996, A2 => n120510, B1 => n120776, B2 
                           => n120504, ZN => n6832);
   U87608 : OAI22_X1 port map( A1 => n98995, A2 => n120510, B1 => n120779, B2 
                           => n120504, ZN => n6833);
   U87609 : OAI22_X1 port map( A1 => n98994, A2 => n120510, B1 => n120782, B2 
                           => n120504, ZN => n6834);
   U87610 : OAI22_X1 port map( A1 => n98993, A2 => n120510, B1 => n120785, B2 
                           => n120504, ZN => n6835);
   U87611 : OAI22_X1 port map( A1 => n98992, A2 => n120510, B1 => n120788, B2 
                           => n120504, ZN => n6836);
   U87612 : OAI22_X1 port map( A1 => n98991, A2 => n120510, B1 => n120791, B2 
                           => n120504, ZN => n6837);
   U87613 : OAI22_X1 port map( A1 => n98990, A2 => n120510, B1 => n120794, B2 
                           => n120504, ZN => n6838);
   U87614 : OAI22_X1 port map( A1 => n98989, A2 => n120510, B1 => n120797, B2 
                           => n120504, ZN => n6839);
   U87615 : OAI22_X1 port map( A1 => n98988, A2 => n120510, B1 => n120800, B2 
                           => n120504, ZN => n6840);
   U87616 : OAI22_X1 port map( A1 => n98987, A2 => n120510, B1 => n120803, B2 
                           => n120504, ZN => n6841);
   U87617 : OAI22_X1 port map( A1 => n98986, A2 => n120511, B1 => n120806, B2 
                           => n120504, ZN => n6842);
   U87618 : OAI22_X1 port map( A1 => n98907, A2 => n120556, B1 => n120629, B2 
                           => n120550, ZN => n7039);
   U87619 : OAI22_X1 port map( A1 => n98906, A2 => n120556, B1 => n120632, B2 
                           => n120550, ZN => n7040);
   U87620 : OAI22_X1 port map( A1 => n98905, A2 => n120556, B1 => n120635, B2 
                           => n120550, ZN => n7041);
   U87621 : OAI22_X1 port map( A1 => n98904, A2 => n120556, B1 => n120638, B2 
                           => n120550, ZN => n7042);
   U87622 : OAI22_X1 port map( A1 => n98903, A2 => n120556, B1 => n120641, B2 
                           => n120550, ZN => n7043);
   U87623 : OAI22_X1 port map( A1 => n98902, A2 => n120556, B1 => n120644, B2 
                           => n120550, ZN => n7044);
   U87624 : OAI22_X1 port map( A1 => n98901, A2 => n120556, B1 => n120647, B2 
                           => n120550, ZN => n7045);
   U87625 : OAI22_X1 port map( A1 => n98900, A2 => n120556, B1 => n120650, B2 
                           => n120550, ZN => n7046);
   U87626 : OAI22_X1 port map( A1 => n98899, A2 => n120556, B1 => n120653, B2 
                           => n120550, ZN => n7047);
   U87627 : OAI22_X1 port map( A1 => n98898, A2 => n120556, B1 => n120656, B2 
                           => n120550, ZN => n7048);
   U87628 : OAI22_X1 port map( A1 => n98897, A2 => n120556, B1 => n120659, B2 
                           => n120550, ZN => n7049);
   U87629 : OAI22_X1 port map( A1 => n98896, A2 => n120557, B1 => n120662, B2 
                           => n120550, ZN => n7050);
   U87630 : OAI22_X1 port map( A1 => n98895, A2 => n120557, B1 => n120665, B2 
                           => n120551, ZN => n7051);
   U87631 : OAI22_X1 port map( A1 => n98894, A2 => n120557, B1 => n120668, B2 
                           => n120551, ZN => n7052);
   U87632 : OAI22_X1 port map( A1 => n98893, A2 => n120557, B1 => n120671, B2 
                           => n120551, ZN => n7053);
   U87633 : OAI22_X1 port map( A1 => n98892, A2 => n120557, B1 => n120674, B2 
                           => n120551, ZN => n7054);
   U87634 : OAI22_X1 port map( A1 => n98891, A2 => n120557, B1 => n120677, B2 
                           => n120551, ZN => n7055);
   U87635 : OAI22_X1 port map( A1 => n98890, A2 => n120557, B1 => n120680, B2 
                           => n120551, ZN => n7056);
   U87636 : OAI22_X1 port map( A1 => n98889, A2 => n120557, B1 => n120683, B2 
                           => n120551, ZN => n7057);
   U87637 : OAI22_X1 port map( A1 => n98888, A2 => n120557, B1 => n120686, B2 
                           => n120551, ZN => n7058);
   U87638 : OAI22_X1 port map( A1 => n98887, A2 => n120557, B1 => n120689, B2 
                           => n120551, ZN => n7059);
   U87639 : OAI22_X1 port map( A1 => n98886, A2 => n120557, B1 => n120692, B2 
                           => n120551, ZN => n7060);
   U87640 : OAI22_X1 port map( A1 => n98885, A2 => n120557, B1 => n120695, B2 
                           => n120551, ZN => n7061);
   U87641 : OAI22_X1 port map( A1 => n98884, A2 => n120558, B1 => n120698, B2 
                           => n120551, ZN => n7062);
   U87642 : OAI22_X1 port map( A1 => n98883, A2 => n120558, B1 => n120701, B2 
                           => n120552, ZN => n7063);
   U87643 : OAI22_X1 port map( A1 => n98882, A2 => n120558, B1 => n120704, B2 
                           => n120552, ZN => n7064);
   U87644 : OAI22_X1 port map( A1 => n98881, A2 => n120558, B1 => n120707, B2 
                           => n120552, ZN => n7065);
   U87645 : OAI22_X1 port map( A1 => n98880, A2 => n120558, B1 => n120710, B2 
                           => n120552, ZN => n7066);
   U87646 : OAI22_X1 port map( A1 => n98879, A2 => n120558, B1 => n120713, B2 
                           => n120552, ZN => n7067);
   U87647 : OAI22_X1 port map( A1 => n98878, A2 => n120558, B1 => n120716, B2 
                           => n120552, ZN => n7068);
   U87648 : OAI22_X1 port map( A1 => n98877, A2 => n120558, B1 => n120719, B2 
                           => n120552, ZN => n7069);
   U87649 : OAI22_X1 port map( A1 => n98876, A2 => n120558, B1 => n120722, B2 
                           => n120552, ZN => n7070);
   U87650 : OAI22_X1 port map( A1 => n98875, A2 => n120558, B1 => n120725, B2 
                           => n120552, ZN => n7071);
   U87651 : OAI22_X1 port map( A1 => n98874, A2 => n120558, B1 => n120728, B2 
                           => n120552, ZN => n7072);
   U87652 : OAI22_X1 port map( A1 => n98873, A2 => n120558, B1 => n120731, B2 
                           => n120552, ZN => n7073);
   U87653 : OAI22_X1 port map( A1 => n98872, A2 => n120559, B1 => n120734, B2 
                           => n120552, ZN => n7074);
   U87654 : OAI22_X1 port map( A1 => n98871, A2 => n120559, B1 => n120737, B2 
                           => n120553, ZN => n7075);
   U87655 : OAI22_X1 port map( A1 => n98870, A2 => n120559, B1 => n120740, B2 
                           => n120553, ZN => n7076);
   U87656 : OAI22_X1 port map( A1 => n98869, A2 => n120559, B1 => n120743, B2 
                           => n120553, ZN => n7077);
   U87657 : OAI22_X1 port map( A1 => n98868, A2 => n120559, B1 => n120746, B2 
                           => n120553, ZN => n7078);
   U87658 : OAI22_X1 port map( A1 => n98867, A2 => n120559, B1 => n120749, B2 
                           => n120553, ZN => n7079);
   U87659 : OAI22_X1 port map( A1 => n98866, A2 => n120559, B1 => n120752, B2 
                           => n120553, ZN => n7080);
   U87660 : OAI22_X1 port map( A1 => n98865, A2 => n120559, B1 => n120755, B2 
                           => n120553, ZN => n7081);
   U87661 : OAI22_X1 port map( A1 => n98864, A2 => n120559, B1 => n120758, B2 
                           => n120553, ZN => n7082);
   U87662 : OAI22_X1 port map( A1 => n98863, A2 => n120559, B1 => n120761, B2 
                           => n120553, ZN => n7083);
   U87663 : OAI22_X1 port map( A1 => n98862, A2 => n120559, B1 => n120764, B2 
                           => n120553, ZN => n7084);
   U87664 : OAI22_X1 port map( A1 => n98861, A2 => n120559, B1 => n120767, B2 
                           => n120553, ZN => n7085);
   U87665 : OAI22_X1 port map( A1 => n98860, A2 => n120560, B1 => n120770, B2 
                           => n120553, ZN => n7086);
   U87666 : OAI22_X1 port map( A1 => n98859, A2 => n120560, B1 => n120773, B2 
                           => n120554, ZN => n7087);
   U87667 : OAI22_X1 port map( A1 => n98858, A2 => n120560, B1 => n120776, B2 
                           => n120554, ZN => n7088);
   U87668 : OAI22_X1 port map( A1 => n98857, A2 => n120560, B1 => n120779, B2 
                           => n120554, ZN => n7089);
   U87669 : OAI22_X1 port map( A1 => n98856, A2 => n120560, B1 => n120782, B2 
                           => n120554, ZN => n7090);
   U87670 : OAI22_X1 port map( A1 => n98855, A2 => n120560, B1 => n120785, B2 
                           => n120554, ZN => n7091);
   U87671 : OAI22_X1 port map( A1 => n98854, A2 => n120560, B1 => n120788, B2 
                           => n120554, ZN => n7092);
   U87672 : OAI22_X1 port map( A1 => n98853, A2 => n120560, B1 => n120791, B2 
                           => n120554, ZN => n7093);
   U87673 : OAI22_X1 port map( A1 => n98852, A2 => n120560, B1 => n120794, B2 
                           => n120554, ZN => n7094);
   U87674 : OAI22_X1 port map( A1 => n98851, A2 => n120560, B1 => n120797, B2 
                           => n120554, ZN => n7095);
   U87675 : OAI22_X1 port map( A1 => n98850, A2 => n120560, B1 => n120800, B2 
                           => n120554, ZN => n7096);
   U87676 : OAI22_X1 port map( A1 => n98849, A2 => n120560, B1 => n120803, B2 
                           => n120554, ZN => n7097);
   U87677 : OAI22_X1 port map( A1 => n98848, A2 => n120561, B1 => n120806, B2 
                           => n120554, ZN => n7098);
   U87678 : OAI22_X1 port map( A1 => n98582, A2 => n120617, B1 => n120629, B2 
                           => n120611, ZN => n7359);
   U87679 : OAI22_X1 port map( A1 => n98581, A2 => n120617, B1 => n120632, B2 
                           => n120611, ZN => n7360);
   U87680 : OAI22_X1 port map( A1 => n98580, A2 => n120617, B1 => n120635, B2 
                           => n120611, ZN => n7361);
   U87681 : OAI22_X1 port map( A1 => n98579, A2 => n120617, B1 => n120638, B2 
                           => n120611, ZN => n7362);
   U87682 : OAI22_X1 port map( A1 => n98578, A2 => n120617, B1 => n120641, B2 
                           => n120611, ZN => n7363);
   U87683 : OAI22_X1 port map( A1 => n98577, A2 => n120617, B1 => n120644, B2 
                           => n120611, ZN => n7364);
   U87684 : OAI22_X1 port map( A1 => n98576, A2 => n120617, B1 => n120647, B2 
                           => n120611, ZN => n7365);
   U87685 : OAI22_X1 port map( A1 => n98575, A2 => n120617, B1 => n120650, B2 
                           => n120611, ZN => n7366);
   U87686 : OAI22_X1 port map( A1 => n98574, A2 => n120617, B1 => n120653, B2 
                           => n120611, ZN => n7367);
   U87687 : OAI22_X1 port map( A1 => n98573, A2 => n120617, B1 => n120656, B2 
                           => n120611, ZN => n7368);
   U87688 : OAI22_X1 port map( A1 => n98572, A2 => n120617, B1 => n120659, B2 
                           => n120611, ZN => n7369);
   U87689 : OAI22_X1 port map( A1 => n98571, A2 => n120618, B1 => n120662, B2 
                           => n120611, ZN => n7370);
   U87690 : OAI22_X1 port map( A1 => n98570, A2 => n120618, B1 => n120665, B2 
                           => n120612, ZN => n7371);
   U87691 : OAI22_X1 port map( A1 => n98569, A2 => n120618, B1 => n120668, B2 
                           => n120612, ZN => n7372);
   U87692 : OAI22_X1 port map( A1 => n98568, A2 => n120618, B1 => n120671, B2 
                           => n120612, ZN => n7373);
   U87693 : OAI22_X1 port map( A1 => n98567, A2 => n120618, B1 => n120674, B2 
                           => n120612, ZN => n7374);
   U87694 : OAI22_X1 port map( A1 => n98566, A2 => n120618, B1 => n120677, B2 
                           => n120612, ZN => n7375);
   U87695 : OAI22_X1 port map( A1 => n98565, A2 => n120618, B1 => n120680, B2 
                           => n120612, ZN => n7376);
   U87696 : OAI22_X1 port map( A1 => n98564, A2 => n120618, B1 => n120683, B2 
                           => n120612, ZN => n7377);
   U87697 : OAI22_X1 port map( A1 => n98563, A2 => n120618, B1 => n120686, B2 
                           => n120612, ZN => n7378);
   U87698 : OAI22_X1 port map( A1 => n98562, A2 => n120618, B1 => n120689, B2 
                           => n120612, ZN => n7379);
   U87699 : OAI22_X1 port map( A1 => n98561, A2 => n120618, B1 => n120692, B2 
                           => n120612, ZN => n7380);
   U87700 : OAI22_X1 port map( A1 => n98560, A2 => n120618, B1 => n120695, B2 
                           => n120612, ZN => n7381);
   U87701 : OAI22_X1 port map( A1 => n98559, A2 => n120619, B1 => n120698, B2 
                           => n120612, ZN => n7382);
   U87702 : OAI22_X1 port map( A1 => n98558, A2 => n120619, B1 => n120701, B2 
                           => n120613, ZN => n7383);
   U87703 : OAI22_X1 port map( A1 => n98557, A2 => n120619, B1 => n120704, B2 
                           => n120613, ZN => n7384);
   U87704 : OAI22_X1 port map( A1 => n98556, A2 => n120619, B1 => n120707, B2 
                           => n120613, ZN => n7385);
   U87705 : OAI22_X1 port map( A1 => n98555, A2 => n120619, B1 => n120710, B2 
                           => n120613, ZN => n7386);
   U87706 : OAI22_X1 port map( A1 => n98554, A2 => n120619, B1 => n120713, B2 
                           => n120613, ZN => n7387);
   U87707 : OAI22_X1 port map( A1 => n98553, A2 => n120619, B1 => n120716, B2 
                           => n120613, ZN => n7388);
   U87708 : OAI22_X1 port map( A1 => n98552, A2 => n120619, B1 => n120719, B2 
                           => n120613, ZN => n7389);
   U87709 : OAI22_X1 port map( A1 => n98551, A2 => n120619, B1 => n120722, B2 
                           => n120613, ZN => n7390);
   U87710 : OAI22_X1 port map( A1 => n98550, A2 => n120619, B1 => n120725, B2 
                           => n120613, ZN => n7391);
   U87711 : OAI22_X1 port map( A1 => n98549, A2 => n120619, B1 => n120728, B2 
                           => n120613, ZN => n7392);
   U87712 : OAI22_X1 port map( A1 => n98548, A2 => n120619, B1 => n120731, B2 
                           => n120613, ZN => n7393);
   U87713 : OAI22_X1 port map( A1 => n98547, A2 => n120620, B1 => n120734, B2 
                           => n120613, ZN => n7394);
   U87714 : OAI22_X1 port map( A1 => n98546, A2 => n120620, B1 => n120737, B2 
                           => n120614, ZN => n7395);
   U87715 : OAI22_X1 port map( A1 => n98545, A2 => n120620, B1 => n120740, B2 
                           => n120614, ZN => n7396);
   U87716 : OAI22_X1 port map( A1 => n98544, A2 => n120620, B1 => n120743, B2 
                           => n120614, ZN => n7397);
   U87717 : OAI22_X1 port map( A1 => n98543, A2 => n120620, B1 => n120746, B2 
                           => n120614, ZN => n7398);
   U87718 : OAI22_X1 port map( A1 => n98542, A2 => n120620, B1 => n120749, B2 
                           => n120614, ZN => n7399);
   U87719 : OAI22_X1 port map( A1 => n98541, A2 => n120620, B1 => n120752, B2 
                           => n120614, ZN => n7400);
   U87720 : OAI22_X1 port map( A1 => n98540, A2 => n120620, B1 => n120755, B2 
                           => n120614, ZN => n7401);
   U87721 : OAI22_X1 port map( A1 => n98539, A2 => n120620, B1 => n120758, B2 
                           => n120614, ZN => n7402);
   U87722 : OAI22_X1 port map( A1 => n98538, A2 => n120620, B1 => n120761, B2 
                           => n120614, ZN => n7403);
   U87723 : OAI22_X1 port map( A1 => n98537, A2 => n120620, B1 => n120764, B2 
                           => n120614, ZN => n7404);
   U87724 : OAI22_X1 port map( A1 => n98536, A2 => n120620, B1 => n120767, B2 
                           => n120614, ZN => n7405);
   U87725 : OAI22_X1 port map( A1 => n98535, A2 => n120621, B1 => n120770, B2 
                           => n120614, ZN => n7406);
   U87726 : OAI22_X1 port map( A1 => n98534, A2 => n120621, B1 => n120773, B2 
                           => n120615, ZN => n7407);
   U87727 : OAI22_X1 port map( A1 => n98533, A2 => n120621, B1 => n120776, B2 
                           => n120615, ZN => n7408);
   U87728 : OAI22_X1 port map( A1 => n98532, A2 => n120621, B1 => n120779, B2 
                           => n120615, ZN => n7409);
   U87729 : OAI22_X1 port map( A1 => n98531, A2 => n120621, B1 => n120782, B2 
                           => n120615, ZN => n7410);
   U87730 : OAI22_X1 port map( A1 => n98530, A2 => n120621, B1 => n120785, B2 
                           => n120615, ZN => n7411);
   U87731 : OAI22_X1 port map( A1 => n98529, A2 => n120621, B1 => n120788, B2 
                           => n120615, ZN => n7412);
   U87732 : OAI22_X1 port map( A1 => n98528, A2 => n120621, B1 => n120791, B2 
                           => n120615, ZN => n7413);
   U87733 : OAI22_X1 port map( A1 => n98527, A2 => n120621, B1 => n120794, B2 
                           => n120615, ZN => n7414);
   U87734 : OAI22_X1 port map( A1 => n98526, A2 => n120621, B1 => n120797, B2 
                           => n120615, ZN => n7415);
   U87735 : OAI22_X1 port map( A1 => n98525, A2 => n120621, B1 => n120800, B2 
                           => n120615, ZN => n7416);
   U87736 : OAI22_X1 port map( A1 => n98524, A2 => n120621, B1 => n120803, B2 
                           => n120615, ZN => n7417);
   U87737 : OAI22_X1 port map( A1 => n98523, A2 => n120622, B1 => n120806, B2 
                           => n120615, ZN => n7418);
   U87738 : OAI22_X1 port map( A1 => n98712, A2 => n120593, B1 => n120629, B2 
                           => n120587, ZN => n7231);
   U87739 : OAI22_X1 port map( A1 => n98711, A2 => n120593, B1 => n120632, B2 
                           => n120587, ZN => n7232);
   U87740 : OAI22_X1 port map( A1 => n98710, A2 => n120593, B1 => n120635, B2 
                           => n120587, ZN => n7233);
   U87741 : OAI22_X1 port map( A1 => n98709, A2 => n120593, B1 => n120638, B2 
                           => n120587, ZN => n7234);
   U87742 : OAI22_X1 port map( A1 => n98708, A2 => n120593, B1 => n120641, B2 
                           => n120587, ZN => n7235);
   U87743 : OAI22_X1 port map( A1 => n98707, A2 => n120593, B1 => n120644, B2 
                           => n120587, ZN => n7236);
   U87744 : OAI22_X1 port map( A1 => n98706, A2 => n120593, B1 => n120647, B2 
                           => n120587, ZN => n7237);
   U87745 : OAI22_X1 port map( A1 => n98705, A2 => n120593, B1 => n120650, B2 
                           => n120587, ZN => n7238);
   U87746 : OAI22_X1 port map( A1 => n98704, A2 => n120593, B1 => n120653, B2 
                           => n120587, ZN => n7239);
   U87747 : OAI22_X1 port map( A1 => n98703, A2 => n120593, B1 => n120656, B2 
                           => n120587, ZN => n7240);
   U87748 : OAI22_X1 port map( A1 => n98702, A2 => n120593, B1 => n120659, B2 
                           => n120587, ZN => n7241);
   U87749 : OAI22_X1 port map( A1 => n98701, A2 => n120594, B1 => n120662, B2 
                           => n120587, ZN => n7242);
   U87750 : OAI22_X1 port map( A1 => n98700, A2 => n120594, B1 => n120665, B2 
                           => n120588, ZN => n7243);
   U87751 : OAI22_X1 port map( A1 => n98699, A2 => n120594, B1 => n120668, B2 
                           => n120588, ZN => n7244);
   U87752 : OAI22_X1 port map( A1 => n98698, A2 => n120594, B1 => n120671, B2 
                           => n120588, ZN => n7245);
   U87753 : OAI22_X1 port map( A1 => n98697, A2 => n120594, B1 => n120674, B2 
                           => n120588, ZN => n7246);
   U87754 : OAI22_X1 port map( A1 => n98696, A2 => n120594, B1 => n120677, B2 
                           => n120588, ZN => n7247);
   U87755 : OAI22_X1 port map( A1 => n98695, A2 => n120594, B1 => n120680, B2 
                           => n120588, ZN => n7248);
   U87756 : OAI22_X1 port map( A1 => n98694, A2 => n120594, B1 => n120683, B2 
                           => n120588, ZN => n7249);
   U87757 : OAI22_X1 port map( A1 => n98693, A2 => n120594, B1 => n120686, B2 
                           => n120588, ZN => n7250);
   U87758 : OAI22_X1 port map( A1 => n98692, A2 => n120594, B1 => n120689, B2 
                           => n120588, ZN => n7251);
   U87759 : OAI22_X1 port map( A1 => n98691, A2 => n120594, B1 => n120692, B2 
                           => n120588, ZN => n7252);
   U87760 : OAI22_X1 port map( A1 => n98690, A2 => n120594, B1 => n120695, B2 
                           => n120588, ZN => n7253);
   U87761 : OAI22_X1 port map( A1 => n98689, A2 => n120595, B1 => n120698, B2 
                           => n120588, ZN => n7254);
   U87762 : OAI22_X1 port map( A1 => n98688, A2 => n120595, B1 => n120701, B2 
                           => n120589, ZN => n7255);
   U87763 : OAI22_X1 port map( A1 => n98687, A2 => n120595, B1 => n120704, B2 
                           => n120589, ZN => n7256);
   U87764 : OAI22_X1 port map( A1 => n98686, A2 => n120595, B1 => n120707, B2 
                           => n120589, ZN => n7257);
   U87765 : OAI22_X1 port map( A1 => n98685, A2 => n120595, B1 => n120710, B2 
                           => n120589, ZN => n7258);
   U87766 : OAI22_X1 port map( A1 => n98684, A2 => n120595, B1 => n120713, B2 
                           => n120589, ZN => n7259);
   U87767 : OAI22_X1 port map( A1 => n98683, A2 => n120595, B1 => n120716, B2 
                           => n120589, ZN => n7260);
   U87768 : OAI22_X1 port map( A1 => n98682, A2 => n120595, B1 => n120719, B2 
                           => n120589, ZN => n7261);
   U87769 : OAI22_X1 port map( A1 => n98681, A2 => n120595, B1 => n120722, B2 
                           => n120589, ZN => n7262);
   U87770 : OAI22_X1 port map( A1 => n98680, A2 => n120595, B1 => n120725, B2 
                           => n120589, ZN => n7263);
   U87771 : OAI22_X1 port map( A1 => n98679, A2 => n120595, B1 => n120728, B2 
                           => n120589, ZN => n7264);
   U87772 : OAI22_X1 port map( A1 => n98678, A2 => n120595, B1 => n120731, B2 
                           => n120589, ZN => n7265);
   U87773 : OAI22_X1 port map( A1 => n98677, A2 => n120596, B1 => n120734, B2 
                           => n120589, ZN => n7266);
   U87774 : OAI22_X1 port map( A1 => n98676, A2 => n120596, B1 => n120737, B2 
                           => n120590, ZN => n7267);
   U87775 : OAI22_X1 port map( A1 => n98675, A2 => n120596, B1 => n120740, B2 
                           => n120590, ZN => n7268);
   U87776 : OAI22_X1 port map( A1 => n98674, A2 => n120596, B1 => n120743, B2 
                           => n120590, ZN => n7269);
   U87777 : OAI22_X1 port map( A1 => n98673, A2 => n120596, B1 => n120746, B2 
                           => n120590, ZN => n7270);
   U87778 : OAI22_X1 port map( A1 => n98672, A2 => n120596, B1 => n120749, B2 
                           => n120590, ZN => n7271);
   U87779 : OAI22_X1 port map( A1 => n98671, A2 => n120596, B1 => n120752, B2 
                           => n120590, ZN => n7272);
   U87780 : OAI22_X1 port map( A1 => n98670, A2 => n120596, B1 => n120755, B2 
                           => n120590, ZN => n7273);
   U87781 : OAI22_X1 port map( A1 => n98669, A2 => n120596, B1 => n120758, B2 
                           => n120590, ZN => n7274);
   U87782 : OAI22_X1 port map( A1 => n98668, A2 => n120596, B1 => n120761, B2 
                           => n120590, ZN => n7275);
   U87783 : OAI22_X1 port map( A1 => n98667, A2 => n120596, B1 => n120764, B2 
                           => n120590, ZN => n7276);
   U87784 : OAI22_X1 port map( A1 => n98666, A2 => n120596, B1 => n120767, B2 
                           => n120590, ZN => n7277);
   U87785 : OAI22_X1 port map( A1 => n98665, A2 => n120597, B1 => n120770, B2 
                           => n120590, ZN => n7278);
   U87786 : OAI22_X1 port map( A1 => n98664, A2 => n120597, B1 => n120773, B2 
                           => n120591, ZN => n7279);
   U87787 : OAI22_X1 port map( A1 => n98663, A2 => n120597, B1 => n120776, B2 
                           => n120591, ZN => n7280);
   U87788 : OAI22_X1 port map( A1 => n98662, A2 => n120597, B1 => n120779, B2 
                           => n120591, ZN => n7281);
   U87789 : OAI22_X1 port map( A1 => n98661, A2 => n120597, B1 => n120782, B2 
                           => n120591, ZN => n7282);
   U87790 : OAI22_X1 port map( A1 => n98660, A2 => n120597, B1 => n120785, B2 
                           => n120591, ZN => n7283);
   U87791 : OAI22_X1 port map( A1 => n98659, A2 => n120597, B1 => n120788, B2 
                           => n120591, ZN => n7284);
   U87792 : OAI22_X1 port map( A1 => n98658, A2 => n120597, B1 => n120791, B2 
                           => n120591, ZN => n7285);
   U87793 : OAI22_X1 port map( A1 => n98657, A2 => n120597, B1 => n120794, B2 
                           => n120591, ZN => n7286);
   U87794 : OAI22_X1 port map( A1 => n98656, A2 => n120597, B1 => n120797, B2 
                           => n120591, ZN => n7287);
   U87795 : OAI22_X1 port map( A1 => n98655, A2 => n120597, B1 => n120800, B2 
                           => n120591, ZN => n7288);
   U87796 : OAI22_X1 port map( A1 => n98654, A2 => n120597, B1 => n120803, B2 
                           => n120591, ZN => n7289);
   U87797 : OAI22_X1 port map( A1 => n98653, A2 => n120598, B1 => n120806, B2 
                           => n120591, ZN => n7290);
   U87798 : OAI22_X1 port map( A1 => n98645, A2 => n120605, B1 => n120629, B2 
                           => n120599, ZN => n7295);
   U87799 : OAI22_X1 port map( A1 => n98644, A2 => n120605, B1 => n120632, B2 
                           => n120599, ZN => n7296);
   U87800 : OAI22_X1 port map( A1 => n98643, A2 => n120605, B1 => n120635, B2 
                           => n120599, ZN => n7297);
   U87801 : OAI22_X1 port map( A1 => n98642, A2 => n120605, B1 => n120638, B2 
                           => n120599, ZN => n7298);
   U87802 : OAI22_X1 port map( A1 => n98641, A2 => n120605, B1 => n120641, B2 
                           => n120599, ZN => n7299);
   U87803 : OAI22_X1 port map( A1 => n98640, A2 => n120605, B1 => n120644, B2 
                           => n120599, ZN => n7300);
   U87804 : OAI22_X1 port map( A1 => n98639, A2 => n120605, B1 => n120647, B2 
                           => n120599, ZN => n7301);
   U87805 : OAI22_X1 port map( A1 => n98638, A2 => n120605, B1 => n120650, B2 
                           => n120599, ZN => n7302);
   U87806 : OAI22_X1 port map( A1 => n98637, A2 => n120605, B1 => n120653, B2 
                           => n120599, ZN => n7303);
   U87807 : OAI22_X1 port map( A1 => n98636, A2 => n120605, B1 => n120656, B2 
                           => n120599, ZN => n7304);
   U87808 : OAI22_X1 port map( A1 => n98635, A2 => n120605, B1 => n120659, B2 
                           => n120599, ZN => n7305);
   U87809 : OAI22_X1 port map( A1 => n98634, A2 => n120606, B1 => n120662, B2 
                           => n120599, ZN => n7306);
   U87810 : OAI22_X1 port map( A1 => n98633, A2 => n120606, B1 => n120665, B2 
                           => n120600, ZN => n7307);
   U87811 : OAI22_X1 port map( A1 => n98632, A2 => n120606, B1 => n120668, B2 
                           => n120600, ZN => n7308);
   U87812 : OAI22_X1 port map( A1 => n98631, A2 => n120606, B1 => n120671, B2 
                           => n120600, ZN => n7309);
   U87813 : OAI22_X1 port map( A1 => n98630, A2 => n120606, B1 => n120674, B2 
                           => n120600, ZN => n7310);
   U87814 : OAI22_X1 port map( A1 => n98629, A2 => n120606, B1 => n120677, B2 
                           => n120600, ZN => n7311);
   U87815 : OAI22_X1 port map( A1 => n98628, A2 => n120606, B1 => n120680, B2 
                           => n120600, ZN => n7312);
   U87816 : OAI22_X1 port map( A1 => n98627, A2 => n120606, B1 => n120683, B2 
                           => n120600, ZN => n7313);
   U87817 : OAI22_X1 port map( A1 => n98626, A2 => n120606, B1 => n120686, B2 
                           => n120600, ZN => n7314);
   U87818 : OAI22_X1 port map( A1 => n98625, A2 => n120606, B1 => n120689, B2 
                           => n120600, ZN => n7315);
   U87819 : OAI22_X1 port map( A1 => n98624, A2 => n120606, B1 => n120692, B2 
                           => n120600, ZN => n7316);
   U87820 : OAI22_X1 port map( A1 => n98623, A2 => n120606, B1 => n120695, B2 
                           => n120600, ZN => n7317);
   U87821 : OAI22_X1 port map( A1 => n98622, A2 => n120607, B1 => n120698, B2 
                           => n120600, ZN => n7318);
   U87822 : OAI22_X1 port map( A1 => n98621, A2 => n120607, B1 => n120701, B2 
                           => n120601, ZN => n7319);
   U87823 : OAI22_X1 port map( A1 => n98620, A2 => n120607, B1 => n120704, B2 
                           => n120601, ZN => n7320);
   U87824 : OAI22_X1 port map( A1 => n98619, A2 => n120607, B1 => n120707, B2 
                           => n120601, ZN => n7321);
   U87825 : OAI22_X1 port map( A1 => n98618, A2 => n120607, B1 => n120710, B2 
                           => n120601, ZN => n7322);
   U87826 : OAI22_X1 port map( A1 => n98617, A2 => n120607, B1 => n120713, B2 
                           => n120601, ZN => n7323);
   U87827 : OAI22_X1 port map( A1 => n98616, A2 => n120607, B1 => n120716, B2 
                           => n120601, ZN => n7324);
   U87828 : OAI22_X1 port map( A1 => n98615, A2 => n120607, B1 => n120719, B2 
                           => n120601, ZN => n7325);
   U87829 : OAI22_X1 port map( A1 => n98614, A2 => n120607, B1 => n120722, B2 
                           => n120601, ZN => n7326);
   U87830 : OAI22_X1 port map( A1 => n98613, A2 => n120607, B1 => n120725, B2 
                           => n120601, ZN => n7327);
   U87831 : OAI22_X1 port map( A1 => n98612, A2 => n120607, B1 => n120728, B2 
                           => n120601, ZN => n7328);
   U87832 : OAI22_X1 port map( A1 => n98611, A2 => n120607, B1 => n120731, B2 
                           => n120601, ZN => n7329);
   U87833 : OAI22_X1 port map( A1 => n98610, A2 => n120608, B1 => n120734, B2 
                           => n120601, ZN => n7330);
   U87834 : OAI22_X1 port map( A1 => n98609, A2 => n120608, B1 => n120737, B2 
                           => n120602, ZN => n7331);
   U87835 : OAI22_X1 port map( A1 => n98608, A2 => n120608, B1 => n120740, B2 
                           => n120602, ZN => n7332);
   U87836 : OAI22_X1 port map( A1 => n98607, A2 => n120608, B1 => n120743, B2 
                           => n120602, ZN => n7333);
   U87837 : OAI22_X1 port map( A1 => n98606, A2 => n120608, B1 => n120746, B2 
                           => n120602, ZN => n7334);
   U87838 : OAI22_X1 port map( A1 => n98605, A2 => n120608, B1 => n120749, B2 
                           => n120602, ZN => n7335);
   U87839 : OAI22_X1 port map( A1 => n98604, A2 => n120608, B1 => n120752, B2 
                           => n120602, ZN => n7336);
   U87840 : OAI22_X1 port map( A1 => n98603, A2 => n120608, B1 => n120755, B2 
                           => n120602, ZN => n7337);
   U87841 : OAI22_X1 port map( A1 => n98602, A2 => n120608, B1 => n120758, B2 
                           => n120602, ZN => n7338);
   U87842 : OAI22_X1 port map( A1 => n98601, A2 => n120608, B1 => n120761, B2 
                           => n120602, ZN => n7339);
   U87843 : OAI22_X1 port map( A1 => n98600, A2 => n120608, B1 => n120764, B2 
                           => n120602, ZN => n7340);
   U87844 : OAI22_X1 port map( A1 => n98599, A2 => n120608, B1 => n120767, B2 
                           => n120602, ZN => n7341);
   U87845 : OAI22_X1 port map( A1 => n98598, A2 => n120609, B1 => n120770, B2 
                           => n120602, ZN => n7342);
   U87846 : OAI22_X1 port map( A1 => n98597, A2 => n120609, B1 => n120773, B2 
                           => n120603, ZN => n7343);
   U87847 : OAI22_X1 port map( A1 => n98596, A2 => n120609, B1 => n120776, B2 
                           => n120603, ZN => n7344);
   U87848 : OAI22_X1 port map( A1 => n98595, A2 => n120609, B1 => n120779, B2 
                           => n120603, ZN => n7345);
   U87849 : OAI22_X1 port map( A1 => n98594, A2 => n120609, B1 => n120782, B2 
                           => n120603, ZN => n7346);
   U87850 : OAI22_X1 port map( A1 => n98593, A2 => n120609, B1 => n120785, B2 
                           => n120603, ZN => n7347);
   U87851 : OAI22_X1 port map( A1 => n98592, A2 => n120609, B1 => n120788, B2 
                           => n120603, ZN => n7348);
   U87852 : OAI22_X1 port map( A1 => n98591, A2 => n120609, B1 => n120791, B2 
                           => n120603, ZN => n7349);
   U87853 : OAI22_X1 port map( A1 => n98590, A2 => n120609, B1 => n120794, B2 
                           => n120603, ZN => n7350);
   U87854 : OAI22_X1 port map( A1 => n98589, A2 => n120609, B1 => n120797, B2 
                           => n120603, ZN => n7351);
   U87855 : OAI22_X1 port map( A1 => n98588, A2 => n120609, B1 => n120800, B2 
                           => n120603, ZN => n7352);
   U87856 : OAI22_X1 port map( A1 => n98587, A2 => n120609, B1 => n120803, B2 
                           => n120603, ZN => n7353);
   U87857 : OAI22_X1 port map( A1 => n98586, A2 => n120610, B1 => n120806, B2 
                           => n120603, ZN => n7354);
   U87858 : OAI22_X1 port map( A1 => n99644, A2 => n120360, B1 => n120630, B2 
                           => n120354, ZN => n6015);
   U87859 : OAI22_X1 port map( A1 => n99643, A2 => n120360, B1 => n120633, B2 
                           => n120354, ZN => n6016);
   U87860 : OAI22_X1 port map( A1 => n99642, A2 => n120360, B1 => n120636, B2 
                           => n120354, ZN => n6017);
   U87861 : OAI22_X1 port map( A1 => n99641, A2 => n120360, B1 => n120639, B2 
                           => n120354, ZN => n6018);
   U87862 : OAI22_X1 port map( A1 => n99640, A2 => n120360, B1 => n120642, B2 
                           => n120354, ZN => n6019);
   U87863 : OAI22_X1 port map( A1 => n99639, A2 => n120360, B1 => n120645, B2 
                           => n120354, ZN => n6020);
   U87864 : OAI22_X1 port map( A1 => n99638, A2 => n120360, B1 => n120648, B2 
                           => n120354, ZN => n6021);
   U87865 : OAI22_X1 port map( A1 => n99637, A2 => n120360, B1 => n120651, B2 
                           => n120354, ZN => n6022);
   U87866 : OAI22_X1 port map( A1 => n99636, A2 => n120360, B1 => n120654, B2 
                           => n120354, ZN => n6023);
   U87867 : OAI22_X1 port map( A1 => n99635, A2 => n120360, B1 => n120657, B2 
                           => n120354, ZN => n6024);
   U87868 : OAI22_X1 port map( A1 => n99634, A2 => n120360, B1 => n120660, B2 
                           => n120354, ZN => n6025);
   U87869 : OAI22_X1 port map( A1 => n99633, A2 => n120361, B1 => n120663, B2 
                           => n120354, ZN => n6026);
   U87870 : OAI22_X1 port map( A1 => n99632, A2 => n120361, B1 => n120666, B2 
                           => n120355, ZN => n6027);
   U87871 : OAI22_X1 port map( A1 => n99631, A2 => n120361, B1 => n120669, B2 
                           => n120355, ZN => n6028);
   U87872 : OAI22_X1 port map( A1 => n99630, A2 => n120361, B1 => n120672, B2 
                           => n120355, ZN => n6029);
   U87873 : OAI22_X1 port map( A1 => n99629, A2 => n120361, B1 => n120675, B2 
                           => n120355, ZN => n6030);
   U87874 : OAI22_X1 port map( A1 => n99628, A2 => n120361, B1 => n120678, B2 
                           => n120355, ZN => n6031);
   U87875 : OAI22_X1 port map( A1 => n99627, A2 => n120361, B1 => n120681, B2 
                           => n120355, ZN => n6032);
   U87876 : OAI22_X1 port map( A1 => n99626, A2 => n120361, B1 => n120684, B2 
                           => n120355, ZN => n6033);
   U87877 : OAI22_X1 port map( A1 => n99625, A2 => n120361, B1 => n120687, B2 
                           => n120355, ZN => n6034);
   U87878 : OAI22_X1 port map( A1 => n99624, A2 => n120361, B1 => n120690, B2 
                           => n120355, ZN => n6035);
   U87879 : OAI22_X1 port map( A1 => n99623, A2 => n120361, B1 => n120693, B2 
                           => n120355, ZN => n6036);
   U87880 : OAI22_X1 port map( A1 => n99622, A2 => n120361, B1 => n120696, B2 
                           => n120355, ZN => n6037);
   U87881 : OAI22_X1 port map( A1 => n99621, A2 => n120362, B1 => n120699, B2 
                           => n120355, ZN => n6038);
   U87882 : OAI22_X1 port map( A1 => n99620, A2 => n120362, B1 => n120702, B2 
                           => n120356, ZN => n6039);
   U87883 : OAI22_X1 port map( A1 => n99619, A2 => n120362, B1 => n120705, B2 
                           => n120356, ZN => n6040);
   U87884 : OAI22_X1 port map( A1 => n99618, A2 => n120362, B1 => n120708, B2 
                           => n120356, ZN => n6041);
   U87885 : OAI22_X1 port map( A1 => n99617, A2 => n120362, B1 => n120711, B2 
                           => n120356, ZN => n6042);
   U87886 : OAI22_X1 port map( A1 => n99616, A2 => n120362, B1 => n120714, B2 
                           => n120356, ZN => n6043);
   U87887 : OAI22_X1 port map( A1 => n99615, A2 => n120362, B1 => n120717, B2 
                           => n120356, ZN => n6044);
   U87888 : OAI22_X1 port map( A1 => n99614, A2 => n120362, B1 => n120720, B2 
                           => n120356, ZN => n6045);
   U87889 : OAI22_X1 port map( A1 => n99613, A2 => n120362, B1 => n120723, B2 
                           => n120356, ZN => n6046);
   U87890 : OAI22_X1 port map( A1 => n99612, A2 => n120362, B1 => n120726, B2 
                           => n120356, ZN => n6047);
   U87891 : OAI22_X1 port map( A1 => n99611, A2 => n120362, B1 => n120729, B2 
                           => n120356, ZN => n6048);
   U87892 : OAI22_X1 port map( A1 => n99610, A2 => n120362, B1 => n120732, B2 
                           => n120356, ZN => n6049);
   U87893 : OAI22_X1 port map( A1 => n99609, A2 => n120363, B1 => n120735, B2 
                           => n120356, ZN => n6050);
   U87894 : OAI22_X1 port map( A1 => n99608, A2 => n120363, B1 => n120738, B2 
                           => n120357, ZN => n6051);
   U87895 : OAI22_X1 port map( A1 => n99607, A2 => n120363, B1 => n120741, B2 
                           => n120357, ZN => n6052);
   U87896 : OAI22_X1 port map( A1 => n99606, A2 => n120363, B1 => n120744, B2 
                           => n120357, ZN => n6053);
   U87897 : OAI22_X1 port map( A1 => n99605, A2 => n120363, B1 => n120747, B2 
                           => n120357, ZN => n6054);
   U87898 : OAI22_X1 port map( A1 => n99604, A2 => n120363, B1 => n120750, B2 
                           => n120357, ZN => n6055);
   U87899 : OAI22_X1 port map( A1 => n99603, A2 => n120363, B1 => n120753, B2 
                           => n120357, ZN => n6056);
   U87900 : OAI22_X1 port map( A1 => n99602, A2 => n120363, B1 => n120756, B2 
                           => n120357, ZN => n6057);
   U87901 : OAI22_X1 port map( A1 => n99601, A2 => n120363, B1 => n120759, B2 
                           => n120357, ZN => n6058);
   U87902 : OAI22_X1 port map( A1 => n99600, A2 => n120363, B1 => n120762, B2 
                           => n120357, ZN => n6059);
   U87903 : OAI22_X1 port map( A1 => n99599, A2 => n120363, B1 => n120765, B2 
                           => n120357, ZN => n6060);
   U87904 : OAI22_X1 port map( A1 => n99598, A2 => n120363, B1 => n120768, B2 
                           => n120357, ZN => n6061);
   U87905 : OAI22_X1 port map( A1 => n99597, A2 => n120364, B1 => n120771, B2 
                           => n120357, ZN => n6062);
   U87906 : OAI22_X1 port map( A1 => n99596, A2 => n120364, B1 => n120774, B2 
                           => n120358, ZN => n6063);
   U87907 : OAI22_X1 port map( A1 => n99595, A2 => n120364, B1 => n120777, B2 
                           => n120358, ZN => n6064);
   U87908 : OAI22_X1 port map( A1 => n99594, A2 => n120364, B1 => n120780, B2 
                           => n120358, ZN => n6065);
   U87909 : OAI22_X1 port map( A1 => n99593, A2 => n120364, B1 => n120783, B2 
                           => n120358, ZN => n6066);
   U87910 : OAI22_X1 port map( A1 => n99592, A2 => n120364, B1 => n120786, B2 
                           => n120358, ZN => n6067);
   U87911 : OAI22_X1 port map( A1 => n99591, A2 => n120364, B1 => n120789, B2 
                           => n120358, ZN => n6068);
   U87912 : OAI22_X1 port map( A1 => n99590, A2 => n120364, B1 => n120792, B2 
                           => n120358, ZN => n6069);
   U87913 : OAI22_X1 port map( A1 => n99589, A2 => n120364, B1 => n120795, B2 
                           => n120358, ZN => n6070);
   U87914 : OAI22_X1 port map( A1 => n99588, A2 => n120364, B1 => n120798, B2 
                           => n120358, ZN => n6071);
   U87915 : OAI22_X1 port map( A1 => n99587, A2 => n120364, B1 => n120801, B2 
                           => n120358, ZN => n6072);
   U87916 : OAI22_X1 port map( A1 => n99586, A2 => n120364, B1 => n120804, B2 
                           => n120358, ZN => n6073);
   U87917 : OAI22_X1 port map( A1 => n99585, A2 => n120365, B1 => n120807, B2 
                           => n120358, ZN => n6074);
   U87918 : OAI22_X1 port map( A1 => n120337, A2 => n114370, B1 => n120630, B2 
                           => n120329, ZN => n5887);
   U87919 : OAI22_X1 port map( A1 => n120337, A2 => n114369, B1 => n120633, B2 
                           => n120329, ZN => n5888);
   U87920 : OAI22_X1 port map( A1 => n120337, A2 => n114368, B1 => n120636, B2 
                           => n120329, ZN => n5889);
   U87921 : OAI22_X1 port map( A1 => n120337, A2 => n114367, B1 => n120639, B2 
                           => n120329, ZN => n5890);
   U87922 : OAI22_X1 port map( A1 => n120337, A2 => n114366, B1 => n120642, B2 
                           => n120329, ZN => n5891);
   U87923 : OAI22_X1 port map( A1 => n120337, A2 => n114365, B1 => n120645, B2 
                           => n120329, ZN => n5892);
   U87924 : OAI22_X1 port map( A1 => n120337, A2 => n114364, B1 => n120648, B2 
                           => n120329, ZN => n5893);
   U87925 : OAI22_X1 port map( A1 => n120337, A2 => n114363, B1 => n120651, B2 
                           => n120329, ZN => n5894);
   U87926 : OAI22_X1 port map( A1 => n120337, A2 => n114362, B1 => n120654, B2 
                           => n120329, ZN => n5895);
   U87927 : OAI22_X1 port map( A1 => n120337, A2 => n114361, B1 => n120657, B2 
                           => n120329, ZN => n5896);
   U87928 : OAI22_X1 port map( A1 => n120337, A2 => n114360, B1 => n120660, B2 
                           => n120329, ZN => n5897);
   U87929 : OAI22_X1 port map( A1 => n120337, A2 => n114359, B1 => n120663, B2 
                           => n120329, ZN => n5898);
   U87930 : OAI22_X1 port map( A1 => n120338, A2 => n114358, B1 => n120666, B2 
                           => n120330, ZN => n5899);
   U87931 : OAI22_X1 port map( A1 => n120338, A2 => n114357, B1 => n120669, B2 
                           => n120330, ZN => n5900);
   U87932 : OAI22_X1 port map( A1 => n120338, A2 => n114356, B1 => n120672, B2 
                           => n120330, ZN => n5901);
   U87933 : OAI22_X1 port map( A1 => n120338, A2 => n114355, B1 => n120675, B2 
                           => n120330, ZN => n5902);
   U87934 : OAI22_X1 port map( A1 => n120338, A2 => n114354, B1 => n120678, B2 
                           => n120330, ZN => n5903);
   U87935 : OAI22_X1 port map( A1 => n120338, A2 => n114353, B1 => n120681, B2 
                           => n120330, ZN => n5904);
   U87936 : OAI22_X1 port map( A1 => n120338, A2 => n114352, B1 => n120684, B2 
                           => n120330, ZN => n5905);
   U87937 : OAI22_X1 port map( A1 => n120338, A2 => n114351, B1 => n120687, B2 
                           => n120330, ZN => n5906);
   U87938 : OAI22_X1 port map( A1 => n120338, A2 => n114350, B1 => n120690, B2 
                           => n120330, ZN => n5907);
   U87939 : OAI22_X1 port map( A1 => n120338, A2 => n114349, B1 => n120693, B2 
                           => n120330, ZN => n5908);
   U87940 : OAI22_X1 port map( A1 => n120338, A2 => n114348, B1 => n120696, B2 
                           => n120330, ZN => n5909);
   U87941 : OAI22_X1 port map( A1 => n120338, A2 => n114347, B1 => n120699, B2 
                           => n120330, ZN => n5910);
   U87942 : OAI22_X1 port map( A1 => n120338, A2 => n114346, B1 => n120702, B2 
                           => n120331, ZN => n5911);
   U87943 : OAI22_X1 port map( A1 => n120339, A2 => n114345, B1 => n120705, B2 
                           => n120331, ZN => n5912);
   U87944 : OAI22_X1 port map( A1 => n120339, A2 => n114344, B1 => n120708, B2 
                           => n120331, ZN => n5913);
   U87945 : OAI22_X1 port map( A1 => n120339, A2 => n114343, B1 => n120711, B2 
                           => n120331, ZN => n5914);
   U87946 : OAI22_X1 port map( A1 => n120339, A2 => n114342, B1 => n120714, B2 
                           => n120331, ZN => n5915);
   U87947 : OAI22_X1 port map( A1 => n120339, A2 => n114341, B1 => n120717, B2 
                           => n120331, ZN => n5916);
   U87948 : OAI22_X1 port map( A1 => n120339, A2 => n114340, B1 => n120720, B2 
                           => n120331, ZN => n5917);
   U87949 : OAI22_X1 port map( A1 => n120339, A2 => n114339, B1 => n120723, B2 
                           => n120331, ZN => n5918);
   U87950 : OAI22_X1 port map( A1 => n120339, A2 => n114338, B1 => n120726, B2 
                           => n120331, ZN => n5919);
   U87951 : OAI22_X1 port map( A1 => n120339, A2 => n114337, B1 => n120729, B2 
                           => n120331, ZN => n5920);
   U87952 : OAI22_X1 port map( A1 => n120339, A2 => n114336, B1 => n120732, B2 
                           => n120331, ZN => n5921);
   U87953 : OAI22_X1 port map( A1 => n120339, A2 => n114335, B1 => n120735, B2 
                           => n120331, ZN => n5922);
   U87954 : OAI22_X1 port map( A1 => n120339, A2 => n114334, B1 => n120738, B2 
                           => n120332, ZN => n5923);
   U87955 : OAI22_X1 port map( A1 => n120339, A2 => n114333, B1 => n120741, B2 
                           => n120332, ZN => n5924);
   U87956 : OAI22_X1 port map( A1 => n120340, A2 => n114332, B1 => n120744, B2 
                           => n120332, ZN => n5925);
   U87957 : OAI22_X1 port map( A1 => n120340, A2 => n114331, B1 => n120747, B2 
                           => n120332, ZN => n5926);
   U87958 : OAI22_X1 port map( A1 => n120340, A2 => n114330, B1 => n120750, B2 
                           => n120332, ZN => n5927);
   U87959 : OAI22_X1 port map( A1 => n120340, A2 => n114329, B1 => n120753, B2 
                           => n120332, ZN => n5928);
   U87960 : OAI22_X1 port map( A1 => n120340, A2 => n114328, B1 => n120756, B2 
                           => n120332, ZN => n5929);
   U87961 : OAI22_X1 port map( A1 => n120340, A2 => n114327, B1 => n120759, B2 
                           => n120332, ZN => n5930);
   U87962 : OAI22_X1 port map( A1 => n120340, A2 => n114326, B1 => n120762, B2 
                           => n120332, ZN => n5931);
   U87963 : OAI22_X1 port map( A1 => n120340, A2 => n114325, B1 => n120765, B2 
                           => n120332, ZN => n5932);
   U87964 : OAI22_X1 port map( A1 => n120340, A2 => n114324, B1 => n120768, B2 
                           => n120332, ZN => n5933);
   U87965 : OAI22_X1 port map( A1 => n120340, A2 => n114323, B1 => n120771, B2 
                           => n120332, ZN => n5934);
   U87966 : OAI22_X1 port map( A1 => n120340, A2 => n114322, B1 => n120774, B2 
                           => n120333, ZN => n5935);
   U87967 : OAI22_X1 port map( A1 => n120340, A2 => n114321, B1 => n120777, B2 
                           => n120333, ZN => n5936);
   U87968 : OAI22_X1 port map( A1 => n120340, A2 => n114320, B1 => n120780, B2 
                           => n120333, ZN => n5937);
   U87969 : OAI22_X1 port map( A1 => n120341, A2 => n114319, B1 => n120783, B2 
                           => n120333, ZN => n5938);
   U87970 : OAI22_X1 port map( A1 => n120341, A2 => n114318, B1 => n120786, B2 
                           => n120333, ZN => n5939);
   U87971 : OAI22_X1 port map( A1 => n120341, A2 => n114317, B1 => n120789, B2 
                           => n120333, ZN => n5940);
   U87972 : OAI22_X1 port map( A1 => n120341, A2 => n114316, B1 => n120792, B2 
                           => n120333, ZN => n5941);
   U87973 : OAI22_X1 port map( A1 => n120341, A2 => n114315, B1 => n120795, B2 
                           => n120333, ZN => n5942);
   U87974 : OAI22_X1 port map( A1 => n120341, A2 => n114314, B1 => n120798, B2 
                           => n120333, ZN => n5943);
   U87975 : OAI22_X1 port map( A1 => n120341, A2 => n114313, B1 => n120801, B2 
                           => n120333, ZN => n5944);
   U87976 : OAI22_X1 port map( A1 => n120341, A2 => n114312, B1 => n120804, B2 
                           => n120333, ZN => n5945);
   U87977 : OAI22_X1 port map( A1 => n120341, A2 => n114311, B1 => n120807, B2 
                           => n120333, ZN => n5946);
   U87978 : OAI22_X1 port map( A1 => n99510, A2 => n120397, B1 => n120630, B2 
                           => n120391, ZN => n6207);
   U87979 : OAI22_X1 port map( A1 => n99509, A2 => n120397, B1 => n120633, B2 
                           => n120391, ZN => n6208);
   U87980 : OAI22_X1 port map( A1 => n99508, A2 => n120397, B1 => n120636, B2 
                           => n120391, ZN => n6209);
   U87981 : OAI22_X1 port map( A1 => n99507, A2 => n120397, B1 => n120639, B2 
                           => n120391, ZN => n6210);
   U87982 : OAI22_X1 port map( A1 => n99506, A2 => n120397, B1 => n120642, B2 
                           => n120391, ZN => n6211);
   U87983 : OAI22_X1 port map( A1 => n99505, A2 => n120397, B1 => n120645, B2 
                           => n120391, ZN => n6212);
   U87984 : OAI22_X1 port map( A1 => n99504, A2 => n120397, B1 => n120648, B2 
                           => n120391, ZN => n6213);
   U87985 : OAI22_X1 port map( A1 => n99503, A2 => n120397, B1 => n120651, B2 
                           => n120391, ZN => n6214);
   U87986 : OAI22_X1 port map( A1 => n99502, A2 => n120397, B1 => n120654, B2 
                           => n120391, ZN => n6215);
   U87987 : OAI22_X1 port map( A1 => n99501, A2 => n120397, B1 => n120657, B2 
                           => n120391, ZN => n6216);
   U87988 : OAI22_X1 port map( A1 => n99500, A2 => n120397, B1 => n120660, B2 
                           => n120391, ZN => n6217);
   U87989 : OAI22_X1 port map( A1 => n99499, A2 => n120398, B1 => n120663, B2 
                           => n120391, ZN => n6218);
   U87990 : OAI22_X1 port map( A1 => n99498, A2 => n120398, B1 => n120666, B2 
                           => n120392, ZN => n6219);
   U87991 : OAI22_X1 port map( A1 => n99497, A2 => n120398, B1 => n120669, B2 
                           => n120392, ZN => n6220);
   U87992 : OAI22_X1 port map( A1 => n99496, A2 => n120398, B1 => n120672, B2 
                           => n120392, ZN => n6221);
   U87993 : OAI22_X1 port map( A1 => n99495, A2 => n120398, B1 => n120675, B2 
                           => n120392, ZN => n6222);
   U87994 : OAI22_X1 port map( A1 => n99494, A2 => n120398, B1 => n120678, B2 
                           => n120392, ZN => n6223);
   U87995 : OAI22_X1 port map( A1 => n99493, A2 => n120398, B1 => n120681, B2 
                           => n120392, ZN => n6224);
   U87996 : OAI22_X1 port map( A1 => n99492, A2 => n120398, B1 => n120684, B2 
                           => n120392, ZN => n6225);
   U87997 : OAI22_X1 port map( A1 => n99491, A2 => n120398, B1 => n120687, B2 
                           => n120392, ZN => n6226);
   U87998 : OAI22_X1 port map( A1 => n99490, A2 => n120398, B1 => n120690, B2 
                           => n120392, ZN => n6227);
   U87999 : OAI22_X1 port map( A1 => n99489, A2 => n120398, B1 => n120693, B2 
                           => n120392, ZN => n6228);
   U88000 : OAI22_X1 port map( A1 => n99488, A2 => n120398, B1 => n120696, B2 
                           => n120392, ZN => n6229);
   U88001 : OAI22_X1 port map( A1 => n99487, A2 => n120399, B1 => n120699, B2 
                           => n120392, ZN => n6230);
   U88002 : OAI22_X1 port map( A1 => n99486, A2 => n120399, B1 => n120702, B2 
                           => n120393, ZN => n6231);
   U88003 : OAI22_X1 port map( A1 => n99485, A2 => n120399, B1 => n120705, B2 
                           => n120393, ZN => n6232);
   U88004 : OAI22_X1 port map( A1 => n99484, A2 => n120399, B1 => n120708, B2 
                           => n120393, ZN => n6233);
   U88005 : OAI22_X1 port map( A1 => n99483, A2 => n120399, B1 => n120711, B2 
                           => n120393, ZN => n6234);
   U88006 : OAI22_X1 port map( A1 => n99482, A2 => n120399, B1 => n120714, B2 
                           => n120393, ZN => n6235);
   U88007 : OAI22_X1 port map( A1 => n99481, A2 => n120399, B1 => n120717, B2 
                           => n120393, ZN => n6236);
   U88008 : OAI22_X1 port map( A1 => n99480, A2 => n120399, B1 => n120720, B2 
                           => n120393, ZN => n6237);
   U88009 : OAI22_X1 port map( A1 => n99479, A2 => n120399, B1 => n120723, B2 
                           => n120393, ZN => n6238);
   U88010 : OAI22_X1 port map( A1 => n99478, A2 => n120399, B1 => n120726, B2 
                           => n120393, ZN => n6239);
   U88011 : OAI22_X1 port map( A1 => n99477, A2 => n120399, B1 => n120729, B2 
                           => n120393, ZN => n6240);
   U88012 : OAI22_X1 port map( A1 => n99476, A2 => n120399, B1 => n120732, B2 
                           => n120393, ZN => n6241);
   U88013 : OAI22_X1 port map( A1 => n99475, A2 => n120400, B1 => n120735, B2 
                           => n120393, ZN => n6242);
   U88014 : OAI22_X1 port map( A1 => n99474, A2 => n120400, B1 => n120738, B2 
                           => n120394, ZN => n6243);
   U88015 : OAI22_X1 port map( A1 => n99473, A2 => n120400, B1 => n120741, B2 
                           => n120394, ZN => n6244);
   U88016 : OAI22_X1 port map( A1 => n99472, A2 => n120400, B1 => n120744, B2 
                           => n120394, ZN => n6245);
   U88017 : OAI22_X1 port map( A1 => n99471, A2 => n120400, B1 => n120747, B2 
                           => n120394, ZN => n6246);
   U88018 : OAI22_X1 port map( A1 => n99470, A2 => n120400, B1 => n120750, B2 
                           => n120394, ZN => n6247);
   U88019 : OAI22_X1 port map( A1 => n99469, A2 => n120400, B1 => n120753, B2 
                           => n120394, ZN => n6248);
   U88020 : OAI22_X1 port map( A1 => n99468, A2 => n120400, B1 => n120756, B2 
                           => n120394, ZN => n6249);
   U88021 : OAI22_X1 port map( A1 => n99467, A2 => n120400, B1 => n120759, B2 
                           => n120394, ZN => n6250);
   U88022 : OAI22_X1 port map( A1 => n99466, A2 => n120400, B1 => n120762, B2 
                           => n120394, ZN => n6251);
   U88023 : OAI22_X1 port map( A1 => n99465, A2 => n120400, B1 => n120765, B2 
                           => n120394, ZN => n6252);
   U88024 : OAI22_X1 port map( A1 => n99464, A2 => n120400, B1 => n120768, B2 
                           => n120394, ZN => n6253);
   U88025 : OAI22_X1 port map( A1 => n99463, A2 => n120401, B1 => n120771, B2 
                           => n120394, ZN => n6254);
   U88026 : OAI22_X1 port map( A1 => n99462, A2 => n120401, B1 => n120774, B2 
                           => n120395, ZN => n6255);
   U88027 : OAI22_X1 port map( A1 => n99461, A2 => n120401, B1 => n120777, B2 
                           => n120395, ZN => n6256);
   U88028 : OAI22_X1 port map( A1 => n99460, A2 => n120401, B1 => n120780, B2 
                           => n120395, ZN => n6257);
   U88029 : OAI22_X1 port map( A1 => n99459, A2 => n120401, B1 => n120783, B2 
                           => n120395, ZN => n6258);
   U88030 : OAI22_X1 port map( A1 => n99458, A2 => n120401, B1 => n120786, B2 
                           => n120395, ZN => n6259);
   U88031 : OAI22_X1 port map( A1 => n99457, A2 => n120401, B1 => n120789, B2 
                           => n120395, ZN => n6260);
   U88032 : OAI22_X1 port map( A1 => n99456, A2 => n120401, B1 => n120792, B2 
                           => n120395, ZN => n6261);
   U88033 : OAI22_X1 port map( A1 => n99455, A2 => n120401, B1 => n120795, B2 
                           => n120395, ZN => n6262);
   U88034 : OAI22_X1 port map( A1 => n99454, A2 => n120401, B1 => n120798, B2 
                           => n120395, ZN => n6263);
   U88035 : OAI22_X1 port map( A1 => n99453, A2 => n120401, B1 => n120801, B2 
                           => n120395, ZN => n6264);
   U88036 : OAI22_X1 port map( A1 => n99452, A2 => n120401, B1 => n120804, B2 
                           => n120395, ZN => n6265);
   U88037 : OAI22_X1 port map( A1 => n99451, A2 => n120402, B1 => n120807, B2 
                           => n120395, ZN => n6266);
   U88038 : OAI22_X1 port map( A1 => n90557, A2 => n120388, B1 => n120687, B2 
                           => n120380, ZN => n6162);
   U88039 : OAI22_X1 port map( A1 => n90556, A2 => n120388, B1 => n120690, B2 
                           => n120380, ZN => n6163);
   U88040 : OAI22_X1 port map( A1 => n90555, A2 => n120388, B1 => n120693, B2 
                           => n120380, ZN => n6164);
   U88041 : OAI22_X1 port map( A1 => n90554, A2 => n120388, B1 => n120696, B2 
                           => n120380, ZN => n6165);
   U88042 : OAI22_X1 port map( A1 => n90553, A2 => n120388, B1 => n120699, B2 
                           => n120380, ZN => n6166);
   U88043 : OAI22_X1 port map( A1 => n90552, A2 => n120388, B1 => n120702, B2 
                           => n120381, ZN => n6167);
   U88044 : OAI22_X1 port map( A1 => n90551, A2 => n120388, B1 => n120705, B2 
                           => n120381, ZN => n6168);
   U88045 : OAI22_X1 port map( A1 => n90550, A2 => n120388, B1 => n120708, B2 
                           => n120381, ZN => n6169);
   U88046 : OAI22_X1 port map( A1 => n90549, A2 => n120388, B1 => n120711, B2 
                           => n120381, ZN => n6170);
   U88047 : OAI22_X1 port map( A1 => n90548, A2 => n120388, B1 => n120714, B2 
                           => n120381, ZN => n6171);
   U88048 : OAI22_X1 port map( A1 => n90547, A2 => n120387, B1 => n120717, B2 
                           => n120381, ZN => n6172);
   U88049 : OAI22_X1 port map( A1 => n90546, A2 => n120387, B1 => n120720, B2 
                           => n120381, ZN => n6173);
   U88050 : OAI22_X1 port map( A1 => n90545, A2 => n120387, B1 => n120723, B2 
                           => n120381, ZN => n6174);
   U88051 : OAI22_X1 port map( A1 => n90544, A2 => n120387, B1 => n120726, B2 
                           => n120381, ZN => n6175);
   U88052 : OAI22_X1 port map( A1 => n90543, A2 => n120387, B1 => n120729, B2 
                           => n120381, ZN => n6176);
   U88053 : OAI22_X1 port map( A1 => n90542, A2 => n120387, B1 => n120732, B2 
                           => n120381, ZN => n6177);
   U88054 : OAI22_X1 port map( A1 => n90541, A2 => n120387, B1 => n120735, B2 
                           => n120381, ZN => n6178);
   U88055 : OAI22_X1 port map( A1 => n90540, A2 => n120387, B1 => n120738, B2 
                           => n120382, ZN => n6179);
   U88056 : OAI22_X1 port map( A1 => n90539, A2 => n120387, B1 => n120741, B2 
                           => n120382, ZN => n6180);
   U88057 : OAI22_X1 port map( A1 => n90538, A2 => n120387, B1 => n120744, B2 
                           => n120382, ZN => n6181);
   U88058 : OAI22_X1 port map( A1 => n90537, A2 => n120387, B1 => n120747, B2 
                           => n120382, ZN => n6182);
   U88059 : OAI22_X1 port map( A1 => n90536, A2 => n120386, B1 => n120750, B2 
                           => n120382, ZN => n6183);
   U88060 : OAI22_X1 port map( A1 => n90535, A2 => n120386, B1 => n120753, B2 
                           => n120382, ZN => n6184);
   U88061 : OAI22_X1 port map( A1 => n90534, A2 => n120386, B1 => n120756, B2 
                           => n120382, ZN => n6185);
   U88062 : OAI22_X1 port map( A1 => n90533, A2 => n120386, B1 => n120759, B2 
                           => n120382, ZN => n6186);
   U88063 : OAI22_X1 port map( A1 => n90532, A2 => n120386, B1 => n120762, B2 
                           => n120382, ZN => n6187);
   U88064 : OAI22_X1 port map( A1 => n90531, A2 => n120386, B1 => n120765, B2 
                           => n120382, ZN => n6188);
   U88065 : OAI22_X1 port map( A1 => n90530, A2 => n120386, B1 => n120768, B2 
                           => n120382, ZN => n6189);
   U88066 : OAI22_X1 port map( A1 => n90529, A2 => n120386, B1 => n120771, B2 
                           => n120382, ZN => n6190);
   U88067 : OAI22_X1 port map( A1 => n90528, A2 => n120386, B1 => n120774, B2 
                           => n120383, ZN => n6191);
   U88068 : OAI22_X1 port map( A1 => n90527, A2 => n120386, B1 => n120777, B2 
                           => n120383, ZN => n6192);
   U88069 : OAI22_X1 port map( A1 => n90526, A2 => n120386, B1 => n120780, B2 
                           => n120383, ZN => n6193);
   U88070 : OAI22_X1 port map( A1 => n90525, A2 => n120386, B1 => n120783, B2 
                           => n120383, ZN => n6194);
   U88071 : OAI22_X1 port map( A1 => n90524, A2 => n120385, B1 => n120786, B2 
                           => n120383, ZN => n6195);
   U88072 : OAI22_X1 port map( A1 => n90523, A2 => n120385, B1 => n120789, B2 
                           => n120383, ZN => n6196);
   U88073 : OAI22_X1 port map( A1 => n90522, A2 => n120385, B1 => n120792, B2 
                           => n120383, ZN => n6197);
   U88074 : OAI22_X1 port map( A1 => n90521, A2 => n120385, B1 => n120795, B2 
                           => n120383, ZN => n6198);
   U88075 : OAI22_X1 port map( A1 => n90520, A2 => n120385, B1 => n120798, B2 
                           => n120383, ZN => n6199);
   U88076 : OAI22_X1 port map( A1 => n90519, A2 => n120385, B1 => n120801, B2 
                           => n120383, ZN => n6200);
   U88077 : OAI22_X1 port map( A1 => n90518, A2 => n120385, B1 => n120804, B2 
                           => n120383, ZN => n6201);
   U88078 : OAI22_X1 port map( A1 => n90517, A2 => n120385, B1 => n120807, B2 
                           => n120383, ZN => n6202);
   U88079 : OAI22_X1 port map( A1 => n90370, A2 => n120434, B1 => n120630, B2 
                           => n120428, ZN => n6399);
   U88080 : OAI22_X1 port map( A1 => n90369, A2 => n120434, B1 => n120633, B2 
                           => n120428, ZN => n6400);
   U88081 : OAI22_X1 port map( A1 => n90368, A2 => n120434, B1 => n120636, B2 
                           => n120428, ZN => n6401);
   U88082 : OAI22_X1 port map( A1 => n90367, A2 => n120434, B1 => n120639, B2 
                           => n120428, ZN => n6402);
   U88083 : OAI22_X1 port map( A1 => n90366, A2 => n120434, B1 => n120642, B2 
                           => n120428, ZN => n6403);
   U88084 : OAI22_X1 port map( A1 => n90365, A2 => n120434, B1 => n120645, B2 
                           => n120428, ZN => n6404);
   U88085 : OAI22_X1 port map( A1 => n90364, A2 => n120434, B1 => n120648, B2 
                           => n120428, ZN => n6405);
   U88086 : OAI22_X1 port map( A1 => n90363, A2 => n120434, B1 => n120651, B2 
                           => n120428, ZN => n6406);
   U88087 : OAI22_X1 port map( A1 => n90362, A2 => n120434, B1 => n120654, B2 
                           => n120428, ZN => n6407);
   U88088 : OAI22_X1 port map( A1 => n90361, A2 => n120434, B1 => n120657, B2 
                           => n120428, ZN => n6408);
   U88089 : OAI22_X1 port map( A1 => n90360, A2 => n120434, B1 => n120660, B2 
                           => n120428, ZN => n6409);
   U88090 : OAI22_X1 port map( A1 => n90359, A2 => n120435, B1 => n120663, B2 
                           => n120428, ZN => n6410);
   U88091 : OAI22_X1 port map( A1 => n90358, A2 => n120435, B1 => n120666, B2 
                           => n120429, ZN => n6411);
   U88092 : OAI22_X1 port map( A1 => n90357, A2 => n120435, B1 => n120669, B2 
                           => n120429, ZN => n6412);
   U88093 : OAI22_X1 port map( A1 => n90356, A2 => n120435, B1 => n120672, B2 
                           => n120429, ZN => n6413);
   U88094 : OAI22_X1 port map( A1 => n90355, A2 => n120435, B1 => n120675, B2 
                           => n120429, ZN => n6414);
   U88095 : OAI22_X1 port map( A1 => n90354, A2 => n120435, B1 => n120678, B2 
                           => n120429, ZN => n6415);
   U88096 : OAI22_X1 port map( A1 => n90353, A2 => n120435, B1 => n120681, B2 
                           => n120429, ZN => n6416);
   U88097 : OAI22_X1 port map( A1 => n90352, A2 => n120435, B1 => n120684, B2 
                           => n120429, ZN => n6417);
   U88098 : OAI22_X1 port map( A1 => n90351, A2 => n120435, B1 => n120687, B2 
                           => n120429, ZN => n6418);
   U88099 : OAI22_X1 port map( A1 => n90350, A2 => n120435, B1 => n120690, B2 
                           => n120429, ZN => n6419);
   U88100 : OAI22_X1 port map( A1 => n90349, A2 => n120435, B1 => n120693, B2 
                           => n120429, ZN => n6420);
   U88101 : OAI22_X1 port map( A1 => n90348, A2 => n120435, B1 => n120696, B2 
                           => n120429, ZN => n6421);
   U88102 : OAI22_X1 port map( A1 => n90347, A2 => n120436, B1 => n120699, B2 
                           => n120429, ZN => n6422);
   U88103 : OAI22_X1 port map( A1 => n90346, A2 => n120436, B1 => n120702, B2 
                           => n120430, ZN => n6423);
   U88104 : OAI22_X1 port map( A1 => n90345, A2 => n120436, B1 => n120705, B2 
                           => n120430, ZN => n6424);
   U88105 : OAI22_X1 port map( A1 => n90344, A2 => n120436, B1 => n120708, B2 
                           => n120430, ZN => n6425);
   U88106 : OAI22_X1 port map( A1 => n90343, A2 => n120436, B1 => n120711, B2 
                           => n120430, ZN => n6426);
   U88107 : OAI22_X1 port map( A1 => n90342, A2 => n120436, B1 => n120714, B2 
                           => n120430, ZN => n6427);
   U88108 : OAI22_X1 port map( A1 => n90341, A2 => n120436, B1 => n120717, B2 
                           => n120430, ZN => n6428);
   U88109 : OAI22_X1 port map( A1 => n90340, A2 => n120436, B1 => n120720, B2 
                           => n120430, ZN => n6429);
   U88110 : OAI22_X1 port map( A1 => n90339, A2 => n120436, B1 => n120723, B2 
                           => n120430, ZN => n6430);
   U88111 : OAI22_X1 port map( A1 => n90338, A2 => n120436, B1 => n120726, B2 
                           => n120430, ZN => n6431);
   U88112 : OAI22_X1 port map( A1 => n90337, A2 => n120436, B1 => n120729, B2 
                           => n120430, ZN => n6432);
   U88113 : OAI22_X1 port map( A1 => n90336, A2 => n120436, B1 => n120732, B2 
                           => n120430, ZN => n6433);
   U88114 : OAI22_X1 port map( A1 => n90335, A2 => n120437, B1 => n120735, B2 
                           => n120430, ZN => n6434);
   U88115 : OAI22_X1 port map( A1 => n90334, A2 => n120437, B1 => n120738, B2 
                           => n120431, ZN => n6435);
   U88116 : OAI22_X1 port map( A1 => n90333, A2 => n120437, B1 => n120741, B2 
                           => n120431, ZN => n6436);
   U88117 : OAI22_X1 port map( A1 => n90332, A2 => n120437, B1 => n120744, B2 
                           => n120431, ZN => n6437);
   U88118 : OAI22_X1 port map( A1 => n90331, A2 => n120437, B1 => n120747, B2 
                           => n120431, ZN => n6438);
   U88119 : OAI22_X1 port map( A1 => n90330, A2 => n120437, B1 => n120750, B2 
                           => n120431, ZN => n6439);
   U88120 : OAI22_X1 port map( A1 => n90329, A2 => n120437, B1 => n120753, B2 
                           => n120431, ZN => n6440);
   U88121 : OAI22_X1 port map( A1 => n90328, A2 => n120437, B1 => n120756, B2 
                           => n120431, ZN => n6441);
   U88122 : OAI22_X1 port map( A1 => n90327, A2 => n120437, B1 => n120759, B2 
                           => n120431, ZN => n6442);
   U88123 : OAI22_X1 port map( A1 => n90326, A2 => n120437, B1 => n120762, B2 
                           => n120431, ZN => n6443);
   U88124 : OAI22_X1 port map( A1 => n90325, A2 => n120437, B1 => n120765, B2 
                           => n120431, ZN => n6444);
   U88125 : OAI22_X1 port map( A1 => n90324, A2 => n120437, B1 => n120768, B2 
                           => n120431, ZN => n6445);
   U88126 : OAI22_X1 port map( A1 => n90323, A2 => n120438, B1 => n120771, B2 
                           => n120431, ZN => n6446);
   U88127 : OAI22_X1 port map( A1 => n90322, A2 => n120438, B1 => n120774, B2 
                           => n120432, ZN => n6447);
   U88128 : OAI22_X1 port map( A1 => n90321, A2 => n120438, B1 => n120777, B2 
                           => n120432, ZN => n6448);
   U88129 : OAI22_X1 port map( A1 => n90320, A2 => n120438, B1 => n120780, B2 
                           => n120432, ZN => n6449);
   U88130 : OAI22_X1 port map( A1 => n90319, A2 => n120438, B1 => n120783, B2 
                           => n120432, ZN => n6450);
   U88131 : OAI22_X1 port map( A1 => n90318, A2 => n120438, B1 => n120786, B2 
                           => n120432, ZN => n6451);
   U88132 : OAI22_X1 port map( A1 => n90317, A2 => n120438, B1 => n120789, B2 
                           => n120432, ZN => n6452);
   U88133 : OAI22_X1 port map( A1 => n90316, A2 => n120438, B1 => n120792, B2 
                           => n120432, ZN => n6453);
   U88134 : OAI22_X1 port map( A1 => n90315, A2 => n120438, B1 => n120795, B2 
                           => n120432, ZN => n6454);
   U88135 : OAI22_X1 port map( A1 => n90314, A2 => n120438, B1 => n120798, B2 
                           => n120432, ZN => n6455);
   U88136 : OAI22_X1 port map( A1 => n90313, A2 => n120438, B1 => n120801, B2 
                           => n120432, ZN => n6456);
   U88137 : OAI22_X1 port map( A1 => n90312, A2 => n120438, B1 => n120804, B2 
                           => n120432, ZN => n6457);
   U88138 : OAI22_X1 port map( A1 => n90311, A2 => n120439, B1 => n120807, B2 
                           => n120432, ZN => n6458);
   U88139 : OAI22_X1 port map( A1 => n90437, A2 => n120422, B1 => n120630, B2 
                           => n120416, ZN => n6335);
   U88140 : OAI22_X1 port map( A1 => n90436, A2 => n120422, B1 => n120633, B2 
                           => n120416, ZN => n6336);
   U88141 : OAI22_X1 port map( A1 => n90435, A2 => n120422, B1 => n120636, B2 
                           => n120416, ZN => n6337);
   U88142 : OAI22_X1 port map( A1 => n90434, A2 => n120422, B1 => n120639, B2 
                           => n120416, ZN => n6338);
   U88143 : OAI22_X1 port map( A1 => n90433, A2 => n120422, B1 => n120642, B2 
                           => n120416, ZN => n6339);
   U88144 : OAI22_X1 port map( A1 => n90432, A2 => n120422, B1 => n120645, B2 
                           => n120416, ZN => n6340);
   U88145 : OAI22_X1 port map( A1 => n90431, A2 => n120422, B1 => n120648, B2 
                           => n120416, ZN => n6341);
   U88146 : OAI22_X1 port map( A1 => n90430, A2 => n120422, B1 => n120651, B2 
                           => n120416, ZN => n6342);
   U88147 : OAI22_X1 port map( A1 => n90429, A2 => n120422, B1 => n120654, B2 
                           => n120416, ZN => n6343);
   U88148 : OAI22_X1 port map( A1 => n90428, A2 => n120422, B1 => n120657, B2 
                           => n120416, ZN => n6344);
   U88149 : OAI22_X1 port map( A1 => n90427, A2 => n120422, B1 => n120660, B2 
                           => n120416, ZN => n6345);
   U88150 : OAI22_X1 port map( A1 => n90426, A2 => n120423, B1 => n120663, B2 
                           => n120416, ZN => n6346);
   U88151 : OAI22_X1 port map( A1 => n90425, A2 => n120423, B1 => n120666, B2 
                           => n120417, ZN => n6347);
   U88152 : OAI22_X1 port map( A1 => n90424, A2 => n120423, B1 => n120669, B2 
                           => n120417, ZN => n6348);
   U88153 : OAI22_X1 port map( A1 => n90423, A2 => n120423, B1 => n120672, B2 
                           => n120417, ZN => n6349);
   U88154 : OAI22_X1 port map( A1 => n90422, A2 => n120423, B1 => n120675, B2 
                           => n120417, ZN => n6350);
   U88155 : OAI22_X1 port map( A1 => n90421, A2 => n120423, B1 => n120678, B2 
                           => n120417, ZN => n6351);
   U88156 : OAI22_X1 port map( A1 => n90420, A2 => n120423, B1 => n120681, B2 
                           => n120417, ZN => n6352);
   U88157 : OAI22_X1 port map( A1 => n90419, A2 => n120423, B1 => n120684, B2 
                           => n120417, ZN => n6353);
   U88158 : OAI22_X1 port map( A1 => n90418, A2 => n120423, B1 => n120687, B2 
                           => n120417, ZN => n6354);
   U88159 : OAI22_X1 port map( A1 => n90417, A2 => n120423, B1 => n120690, B2 
                           => n120417, ZN => n6355);
   U88160 : OAI22_X1 port map( A1 => n90416, A2 => n120423, B1 => n120693, B2 
                           => n120417, ZN => n6356);
   U88161 : OAI22_X1 port map( A1 => n90415, A2 => n120423, B1 => n120696, B2 
                           => n120417, ZN => n6357);
   U88162 : OAI22_X1 port map( A1 => n90414, A2 => n120424, B1 => n120699, B2 
                           => n120417, ZN => n6358);
   U88163 : OAI22_X1 port map( A1 => n90413, A2 => n120424, B1 => n120702, B2 
                           => n120418, ZN => n6359);
   U88164 : OAI22_X1 port map( A1 => n90412, A2 => n120424, B1 => n120705, B2 
                           => n120418, ZN => n6360);
   U88165 : OAI22_X1 port map( A1 => n90411, A2 => n120424, B1 => n120708, B2 
                           => n120418, ZN => n6361);
   U88166 : OAI22_X1 port map( A1 => n90410, A2 => n120424, B1 => n120711, B2 
                           => n120418, ZN => n6362);
   U88167 : OAI22_X1 port map( A1 => n90409, A2 => n120424, B1 => n120714, B2 
                           => n120418, ZN => n6363);
   U88168 : OAI22_X1 port map( A1 => n90408, A2 => n120424, B1 => n120717, B2 
                           => n120418, ZN => n6364);
   U88169 : OAI22_X1 port map( A1 => n90407, A2 => n120424, B1 => n120720, B2 
                           => n120418, ZN => n6365);
   U88170 : OAI22_X1 port map( A1 => n90406, A2 => n120424, B1 => n120723, B2 
                           => n120418, ZN => n6366);
   U88171 : OAI22_X1 port map( A1 => n90405, A2 => n120424, B1 => n120726, B2 
                           => n120418, ZN => n6367);
   U88172 : OAI22_X1 port map( A1 => n90404, A2 => n120424, B1 => n120729, B2 
                           => n120418, ZN => n6368);
   U88173 : OAI22_X1 port map( A1 => n90403, A2 => n120424, B1 => n120732, B2 
                           => n120418, ZN => n6369);
   U88174 : OAI22_X1 port map( A1 => n90402, A2 => n120425, B1 => n120735, B2 
                           => n120418, ZN => n6370);
   U88175 : OAI22_X1 port map( A1 => n90401, A2 => n120425, B1 => n120738, B2 
                           => n120419, ZN => n6371);
   U88176 : OAI22_X1 port map( A1 => n90400, A2 => n120425, B1 => n120741, B2 
                           => n120419, ZN => n6372);
   U88177 : OAI22_X1 port map( A1 => n90399, A2 => n120425, B1 => n120744, B2 
                           => n120419, ZN => n6373);
   U88178 : OAI22_X1 port map( A1 => n90398, A2 => n120425, B1 => n120747, B2 
                           => n120419, ZN => n6374);
   U88179 : OAI22_X1 port map( A1 => n90397, A2 => n120425, B1 => n120750, B2 
                           => n120419, ZN => n6375);
   U88180 : OAI22_X1 port map( A1 => n90396, A2 => n120425, B1 => n120753, B2 
                           => n120419, ZN => n6376);
   U88181 : OAI22_X1 port map( A1 => n90395, A2 => n120425, B1 => n120756, B2 
                           => n120419, ZN => n6377);
   U88182 : OAI22_X1 port map( A1 => n90394, A2 => n120425, B1 => n120759, B2 
                           => n120419, ZN => n6378);
   U88183 : OAI22_X1 port map( A1 => n90393, A2 => n120425, B1 => n120762, B2 
                           => n120419, ZN => n6379);
   U88184 : OAI22_X1 port map( A1 => n90392, A2 => n120425, B1 => n120765, B2 
                           => n120419, ZN => n6380);
   U88185 : OAI22_X1 port map( A1 => n90391, A2 => n120425, B1 => n120768, B2 
                           => n120419, ZN => n6381);
   U88186 : OAI22_X1 port map( A1 => n90390, A2 => n120426, B1 => n120771, B2 
                           => n120419, ZN => n6382);
   U88187 : OAI22_X1 port map( A1 => n90389, A2 => n120426, B1 => n120774, B2 
                           => n120420, ZN => n6383);
   U88188 : OAI22_X1 port map( A1 => n90388, A2 => n120426, B1 => n120777, B2 
                           => n120420, ZN => n6384);
   U88189 : OAI22_X1 port map( A1 => n90387, A2 => n120426, B1 => n120780, B2 
                           => n120420, ZN => n6385);
   U88190 : OAI22_X1 port map( A1 => n90386, A2 => n120426, B1 => n120783, B2 
                           => n120420, ZN => n6386);
   U88191 : OAI22_X1 port map( A1 => n90385, A2 => n120426, B1 => n120786, B2 
                           => n120420, ZN => n6387);
   U88192 : OAI22_X1 port map( A1 => n90384, A2 => n120426, B1 => n120789, B2 
                           => n120420, ZN => n6388);
   U88193 : OAI22_X1 port map( A1 => n90383, A2 => n120426, B1 => n120792, B2 
                           => n120420, ZN => n6389);
   U88194 : OAI22_X1 port map( A1 => n90382, A2 => n120426, B1 => n120795, B2 
                           => n120420, ZN => n6390);
   U88195 : OAI22_X1 port map( A1 => n90381, A2 => n120426, B1 => n120798, B2 
                           => n120420, ZN => n6391);
   U88196 : OAI22_X1 port map( A1 => n90380, A2 => n120426, B1 => n120801, B2 
                           => n120420, ZN => n6392);
   U88197 : OAI22_X1 port map( A1 => n90379, A2 => n120426, B1 => n120804, B2 
                           => n120420, ZN => n6393);
   U88198 : OAI22_X1 port map( A1 => n90378, A2 => n120427, B1 => n120807, B2 
                           => n120420, ZN => n6394);
   U88199 : OAI22_X1 port map( A1 => n90775, A2 => n120348, B1 => n120630, B2 
                           => n120342, ZN => n5951);
   U88200 : OAI22_X1 port map( A1 => n90774, A2 => n120348, B1 => n120633, B2 
                           => n120342, ZN => n5952);
   U88201 : OAI22_X1 port map( A1 => n90773, A2 => n120348, B1 => n120636, B2 
                           => n120342, ZN => n5953);
   U88202 : OAI22_X1 port map( A1 => n90772, A2 => n120348, B1 => n120639, B2 
                           => n120342, ZN => n5954);
   U88203 : OAI22_X1 port map( A1 => n90771, A2 => n120348, B1 => n120642, B2 
                           => n120342, ZN => n5955);
   U88204 : OAI22_X1 port map( A1 => n90770, A2 => n120348, B1 => n120645, B2 
                           => n120342, ZN => n5956);
   U88205 : OAI22_X1 port map( A1 => n90769, A2 => n120348, B1 => n120648, B2 
                           => n120342, ZN => n5957);
   U88206 : OAI22_X1 port map( A1 => n90768, A2 => n120348, B1 => n120651, B2 
                           => n120342, ZN => n5958);
   U88207 : OAI22_X1 port map( A1 => n90767, A2 => n120348, B1 => n120654, B2 
                           => n120342, ZN => n5959);
   U88208 : OAI22_X1 port map( A1 => n90766, A2 => n120348, B1 => n120657, B2 
                           => n120342, ZN => n5960);
   U88209 : OAI22_X1 port map( A1 => n90765, A2 => n120348, B1 => n120660, B2 
                           => n120342, ZN => n5961);
   U88210 : OAI22_X1 port map( A1 => n90764, A2 => n120349, B1 => n120663, B2 
                           => n120342, ZN => n5962);
   U88211 : OAI22_X1 port map( A1 => n90763, A2 => n120349, B1 => n120666, B2 
                           => n120343, ZN => n5963);
   U88212 : OAI22_X1 port map( A1 => n90762, A2 => n120349, B1 => n120669, B2 
                           => n120343, ZN => n5964);
   U88213 : OAI22_X1 port map( A1 => n90761, A2 => n120349, B1 => n120672, B2 
                           => n120343, ZN => n5965);
   U88214 : OAI22_X1 port map( A1 => n90760, A2 => n120349, B1 => n120675, B2 
                           => n120343, ZN => n5966);
   U88215 : OAI22_X1 port map( A1 => n90759, A2 => n120349, B1 => n120678, B2 
                           => n120343, ZN => n5967);
   U88216 : OAI22_X1 port map( A1 => n90758, A2 => n120349, B1 => n120681, B2 
                           => n120343, ZN => n5968);
   U88217 : OAI22_X1 port map( A1 => n90757, A2 => n120349, B1 => n120684, B2 
                           => n120343, ZN => n5969);
   U88218 : OAI22_X1 port map( A1 => n90756, A2 => n120349, B1 => n120687, B2 
                           => n120343, ZN => n5970);
   U88219 : OAI22_X1 port map( A1 => n90755, A2 => n120349, B1 => n120690, B2 
                           => n120343, ZN => n5971);
   U88220 : OAI22_X1 port map( A1 => n90754, A2 => n120349, B1 => n120693, B2 
                           => n120343, ZN => n5972);
   U88221 : OAI22_X1 port map( A1 => n90753, A2 => n120349, B1 => n120696, B2 
                           => n120343, ZN => n5973);
   U88222 : OAI22_X1 port map( A1 => n90752, A2 => n120350, B1 => n120699, B2 
                           => n120343, ZN => n5974);
   U88223 : OAI22_X1 port map( A1 => n90751, A2 => n120350, B1 => n120702, B2 
                           => n120344, ZN => n5975);
   U88224 : OAI22_X1 port map( A1 => n90750, A2 => n120350, B1 => n120705, B2 
                           => n120344, ZN => n5976);
   U88225 : OAI22_X1 port map( A1 => n90749, A2 => n120350, B1 => n120708, B2 
                           => n120344, ZN => n5977);
   U88226 : OAI22_X1 port map( A1 => n90748, A2 => n120350, B1 => n120711, B2 
                           => n120344, ZN => n5978);
   U88227 : OAI22_X1 port map( A1 => n90747, A2 => n120350, B1 => n120714, B2 
                           => n120344, ZN => n5979);
   U88228 : OAI22_X1 port map( A1 => n90746, A2 => n120350, B1 => n120717, B2 
                           => n120344, ZN => n5980);
   U88229 : OAI22_X1 port map( A1 => n90745, A2 => n120350, B1 => n120720, B2 
                           => n120344, ZN => n5981);
   U88230 : OAI22_X1 port map( A1 => n90744, A2 => n120350, B1 => n120723, B2 
                           => n120344, ZN => n5982);
   U88231 : OAI22_X1 port map( A1 => n90743, A2 => n120350, B1 => n120726, B2 
                           => n120344, ZN => n5983);
   U88232 : OAI22_X1 port map( A1 => n90742, A2 => n120350, B1 => n120729, B2 
                           => n120344, ZN => n5984);
   U88233 : OAI22_X1 port map( A1 => n90741, A2 => n120350, B1 => n120732, B2 
                           => n120344, ZN => n5985);
   U88234 : OAI22_X1 port map( A1 => n90740, A2 => n120351, B1 => n120735, B2 
                           => n120344, ZN => n5986);
   U88235 : OAI22_X1 port map( A1 => n90739, A2 => n120351, B1 => n120738, B2 
                           => n120345, ZN => n5987);
   U88236 : OAI22_X1 port map( A1 => n90738, A2 => n120351, B1 => n120741, B2 
                           => n120345, ZN => n5988);
   U88237 : OAI22_X1 port map( A1 => n90737, A2 => n120351, B1 => n120744, B2 
                           => n120345, ZN => n5989);
   U88238 : OAI22_X1 port map( A1 => n90736, A2 => n120351, B1 => n120747, B2 
                           => n120345, ZN => n5990);
   U88239 : OAI22_X1 port map( A1 => n90735, A2 => n120351, B1 => n120750, B2 
                           => n120345, ZN => n5991);
   U88240 : OAI22_X1 port map( A1 => n90734, A2 => n120351, B1 => n120753, B2 
                           => n120345, ZN => n5992);
   U88241 : OAI22_X1 port map( A1 => n90733, A2 => n120351, B1 => n120756, B2 
                           => n120345, ZN => n5993);
   U88242 : OAI22_X1 port map( A1 => n90732, A2 => n120351, B1 => n120759, B2 
                           => n120345, ZN => n5994);
   U88243 : OAI22_X1 port map( A1 => n90731, A2 => n120351, B1 => n120762, B2 
                           => n120345, ZN => n5995);
   U88244 : OAI22_X1 port map( A1 => n90730, A2 => n120351, B1 => n120765, B2 
                           => n120345, ZN => n5996);
   U88245 : OAI22_X1 port map( A1 => n90729, A2 => n120351, B1 => n120768, B2 
                           => n120345, ZN => n5997);
   U88246 : OAI22_X1 port map( A1 => n90728, A2 => n120352, B1 => n120771, B2 
                           => n120345, ZN => n5998);
   U88247 : OAI22_X1 port map( A1 => n90727, A2 => n120352, B1 => n120774, B2 
                           => n120346, ZN => n5999);
   U88248 : OAI22_X1 port map( A1 => n90726, A2 => n120352, B1 => n120777, B2 
                           => n120346, ZN => n6000);
   U88249 : OAI22_X1 port map( A1 => n90725, A2 => n120352, B1 => n120780, B2 
                           => n120346, ZN => n6001);
   U88250 : OAI22_X1 port map( A1 => n90724, A2 => n120352, B1 => n120783, B2 
                           => n120346, ZN => n6002);
   U88251 : OAI22_X1 port map( A1 => n90723, A2 => n120352, B1 => n120786, B2 
                           => n120346, ZN => n6003);
   U88252 : OAI22_X1 port map( A1 => n90722, A2 => n120352, B1 => n120789, B2 
                           => n120346, ZN => n6004);
   U88253 : OAI22_X1 port map( A1 => n90721, A2 => n120352, B1 => n120792, B2 
                           => n120346, ZN => n6005);
   U88254 : OAI22_X1 port map( A1 => n90720, A2 => n120352, B1 => n120795, B2 
                           => n120346, ZN => n6006);
   U88255 : OAI22_X1 port map( A1 => n90719, A2 => n120352, B1 => n120798, B2 
                           => n120346, ZN => n6007);
   U88256 : OAI22_X1 port map( A1 => n90718, A2 => n120352, B1 => n120801, B2 
                           => n120346, ZN => n6008);
   U88257 : OAI22_X1 port map( A1 => n90717, A2 => n120352, B1 => n120804, B2 
                           => n120346, ZN => n6009);
   U88258 : OAI22_X1 port map( A1 => n90716, A2 => n120353, B1 => n120807, B2 
                           => n120346, ZN => n6010);
   U88259 : OAI22_X1 port map( A1 => n90095, A2 => n120531, B1 => n120629, B2 
                           => n120525, ZN => n6911);
   U88260 : OAI22_X1 port map( A1 => n90094, A2 => n120531, B1 => n120632, B2 
                           => n120525, ZN => n6912);
   U88261 : OAI22_X1 port map( A1 => n90093, A2 => n120531, B1 => n120635, B2 
                           => n120525, ZN => n6913);
   U88262 : OAI22_X1 port map( A1 => n90092, A2 => n120531, B1 => n120638, B2 
                           => n120525, ZN => n6914);
   U88263 : OAI22_X1 port map( A1 => n90091, A2 => n120531, B1 => n120641, B2 
                           => n120525, ZN => n6915);
   U88264 : OAI22_X1 port map( A1 => n90090, A2 => n120531, B1 => n120644, B2 
                           => n120525, ZN => n6916);
   U88265 : OAI22_X1 port map( A1 => n90089, A2 => n120531, B1 => n120647, B2 
                           => n120525, ZN => n6917);
   U88266 : OAI22_X1 port map( A1 => n90088, A2 => n120531, B1 => n120650, B2 
                           => n120525, ZN => n6918);
   U88267 : OAI22_X1 port map( A1 => n90087, A2 => n120531, B1 => n120653, B2 
                           => n120525, ZN => n6919);
   U88268 : OAI22_X1 port map( A1 => n90086, A2 => n120531, B1 => n120656, B2 
                           => n120525, ZN => n6920);
   U88269 : OAI22_X1 port map( A1 => n90085, A2 => n120531, B1 => n120659, B2 
                           => n120525, ZN => n6921);
   U88270 : OAI22_X1 port map( A1 => n90084, A2 => n120532, B1 => n120662, B2 
                           => n120525, ZN => n6922);
   U88271 : OAI22_X1 port map( A1 => n90083, A2 => n120532, B1 => n120665, B2 
                           => n120526, ZN => n6923);
   U88272 : OAI22_X1 port map( A1 => n90082, A2 => n120532, B1 => n120668, B2 
                           => n120526, ZN => n6924);
   U88273 : OAI22_X1 port map( A1 => n90081, A2 => n120532, B1 => n120671, B2 
                           => n120526, ZN => n6925);
   U88274 : OAI22_X1 port map( A1 => n90080, A2 => n120532, B1 => n120674, B2 
                           => n120526, ZN => n6926);
   U88275 : OAI22_X1 port map( A1 => n90079, A2 => n120532, B1 => n120677, B2 
                           => n120526, ZN => n6927);
   U88276 : OAI22_X1 port map( A1 => n90078, A2 => n120532, B1 => n120680, B2 
                           => n120526, ZN => n6928);
   U88277 : OAI22_X1 port map( A1 => n90077, A2 => n120532, B1 => n120683, B2 
                           => n120526, ZN => n6929);
   U88278 : OAI22_X1 port map( A1 => n90076, A2 => n120532, B1 => n120686, B2 
                           => n120526, ZN => n6930);
   U88279 : OAI22_X1 port map( A1 => n90075, A2 => n120532, B1 => n120689, B2 
                           => n120526, ZN => n6931);
   U88280 : OAI22_X1 port map( A1 => n90074, A2 => n120532, B1 => n120692, B2 
                           => n120526, ZN => n6932);
   U88281 : OAI22_X1 port map( A1 => n90073, A2 => n120532, B1 => n120695, B2 
                           => n120526, ZN => n6933);
   U88282 : OAI22_X1 port map( A1 => n90072, A2 => n120533, B1 => n120698, B2 
                           => n120526, ZN => n6934);
   U88283 : OAI22_X1 port map( A1 => n90071, A2 => n120533, B1 => n120701, B2 
                           => n120527, ZN => n6935);
   U88284 : OAI22_X1 port map( A1 => n90070, A2 => n120533, B1 => n120704, B2 
                           => n120527, ZN => n6936);
   U88285 : OAI22_X1 port map( A1 => n90069, A2 => n120533, B1 => n120707, B2 
                           => n120527, ZN => n6937);
   U88286 : OAI22_X1 port map( A1 => n90068, A2 => n120533, B1 => n120710, B2 
                           => n120527, ZN => n6938);
   U88287 : OAI22_X1 port map( A1 => n90067, A2 => n120533, B1 => n120713, B2 
                           => n120527, ZN => n6939);
   U88288 : OAI22_X1 port map( A1 => n90066, A2 => n120533, B1 => n120716, B2 
                           => n120527, ZN => n6940);
   U88289 : OAI22_X1 port map( A1 => n90065, A2 => n120533, B1 => n120719, B2 
                           => n120527, ZN => n6941);
   U88290 : OAI22_X1 port map( A1 => n90064, A2 => n120533, B1 => n120722, B2 
                           => n120527, ZN => n6942);
   U88291 : OAI22_X1 port map( A1 => n90063, A2 => n120533, B1 => n120725, B2 
                           => n120527, ZN => n6943);
   U88292 : OAI22_X1 port map( A1 => n90062, A2 => n120533, B1 => n120728, B2 
                           => n120527, ZN => n6944);
   U88293 : OAI22_X1 port map( A1 => n90061, A2 => n120533, B1 => n120731, B2 
                           => n120527, ZN => n6945);
   U88294 : OAI22_X1 port map( A1 => n90060, A2 => n120534, B1 => n120734, B2 
                           => n120527, ZN => n6946);
   U88295 : OAI22_X1 port map( A1 => n90059, A2 => n120534, B1 => n120737, B2 
                           => n120528, ZN => n6947);
   U88296 : OAI22_X1 port map( A1 => n90058, A2 => n120534, B1 => n120740, B2 
                           => n120528, ZN => n6948);
   U88297 : OAI22_X1 port map( A1 => n90057, A2 => n120534, B1 => n120743, B2 
                           => n120528, ZN => n6949);
   U88298 : OAI22_X1 port map( A1 => n90056, A2 => n120534, B1 => n120746, B2 
                           => n120528, ZN => n6950);
   U88299 : OAI22_X1 port map( A1 => n90055, A2 => n120534, B1 => n120749, B2 
                           => n120528, ZN => n6951);
   U88300 : OAI22_X1 port map( A1 => n90054, A2 => n120534, B1 => n120752, B2 
                           => n120528, ZN => n6952);
   U88301 : OAI22_X1 port map( A1 => n90053, A2 => n120534, B1 => n120755, B2 
                           => n120528, ZN => n6953);
   U88302 : OAI22_X1 port map( A1 => n90052, A2 => n120534, B1 => n120758, B2 
                           => n120528, ZN => n6954);
   U88303 : OAI22_X1 port map( A1 => n90051, A2 => n120534, B1 => n120761, B2 
                           => n120528, ZN => n6955);
   U88304 : OAI22_X1 port map( A1 => n90050, A2 => n120534, B1 => n120764, B2 
                           => n120528, ZN => n6956);
   U88305 : OAI22_X1 port map( A1 => n90049, A2 => n120534, B1 => n120767, B2 
                           => n120528, ZN => n6957);
   U88306 : OAI22_X1 port map( A1 => n90048, A2 => n120535, B1 => n120770, B2 
                           => n120528, ZN => n6958);
   U88307 : OAI22_X1 port map( A1 => n90047, A2 => n120535, B1 => n120773, B2 
                           => n120529, ZN => n6959);
   U88308 : OAI22_X1 port map( A1 => n90046, A2 => n120535, B1 => n120776, B2 
                           => n120529, ZN => n6960);
   U88309 : OAI22_X1 port map( A1 => n90045, A2 => n120535, B1 => n120779, B2 
                           => n120529, ZN => n6961);
   U88310 : OAI22_X1 port map( A1 => n90044, A2 => n120535, B1 => n120782, B2 
                           => n120529, ZN => n6962);
   U88311 : OAI22_X1 port map( A1 => n90043, A2 => n120535, B1 => n120785, B2 
                           => n120529, ZN => n6963);
   U88312 : OAI22_X1 port map( A1 => n90042, A2 => n120535, B1 => n120788, B2 
                           => n120529, ZN => n6964);
   U88313 : OAI22_X1 port map( A1 => n90041, A2 => n120535, B1 => n120791, B2 
                           => n120529, ZN => n6965);
   U88314 : OAI22_X1 port map( A1 => n90040, A2 => n120535, B1 => n120794, B2 
                           => n120529, ZN => n6966);
   U88315 : OAI22_X1 port map( A1 => n90039, A2 => n120535, B1 => n120797, B2 
                           => n120529, ZN => n6967);
   U88316 : OAI22_X1 port map( A1 => n90038, A2 => n120535, B1 => n120800, B2 
                           => n120529, ZN => n6968);
   U88317 : OAI22_X1 port map( A1 => n90037, A2 => n120535, B1 => n120803, B2 
                           => n120529, ZN => n6969);
   U88318 : OAI22_X1 port map( A1 => n90036, A2 => n120536, B1 => n120806, B2 
                           => n120529, ZN => n6970);
   U88319 : INV_X1 port map( A => ADD_RD2(3), ZN => n117958);
   U88320 : INV_X1 port map( A => ADD_RD1(4), ZN => n116471);
   U88321 : INV_X1 port map( A => ADD_RD2(0), ZN => n117967);
   U88322 : INV_X1 port map( A => ADD_RD1(3), ZN => n116470);
   U88323 : INV_X1 port map( A => ADD_RD2(4), ZN => n117970);
   U88324 : INV_X1 port map( A => ADD_RD1(0), ZN => n116469);
   U88325 : NAND4_X1 port map( A1 => n117693, A2 => n117694, A3 => n117695, A4 
                           => n117696, ZN => n5322);
   U88326 : AOI221_X1 port map( B1 => n119886, B2 => n118798, C1 => n119880, C2
                           => n109990, A => n117713, ZN => n117694);
   U88327 : AOI221_X1 port map( B1 => n119862, B2 => n95440, C1 => n119856, C2 
                           => n118396, A => n117714, ZN => n117693);
   U88328 : NOR4_X1 port map( A1 => n117709, A2 => n117710, A3 => n117711, A4 
                           => n117712, ZN => n117695);
   U88329 : NAND4_X1 port map( A1 => n117671, A2 => n117672, A3 => n117673, A4 
                           => n117674, ZN => n5323);
   U88330 : AOI221_X1 port map( B1 => n119887, B2 => n118799, C1 => n119881, C2
                           => n109991, A => n117691, ZN => n117672);
   U88331 : AOI221_X1 port map( B1 => n119863, B2 => n95441, C1 => n119857, C2 
                           => n118397, A => n117692, ZN => n117671);
   U88332 : NOR4_X1 port map( A1 => n117687, A2 => n117688, A3 => n117689, A4 
                           => n117690, ZN => n117673);
   U88333 : NAND4_X1 port map( A1 => n117649, A2 => n117650, A3 => n117651, A4 
                           => n117652, ZN => n5324);
   U88334 : AOI221_X1 port map( B1 => n119887, B2 => n118800, C1 => n119881, C2
                           => n109992, A => n117669, ZN => n117650);
   U88335 : AOI221_X1 port map( B1 => n119863, B2 => n95442, C1 => n119857, C2 
                           => n118398, A => n117670, ZN => n117649);
   U88336 : NOR4_X1 port map( A1 => n117665, A2 => n117666, A3 => n117667, A4 
                           => n117668, ZN => n117651);
   U88337 : NAND4_X1 port map( A1 => n117627, A2 => n117628, A3 => n117629, A4 
                           => n117630, ZN => n5325);
   U88338 : AOI221_X1 port map( B1 => n119887, B2 => n118801, C1 => n119881, C2
                           => n109993, A => n117647, ZN => n117628);
   U88339 : AOI221_X1 port map( B1 => n119863, B2 => n95443, C1 => n119857, C2 
                           => n118399, A => n117648, ZN => n117627);
   U88340 : NOR4_X1 port map( A1 => n117643, A2 => n117644, A3 => n117645, A4 
                           => n117646, ZN => n117629);
   U88341 : NAND4_X1 port map( A1 => n117605, A2 => n117606, A3 => n117607, A4 
                           => n117608, ZN => n5326);
   U88342 : AOI221_X1 port map( B1 => n119887, B2 => n118802, C1 => n119881, C2
                           => n109994, A => n117625, ZN => n117606);
   U88343 : AOI221_X1 port map( B1 => n119863, B2 => n95444, C1 => n119857, C2 
                           => n118400, A => n117626, ZN => n117605);
   U88344 : NOR4_X1 port map( A1 => n117621, A2 => n117622, A3 => n117623, A4 
                           => n117624, ZN => n117607);
   U88345 : NAND4_X1 port map( A1 => n117583, A2 => n117584, A3 => n117585, A4 
                           => n117586, ZN => n5327);
   U88346 : AOI221_X1 port map( B1 => n119887, B2 => n118803, C1 => n119881, C2
                           => n109995, A => n117603, ZN => n117584);
   U88347 : AOI221_X1 port map( B1 => n119863, B2 => n95445, C1 => n119857, C2 
                           => n118401, A => n117604, ZN => n117583);
   U88348 : NOR4_X1 port map( A1 => n117599, A2 => n117600, A3 => n117601, A4 
                           => n117602, ZN => n117585);
   U88349 : NAND4_X1 port map( A1 => n117561, A2 => n117562, A3 => n117563, A4 
                           => n117564, ZN => n5328);
   U88350 : AOI221_X1 port map( B1 => n119887, B2 => n118804, C1 => n119881, C2
                           => n109996, A => n117581, ZN => n117562);
   U88351 : AOI221_X1 port map( B1 => n119863, B2 => n95446, C1 => n119857, C2 
                           => n118402, A => n117582, ZN => n117561);
   U88352 : NOR4_X1 port map( A1 => n117577, A2 => n117578, A3 => n117579, A4 
                           => n117580, ZN => n117563);
   U88353 : NAND4_X1 port map( A1 => n117539, A2 => n117540, A3 => n117541, A4 
                           => n117542, ZN => n5329);
   U88354 : AOI221_X1 port map( B1 => n119887, B2 => n118805, C1 => n119881, C2
                           => n109997, A => n117559, ZN => n117540);
   U88355 : AOI221_X1 port map( B1 => n119863, B2 => n95447, C1 => n119857, C2 
                           => n118403, A => n117560, ZN => n117539);
   U88356 : NOR4_X1 port map( A1 => n117555, A2 => n117556, A3 => n117557, A4 
                           => n117558, ZN => n117541);
   U88357 : NAND4_X1 port map( A1 => n117516, A2 => n117517, A3 => n117518, A4 
                           => n117519, ZN => n5330);
   U88358 : AOI221_X1 port map( B1 => n119887, B2 => n118505, C1 => n119881, C2
                           => n118817, A => n117537, ZN => n117517);
   U88359 : AOI221_X1 port map( B1 => n119863, B2 => n95448, C1 => n119857, C2 
                           => n118404, A => n117538, ZN => n117516);
   U88360 : NOR4_X1 port map( A1 => n117532, A2 => n117533, A3 => n117534, A4 
                           => n117535, ZN => n117518);
   U88361 : NAND4_X1 port map( A1 => n117493, A2 => n117494, A3 => n117495, A4 
                           => n117496, ZN => n5331);
   U88362 : AOI221_X1 port map( B1 => n119887, B2 => n118506, C1 => n119881, C2
                           => n118818, A => n117514, ZN => n117494);
   U88363 : AOI221_X1 port map( B1 => n119863, B2 => n95449, C1 => n119857, C2 
                           => n118405, A => n117515, ZN => n117493);
   U88364 : NOR4_X1 port map( A1 => n117509, A2 => n117510, A3 => n117511, A4 
                           => n117512, ZN => n117495);
   U88365 : NAND4_X1 port map( A1 => n117470, A2 => n117471, A3 => n117472, A4 
                           => n117473, ZN => n5332);
   U88366 : AOI221_X1 port map( B1 => n119887, B2 => n118507, C1 => n119881, C2
                           => n118819, A => n117491, ZN => n117471);
   U88367 : AOI221_X1 port map( B1 => n119863, B2 => n95450, C1 => n119857, C2 
                           => n118406, A => n117492, ZN => n117470);
   U88368 : NOR4_X1 port map( A1 => n117486, A2 => n117487, A3 => n117488, A4 
                           => n117489, ZN => n117472);
   U88369 : NAND4_X1 port map( A1 => n117447, A2 => n117448, A3 => n117449, A4 
                           => n117450, ZN => n5333);
   U88370 : AOI221_X1 port map( B1 => n119887, B2 => n118508, C1 => n119881, C2
                           => n118820, A => n117468, ZN => n117448);
   U88371 : AOI221_X1 port map( B1 => n119863, B2 => n95451, C1 => n119857, C2 
                           => n118407, A => n117469, ZN => n117447);
   U88372 : NOR4_X1 port map( A1 => n117463, A2 => n117464, A3 => n117465, A4 
                           => n117466, ZN => n117449);
   U88373 : NAND4_X1 port map( A1 => n117424, A2 => n117425, A3 => n117426, A4 
                           => n117427, ZN => n5334);
   U88374 : AOI221_X1 port map( B1 => n119887, B2 => n118509, C1 => n119881, C2
                           => n118821, A => n117445, ZN => n117425);
   U88375 : AOI221_X1 port map( B1 => n119863, B2 => n95452, C1 => n119857, C2 
                           => n118408, A => n117446, ZN => n117424);
   U88376 : NOR4_X1 port map( A1 => n117440, A2 => n117441, A3 => n117442, A4 
                           => n117443, ZN => n117426);
   U88377 : NAND4_X1 port map( A1 => n117401, A2 => n117402, A3 => n117403, A4 
                           => n117404, ZN => n5335);
   U88378 : AOI221_X1 port map( B1 => n119888, B2 => n118510, C1 => n119882, C2
                           => n118822, A => n117422, ZN => n117402);
   U88379 : AOI221_X1 port map( B1 => n119864, B2 => n95453, C1 => n119858, C2 
                           => n118409, A => n117423, ZN => n117401);
   U88380 : NOR4_X1 port map( A1 => n117417, A2 => n117418, A3 => n117419, A4 
                           => n117420, ZN => n117403);
   U88381 : NAND4_X1 port map( A1 => n117378, A2 => n117379, A3 => n117380, A4 
                           => n117381, ZN => n5336);
   U88382 : AOI221_X1 port map( B1 => n119888, B2 => n118511, C1 => n119882, C2
                           => n118823, A => n117399, ZN => n117379);
   U88383 : AOI221_X1 port map( B1 => n119864, B2 => n95454, C1 => n119858, C2 
                           => n118410, A => n117400, ZN => n117378);
   U88384 : NOR4_X1 port map( A1 => n117394, A2 => n117395, A3 => n117396, A4 
                           => n117397, ZN => n117380);
   U88385 : NAND4_X1 port map( A1 => n117355, A2 => n117356, A3 => n117357, A4 
                           => n117358, ZN => n5337);
   U88386 : AOI221_X1 port map( B1 => n119888, B2 => n118512, C1 => n119882, C2
                           => n118824, A => n117376, ZN => n117356);
   U88387 : AOI221_X1 port map( B1 => n119864, B2 => n95455, C1 => n119858, C2 
                           => n118411, A => n117377, ZN => n117355);
   U88388 : NOR4_X1 port map( A1 => n117371, A2 => n117372, A3 => n117373, A4 
                           => n117374, ZN => n117357);
   U88389 : NAND4_X1 port map( A1 => n117332, A2 => n117333, A3 => n117334, A4 
                           => n117335, ZN => n5338);
   U88390 : AOI221_X1 port map( B1 => n119888, B2 => n118513, C1 => n119882, C2
                           => n118825, A => n117353, ZN => n117333);
   U88391 : AOI221_X1 port map( B1 => n119864, B2 => n95456, C1 => n119858, C2 
                           => n118412, A => n117354, ZN => n117332);
   U88392 : NOR4_X1 port map( A1 => n117348, A2 => n117349, A3 => n117350, A4 
                           => n117351, ZN => n117334);
   U88393 : NAND4_X1 port map( A1 => n117309, A2 => n117310, A3 => n117311, A4 
                           => n117312, ZN => n5339);
   U88394 : AOI221_X1 port map( B1 => n119888, B2 => n118514, C1 => n119882, C2
                           => n118826, A => n117330, ZN => n117310);
   U88395 : AOI221_X1 port map( B1 => n119864, B2 => n95457, C1 => n119858, C2 
                           => n118413, A => n117331, ZN => n117309);
   U88396 : NOR4_X1 port map( A1 => n117325, A2 => n117326, A3 => n117327, A4 
                           => n117328, ZN => n117311);
   U88397 : NAND4_X1 port map( A1 => n117286, A2 => n117287, A3 => n117288, A4 
                           => n117289, ZN => n5340);
   U88398 : AOI221_X1 port map( B1 => n119888, B2 => n118515, C1 => n119882, C2
                           => n118827, A => n117307, ZN => n117287);
   U88399 : AOI221_X1 port map( B1 => n119864, B2 => n95458, C1 => n119858, C2 
                           => n118414, A => n117308, ZN => n117286);
   U88400 : NOR4_X1 port map( A1 => n117302, A2 => n117303, A3 => n117304, A4 
                           => n117305, ZN => n117288);
   U88401 : NAND4_X1 port map( A1 => n117263, A2 => n117264, A3 => n117265, A4 
                           => n117266, ZN => n5341);
   U88402 : AOI221_X1 port map( B1 => n119888, B2 => n118516, C1 => n119882, C2
                           => n118828, A => n117284, ZN => n117264);
   U88403 : AOI221_X1 port map( B1 => n119864, B2 => n95459, C1 => n119858, C2 
                           => n118415, A => n117285, ZN => n117263);
   U88404 : NOR4_X1 port map( A1 => n117279, A2 => n117280, A3 => n117281, A4 
                           => n117282, ZN => n117265);
   U88405 : NAND4_X1 port map( A1 => n117240, A2 => n117241, A3 => n117242, A4 
                           => n117243, ZN => n5342);
   U88406 : AOI221_X1 port map( B1 => n119888, B2 => n118517, C1 => n119882, C2
                           => n118829, A => n117261, ZN => n117241);
   U88407 : AOI221_X1 port map( B1 => n119864, B2 => n95460, C1 => n119858, C2 
                           => n118416, A => n117262, ZN => n117240);
   U88408 : NOR4_X1 port map( A1 => n117256, A2 => n117257, A3 => n117258, A4 
                           => n117259, ZN => n117242);
   U88409 : NAND4_X1 port map( A1 => n117217, A2 => n117218, A3 => n117219, A4 
                           => n117220, ZN => n5343);
   U88410 : AOI221_X1 port map( B1 => n119888, B2 => n118518, C1 => n119882, C2
                           => n118830, A => n117238, ZN => n117218);
   U88411 : AOI221_X1 port map( B1 => n119864, B2 => n95461, C1 => n119858, C2 
                           => n118417, A => n117239, ZN => n117217);
   U88412 : NOR4_X1 port map( A1 => n117233, A2 => n117234, A3 => n117235, A4 
                           => n117236, ZN => n117219);
   U88413 : NAND4_X1 port map( A1 => n117194, A2 => n117195, A3 => n117196, A4 
                           => n117197, ZN => n5344);
   U88414 : AOI221_X1 port map( B1 => n119888, B2 => n118519, C1 => n119882, C2
                           => n118831, A => n117215, ZN => n117195);
   U88415 : AOI221_X1 port map( B1 => n119864, B2 => n95462, C1 => n119858, C2 
                           => n118418, A => n117216, ZN => n117194);
   U88416 : NOR4_X1 port map( A1 => n117210, A2 => n117211, A3 => n117212, A4 
                           => n117213, ZN => n117196);
   U88417 : NAND4_X1 port map( A1 => n117171, A2 => n117172, A3 => n117173, A4 
                           => n117174, ZN => n5345);
   U88418 : AOI221_X1 port map( B1 => n119888, B2 => n118520, C1 => n119882, C2
                           => n118832, A => n117192, ZN => n117172);
   U88419 : AOI221_X1 port map( B1 => n119864, B2 => n95463, C1 => n119858, C2 
                           => n118419, A => n117193, ZN => n117171);
   U88420 : NOR4_X1 port map( A1 => n117187, A2 => n117188, A3 => n117189, A4 
                           => n117190, ZN => n117173);
   U88421 : NAND4_X1 port map( A1 => n117148, A2 => n117149, A3 => n117150, A4 
                           => n117151, ZN => n5346);
   U88422 : AOI221_X1 port map( B1 => n119888, B2 => n118521, C1 => n119882, C2
                           => n118833, A => n117169, ZN => n117149);
   U88423 : AOI221_X1 port map( B1 => n119864, B2 => n95464, C1 => n119858, C2 
                           => n118420, A => n117170, ZN => n117148);
   U88424 : NOR4_X1 port map( A1 => n117164, A2 => n117165, A3 => n117166, A4 
                           => n117167, ZN => n117150);
   U88425 : NAND4_X1 port map( A1 => n117125, A2 => n117126, A3 => n117127, A4 
                           => n117128, ZN => n5347);
   U88426 : AOI221_X1 port map( B1 => n119889, B2 => n118522, C1 => n119883, C2
                           => n118834, A => n117146, ZN => n117126);
   U88427 : AOI221_X1 port map( B1 => n119865, B2 => n95465, C1 => n119859, C2 
                           => n118421, A => n117147, ZN => n117125);
   U88428 : NOR4_X1 port map( A1 => n117141, A2 => n117142, A3 => n117143, A4 
                           => n117144, ZN => n117127);
   U88429 : NAND4_X1 port map( A1 => n117102, A2 => n117103, A3 => n117104, A4 
                           => n117105, ZN => n5348);
   U88430 : AOI221_X1 port map( B1 => n119889, B2 => n118523, C1 => n119883, C2
                           => n118835, A => n117123, ZN => n117103);
   U88431 : AOI221_X1 port map( B1 => n119865, B2 => n95466, C1 => n119859, C2 
                           => n118422, A => n117124, ZN => n117102);
   U88432 : NOR4_X1 port map( A1 => n117118, A2 => n117119, A3 => n117120, A4 
                           => n117121, ZN => n117104);
   U88433 : NAND4_X1 port map( A1 => n117079, A2 => n117080, A3 => n117081, A4 
                           => n117082, ZN => n5349);
   U88434 : AOI221_X1 port map( B1 => n119889, B2 => n118524, C1 => n119883, C2
                           => n118836, A => n117100, ZN => n117080);
   U88435 : AOI221_X1 port map( B1 => n119865, B2 => n95467, C1 => n119859, C2 
                           => n118423, A => n117101, ZN => n117079);
   U88436 : NOR4_X1 port map( A1 => n117095, A2 => n117096, A3 => n117097, A4 
                           => n117098, ZN => n117081);
   U88437 : NAND4_X1 port map( A1 => n117056, A2 => n117057, A3 => n117058, A4 
                           => n117059, ZN => n5350);
   U88438 : AOI221_X1 port map( B1 => n119889, B2 => n118525, C1 => n119883, C2
                           => n118837, A => n117077, ZN => n117057);
   U88439 : AOI221_X1 port map( B1 => n119865, B2 => n95468, C1 => n119859, C2 
                           => n118424, A => n117078, ZN => n117056);
   U88440 : NOR4_X1 port map( A1 => n117072, A2 => n117073, A3 => n117074, A4 
                           => n117075, ZN => n117058);
   U88441 : NAND4_X1 port map( A1 => n117033, A2 => n117034, A3 => n117035, A4 
                           => n117036, ZN => n5351);
   U88442 : AOI221_X1 port map( B1 => n119889, B2 => n118526, C1 => n119883, C2
                           => n118838, A => n117054, ZN => n117034);
   U88443 : AOI221_X1 port map( B1 => n119865, B2 => n95469, C1 => n119859, C2 
                           => n118425, A => n117055, ZN => n117033);
   U88444 : NOR4_X1 port map( A1 => n117049, A2 => n117050, A3 => n117051, A4 
                           => n117052, ZN => n117035);
   U88445 : NAND4_X1 port map( A1 => n117010, A2 => n117011, A3 => n117012, A4 
                           => n117013, ZN => n5352);
   U88446 : AOI221_X1 port map( B1 => n119889, B2 => n118527, C1 => n119883, C2
                           => n118839, A => n117031, ZN => n117011);
   U88447 : AOI221_X1 port map( B1 => n119865, B2 => n95470, C1 => n119859, C2 
                           => n118426, A => n117032, ZN => n117010);
   U88448 : NOR4_X1 port map( A1 => n117026, A2 => n117027, A3 => n117028, A4 
                           => n117029, ZN => n117012);
   U88449 : NAND4_X1 port map( A1 => n116987, A2 => n116988, A3 => n116989, A4 
                           => n116990, ZN => n5353);
   U88450 : AOI221_X1 port map( B1 => n119889, B2 => n118528, C1 => n119883, C2
                           => n118840, A => n117008, ZN => n116988);
   U88451 : AOI221_X1 port map( B1 => n119865, B2 => n95471, C1 => n119859, C2 
                           => n118427, A => n117009, ZN => n116987);
   U88452 : NOR4_X1 port map( A1 => n117003, A2 => n117004, A3 => n117005, A4 
                           => n117006, ZN => n116989);
   U88453 : NAND4_X1 port map( A1 => n116964, A2 => n116965, A3 => n116966, A4 
                           => n116967, ZN => n5354);
   U88454 : AOI221_X1 port map( B1 => n119889, B2 => n118529, C1 => n119883, C2
                           => n118841, A => n116985, ZN => n116965);
   U88455 : AOI221_X1 port map( B1 => n119865, B2 => n95472, C1 => n119859, C2 
                           => n118428, A => n116986, ZN => n116964);
   U88456 : NOR4_X1 port map( A1 => n116980, A2 => n116981, A3 => n116982, A4 
                           => n116983, ZN => n116966);
   U88457 : NAND4_X1 port map( A1 => n116941, A2 => n116942, A3 => n116943, A4 
                           => n116944, ZN => n5355);
   U88458 : AOI221_X1 port map( B1 => n119889, B2 => n118530, C1 => n119883, C2
                           => n118842, A => n116962, ZN => n116942);
   U88459 : AOI221_X1 port map( B1 => n119865, B2 => n95473, C1 => n119859, C2 
                           => n118429, A => n116963, ZN => n116941);
   U88460 : NOR4_X1 port map( A1 => n116957, A2 => n116958, A3 => n116959, A4 
                           => n116960, ZN => n116943);
   U88461 : NAND4_X1 port map( A1 => n116918, A2 => n116919, A3 => n116920, A4 
                           => n116921, ZN => n5356);
   U88462 : AOI221_X1 port map( B1 => n119889, B2 => n118531, C1 => n119883, C2
                           => n118843, A => n116939, ZN => n116919);
   U88463 : AOI221_X1 port map( B1 => n119865, B2 => n95474, C1 => n119859, C2 
                           => n118430, A => n116940, ZN => n116918);
   U88464 : NOR4_X1 port map( A1 => n116934, A2 => n116935, A3 => n116936, A4 
                           => n116937, ZN => n116920);
   U88465 : NAND4_X1 port map( A1 => n116895, A2 => n116896, A3 => n116897, A4 
                           => n116898, ZN => n5357);
   U88466 : AOI221_X1 port map( B1 => n119889, B2 => n118532, C1 => n119883, C2
                           => n118844, A => n116916, ZN => n116896);
   U88467 : AOI221_X1 port map( B1 => n119865, B2 => n95475, C1 => n119859, C2 
                           => n118431, A => n116917, ZN => n116895);
   U88468 : NOR4_X1 port map( A1 => n116911, A2 => n116912, A3 => n116913, A4 
                           => n116914, ZN => n116897);
   U88469 : NAND4_X1 port map( A1 => n116872, A2 => n116873, A3 => n116874, A4 
                           => n116875, ZN => n5358);
   U88470 : AOI221_X1 port map( B1 => n119889, B2 => n118533, C1 => n119883, C2
                           => n118845, A => n116893, ZN => n116873);
   U88471 : AOI221_X1 port map( B1 => n119865, B2 => n95476, C1 => n119859, C2 
                           => n118432, A => n116894, ZN => n116872);
   U88472 : NOR4_X1 port map( A1 => n116888, A2 => n116889, A3 => n116890, A4 
                           => n116891, ZN => n116874);
   U88473 : NAND4_X1 port map( A1 => n116849, A2 => n116850, A3 => n116851, A4 
                           => n116852, ZN => n5359);
   U88474 : AOI221_X1 port map( B1 => n119890, B2 => n118534, C1 => n119884, C2
                           => n118846, A => n116870, ZN => n116850);
   U88475 : AOI221_X1 port map( B1 => n119866, B2 => n95477, C1 => n119860, C2 
                           => n118433, A => n116871, ZN => n116849);
   U88476 : NOR4_X1 port map( A1 => n116865, A2 => n116866, A3 => n116867, A4 
                           => n116868, ZN => n116851);
   U88477 : NAND4_X1 port map( A1 => n116826, A2 => n116827, A3 => n116828, A4 
                           => n116829, ZN => n5360);
   U88478 : AOI221_X1 port map( B1 => n119890, B2 => n118535, C1 => n119884, C2
                           => n118847, A => n116847, ZN => n116827);
   U88479 : AOI221_X1 port map( B1 => n119866, B2 => n95478, C1 => n119860, C2 
                           => n118434, A => n116848, ZN => n116826);
   U88480 : NOR4_X1 port map( A1 => n116842, A2 => n116843, A3 => n116844, A4 
                           => n116845, ZN => n116828);
   U88481 : NAND4_X1 port map( A1 => n116803, A2 => n116804, A3 => n116805, A4 
                           => n116806, ZN => n5361);
   U88482 : AOI221_X1 port map( B1 => n119890, B2 => n118536, C1 => n119884, C2
                           => n118848, A => n116824, ZN => n116804);
   U88483 : AOI221_X1 port map( B1 => n119866, B2 => n95479, C1 => n119860, C2 
                           => n118435, A => n116825, ZN => n116803);
   U88484 : NOR4_X1 port map( A1 => n116819, A2 => n116820, A3 => n116821, A4 
                           => n116822, ZN => n116805);
   U88485 : NAND4_X1 port map( A1 => n116780, A2 => n116781, A3 => n116782, A4 
                           => n116783, ZN => n5362);
   U88486 : AOI221_X1 port map( B1 => n119890, B2 => n118537, C1 => n119884, C2
                           => n118849, A => n116801, ZN => n116781);
   U88487 : AOI221_X1 port map( B1 => n119866, B2 => n95480, C1 => n119860, C2 
                           => n118436, A => n116802, ZN => n116780);
   U88488 : NOR4_X1 port map( A1 => n116796, A2 => n116797, A3 => n116798, A4 
                           => n116799, ZN => n116782);
   U88489 : NAND4_X1 port map( A1 => n116757, A2 => n116758, A3 => n116759, A4 
                           => n116760, ZN => n5363);
   U88490 : AOI221_X1 port map( B1 => n119890, B2 => n118538, C1 => n119884, C2
                           => n118850, A => n116778, ZN => n116758);
   U88491 : AOI221_X1 port map( B1 => n119866, B2 => n95481, C1 => n119860, C2 
                           => n118437, A => n116779, ZN => n116757);
   U88492 : NOR4_X1 port map( A1 => n116773, A2 => n116774, A3 => n116775, A4 
                           => n116776, ZN => n116759);
   U88493 : NAND4_X1 port map( A1 => n116734, A2 => n116735, A3 => n116736, A4 
                           => n116737, ZN => n5364);
   U88494 : AOI221_X1 port map( B1 => n119890, B2 => n118539, C1 => n119884, C2
                           => n118851, A => n116755, ZN => n116735);
   U88495 : AOI221_X1 port map( B1 => n119866, B2 => n95482, C1 => n119860, C2 
                           => n118438, A => n116756, ZN => n116734);
   U88496 : NOR4_X1 port map( A1 => n116750, A2 => n116751, A3 => n116752, A4 
                           => n116753, ZN => n116736);
   U88497 : NAND4_X1 port map( A1 => n116711, A2 => n116712, A3 => n116713, A4 
                           => n116714, ZN => n5365);
   U88498 : AOI221_X1 port map( B1 => n119890, B2 => n118540, C1 => n119884, C2
                           => n118852, A => n116732, ZN => n116712);
   U88499 : AOI221_X1 port map( B1 => n119866, B2 => n95483, C1 => n119860, C2 
                           => n118439, A => n116733, ZN => n116711);
   U88500 : NOR4_X1 port map( A1 => n116727, A2 => n116728, A3 => n116729, A4 
                           => n116730, ZN => n116713);
   U88501 : NAND4_X1 port map( A1 => n116688, A2 => n116689, A3 => n116690, A4 
                           => n116691, ZN => n5366);
   U88502 : AOI221_X1 port map( B1 => n119890, B2 => n118541, C1 => n119884, C2
                           => n118853, A => n116709, ZN => n116689);
   U88503 : AOI221_X1 port map( B1 => n119866, B2 => n95484, C1 => n119860, C2 
                           => n118440, A => n116710, ZN => n116688);
   U88504 : NOR4_X1 port map( A1 => n116704, A2 => n116705, A3 => n116706, A4 
                           => n116707, ZN => n116690);
   U88505 : NAND4_X1 port map( A1 => n116665, A2 => n116666, A3 => n116667, A4 
                           => n116668, ZN => n5367);
   U88506 : AOI221_X1 port map( B1 => n119890, B2 => n118542, C1 => n119884, C2
                           => n118854, A => n116686, ZN => n116666);
   U88507 : AOI221_X1 port map( B1 => n119866, B2 => n95485, C1 => n119860, C2 
                           => n118441, A => n116687, ZN => n116665);
   U88508 : NOR4_X1 port map( A1 => n116681, A2 => n116682, A3 => n116683, A4 
                           => n116684, ZN => n116667);
   U88509 : NAND4_X1 port map( A1 => n116642, A2 => n116643, A3 => n116644, A4 
                           => n116645, ZN => n5368);
   U88510 : AOI221_X1 port map( B1 => n119890, B2 => n118543, C1 => n119884, C2
                           => n118855, A => n116663, ZN => n116643);
   U88511 : AOI221_X1 port map( B1 => n119866, B2 => n95486, C1 => n119860, C2 
                           => n118442, A => n116664, ZN => n116642);
   U88512 : NOR4_X1 port map( A1 => n116658, A2 => n116659, A3 => n116660, A4 
                           => n116661, ZN => n116644);
   U88513 : NAND4_X1 port map( A1 => n116619, A2 => n116620, A3 => n116621, A4 
                           => n116622, ZN => n5369);
   U88514 : AOI221_X1 port map( B1 => n119890, B2 => n118544, C1 => n119884, C2
                           => n118856, A => n116640, ZN => n116620);
   U88515 : AOI221_X1 port map( B1 => n119866, B2 => n95487, C1 => n119860, C2 
                           => n118443, A => n116641, ZN => n116619);
   U88516 : NOR4_X1 port map( A1 => n116635, A2 => n116636, A3 => n116637, A4 
                           => n116638, ZN => n116621);
   U88517 : NAND4_X1 port map( A1 => n116596, A2 => n116597, A3 => n116598, A4 
                           => n116599, ZN => n5370);
   U88518 : AOI221_X1 port map( B1 => n119890, B2 => n118545, C1 => n119884, C2
                           => n118857, A => n116617, ZN => n116597);
   U88519 : AOI221_X1 port map( B1 => n119866, B2 => n95488, C1 => n119860, C2 
                           => n118444, A => n116618, ZN => n116596);
   U88520 : NOR4_X1 port map( A1 => n116612, A2 => n116613, A3 => n116614, A4 
                           => n116615, ZN => n116598);
   U88521 : NAND4_X1 port map( A1 => n114757, A2 => n114758, A3 => n114759, A4 
                           => n114760, ZN => n5495);
   U88522 : AOI221_X1 port map( B1 => n120065, B2 => n119174, C1 => n120059, C2
                           => n117985, A => n114781, ZN => n114757);
   U88523 : NOR4_X1 port map( A1 => n114761, A2 => n114762, A3 => n114763, A4 
                           => n114764, ZN => n114760);
   U88524 : NOR4_X1 port map( A1 => n114773, A2 => n114774, A3 => n114775, A4 
                           => n114776, ZN => n114759);
   U88525 : NAND4_X1 port map( A1 => n114731, A2 => n114732, A3 => n114733, A4 
                           => n114734, ZN => n5497);
   U88526 : AOI221_X1 port map( B1 => n120065, B2 => n119175, C1 => n120059, C2
                           => n117986, A => n114755, ZN => n114731);
   U88527 : NOR4_X1 port map( A1 => n114735, A2 => n114736, A3 => n114737, A4 
                           => n114738, ZN => n114734);
   U88528 : NOR4_X1 port map( A1 => n114747, A2 => n114748, A3 => n114749, A4 
                           => n114750, ZN => n114733);
   U88529 : NAND4_X1 port map( A1 => n114705, A2 => n114706, A3 => n114707, A4 
                           => n114708, ZN => n5499);
   U88530 : AOI221_X1 port map( B1 => n120065, B2 => n119176, C1 => n120059, C2
                           => n117987, A => n114729, ZN => n114705);
   U88531 : NOR4_X1 port map( A1 => n114709, A2 => n114710, A3 => n114711, A4 
                           => n114712, ZN => n114708);
   U88532 : NOR4_X1 port map( A1 => n114721, A2 => n114722, A3 => n114723, A4 
                           => n114724, ZN => n114707);
   U88533 : NAND4_X1 port map( A1 => n114646, A2 => n114647, A3 => n114648, A4 
                           => n114649, ZN => n5501);
   U88534 : AOI221_X1 port map( B1 => n120065, B2 => n119177, C1 => n120059, C2
                           => n117988, A => n114701, ZN => n114646);
   U88535 : NOR4_X1 port map( A1 => n114650, A2 => n114651, A3 => n114652, A4 
                           => n114653, ZN => n114649);
   U88536 : NOR4_X1 port map( A1 => n114678, A2 => n114679, A3 => n114680, A4 
                           => n114681, ZN => n114648);
   U88537 : NAND4_X1 port map( A1 => n116575, A2 => n116576, A3 => n116577, A4 
                           => n116578, ZN => n5371);
   U88538 : NOR4_X1 port map( A1 => n116589, A2 => n116590, A3 => n116591, A4 
                           => n116592, ZN => n116577);
   U88539 : AOI221_X1 port map( B1 => n119891, B2 => n109895, C1 => n119885, C2
                           => n118858, A => n116594, ZN => n116576);
   U88540 : NOR4_X1 port map( A1 => n116579, A2 => n116580, A3 => n116581, A4 
                           => n116582, ZN => n116578);
   U88541 : NAND4_X1 port map( A1 => n116554, A2 => n116555, A3 => n116556, A4 
                           => n116557, ZN => n5372);
   U88542 : NOR4_X1 port map( A1 => n116568, A2 => n116569, A3 => n116570, A4 
                           => n116571, ZN => n116556);
   U88543 : AOI221_X1 port map( B1 => n119891, B2 => n109896, C1 => n119885, C2
                           => n118859, A => n116573, ZN => n116555);
   U88544 : NOR4_X1 port map( A1 => n116558, A2 => n116559, A3 => n116560, A4 
                           => n116561, ZN => n116557);
   U88545 : NAND4_X1 port map( A1 => n116533, A2 => n116534, A3 => n116535, A4 
                           => n116536, ZN => n5373);
   U88546 : NOR4_X1 port map( A1 => n116547, A2 => n116548, A3 => n116549, A4 
                           => n116550, ZN => n116535);
   U88547 : AOI221_X1 port map( B1 => n119891, B2 => n109897, C1 => n119885, C2
                           => n118860, A => n116552, ZN => n116534);
   U88548 : NOR4_X1 port map( A1 => n116537, A2 => n116538, A3 => n116539, A4 
                           => n116540, ZN => n116536);
   U88549 : NAND4_X1 port map( A1 => n116479, A2 => n116480, A3 => n116481, A4 
                           => n116482, ZN => n5374);
   U88550 : NOR4_X1 port map( A1 => n116509, A2 => n116510, A3 => n116511, A4 
                           => n116512, ZN => n116481);
   U88551 : AOI221_X1 port map( B1 => n119891, B2 => n109898, C1 => n119885, C2
                           => n118861, A => n116525, ZN => n116480);
   U88552 : NOR4_X1 port map( A1 => n116483, A2 => n116484, A3 => n116485, A4 
                           => n116486, ZN => n116482);
   U88553 : NAND4_X1 port map( A1 => n115147, A2 => n115148, A3 => n115149, A4 
                           => n115150, ZN => n5467);
   U88554 : AOI221_X1 port map( B1 => n120063, B2 => n119178, C1 => n120057, C2
                           => n118431, A => n115173, ZN => n115147);
   U88555 : AOI221_X1 port map( B1 => n120087, B2 => n118986, C1 => n120081, C2
                           => n118550, A => n115171, ZN => n115148);
   U88556 : NOR4_X1 port map( A1 => n115165, A2 => n115166, A3 => n115167, A4 
                           => n115168, ZN => n115149);
   U88557 : NAND4_X1 port map( A1 => n115119, A2 => n115120, A3 => n115121, A4 
                           => n115122, ZN => n5469);
   U88558 : AOI221_X1 port map( B1 => n120063, B2 => n119179, C1 => n120057, C2
                           => n118432, A => n115145, ZN => n115119);
   U88559 : AOI221_X1 port map( B1 => n120087, B2 => n118987, C1 => n120081, C2
                           => n118551, A => n115143, ZN => n115120);
   U88560 : NOR4_X1 port map( A1 => n115137, A2 => n115138, A3 => n115139, A4 
                           => n115140, ZN => n115121);
   U88561 : NAND4_X1 port map( A1 => n115091, A2 => n115092, A3 => n115093, A4 
                           => n115094, ZN => n5471);
   U88562 : AOI221_X1 port map( B1 => n120064, B2 => n119180, C1 => n120058, C2
                           => n118433, A => n115117, ZN => n115091);
   U88563 : AOI221_X1 port map( B1 => n120088, B2 => n118988, C1 => n120082, C2
                           => n118552, A => n115115, ZN => n115092);
   U88564 : NOR4_X1 port map( A1 => n115109, A2 => n115110, A3 => n115111, A4 
                           => n115112, ZN => n115093);
   U88565 : NAND4_X1 port map( A1 => n115063, A2 => n115064, A3 => n115065, A4 
                           => n115066, ZN => n5473);
   U88566 : AOI221_X1 port map( B1 => n120064, B2 => n119181, C1 => n120058, C2
                           => n118434, A => n115089, ZN => n115063);
   U88567 : AOI221_X1 port map( B1 => n120088, B2 => n118989, C1 => n120082, C2
                           => n118553, A => n115087, ZN => n115064);
   U88568 : NOR4_X1 port map( A1 => n115081, A2 => n115082, A3 => n115083, A4 
                           => n115084, ZN => n115065);
   U88569 : NAND4_X1 port map( A1 => n115035, A2 => n115036, A3 => n115037, A4 
                           => n115038, ZN => n5475);
   U88570 : AOI221_X1 port map( B1 => n120064, B2 => n119182, C1 => n120058, C2
                           => n118435, A => n115061, ZN => n115035);
   U88571 : AOI221_X1 port map( B1 => n120088, B2 => n118990, C1 => n120082, C2
                           => n118554, A => n115059, ZN => n115036);
   U88572 : NOR4_X1 port map( A1 => n115053, A2 => n115054, A3 => n115055, A4 
                           => n115056, ZN => n115037);
   U88573 : NAND4_X1 port map( A1 => n115007, A2 => n115008, A3 => n115009, A4 
                           => n115010, ZN => n5477);
   U88574 : AOI221_X1 port map( B1 => n120064, B2 => n119183, C1 => n120058, C2
                           => n118436, A => n115033, ZN => n115007);
   U88575 : AOI221_X1 port map( B1 => n120088, B2 => n118991, C1 => n120082, C2
                           => n118555, A => n115031, ZN => n115008);
   U88576 : NOR4_X1 port map( A1 => n115025, A2 => n115026, A3 => n115027, A4 
                           => n115028, ZN => n115009);
   U88577 : NAND4_X1 port map( A1 => n114979, A2 => n114980, A3 => n114981, A4 
                           => n114982, ZN => n5479);
   U88578 : AOI221_X1 port map( B1 => n120064, B2 => n119184, C1 => n120058, C2
                           => n118437, A => n115005, ZN => n114979);
   U88579 : AOI221_X1 port map( B1 => n120088, B2 => n118992, C1 => n120082, C2
                           => n118556, A => n115003, ZN => n114980);
   U88580 : NOR4_X1 port map( A1 => n114997, A2 => n114998, A3 => n114999, A4 
                           => n115000, ZN => n114981);
   U88581 : NAND4_X1 port map( A1 => n114951, A2 => n114952, A3 => n114953, A4 
                           => n114954, ZN => n5481);
   U88582 : AOI221_X1 port map( B1 => n120064, B2 => n119185, C1 => n120058, C2
                           => n118438, A => n114977, ZN => n114951);
   U88583 : AOI221_X1 port map( B1 => n120088, B2 => n118993, C1 => n120082, C2
                           => n118557, A => n114975, ZN => n114952);
   U88584 : NOR4_X1 port map( A1 => n114969, A2 => n114970, A3 => n114971, A4 
                           => n114972, ZN => n114953);
   U88585 : NAND4_X1 port map( A1 => n114923, A2 => n114924, A3 => n114925, A4 
                           => n114926, ZN => n5483);
   U88586 : AOI221_X1 port map( B1 => n120064, B2 => n119186, C1 => n120058, C2
                           => n118439, A => n114949, ZN => n114923);
   U88587 : AOI221_X1 port map( B1 => n120088, B2 => n118994, C1 => n120082, C2
                           => n118558, A => n114947, ZN => n114924);
   U88588 : NOR4_X1 port map( A1 => n114941, A2 => n114942, A3 => n114943, A4 
                           => n114944, ZN => n114925);
   U88589 : NAND4_X1 port map( A1 => n114895, A2 => n114896, A3 => n114897, A4 
                           => n114898, ZN => n5485);
   U88590 : AOI221_X1 port map( B1 => n120064, B2 => n119187, C1 => n120058, C2
                           => n118440, A => n114921, ZN => n114895);
   U88591 : AOI221_X1 port map( B1 => n120088, B2 => n118995, C1 => n120082, C2
                           => n118559, A => n114919, ZN => n114896);
   U88592 : NOR4_X1 port map( A1 => n114913, A2 => n114914, A3 => n114915, A4 
                           => n114916, ZN => n114897);
   U88593 : NAND4_X1 port map( A1 => n114867, A2 => n114868, A3 => n114869, A4 
                           => n114870, ZN => n5487);
   U88594 : AOI221_X1 port map( B1 => n120064, B2 => n119188, C1 => n120058, C2
                           => n118441, A => n114893, ZN => n114867);
   U88595 : AOI221_X1 port map( B1 => n120088, B2 => n118996, C1 => n120082, C2
                           => n118560, A => n114891, ZN => n114868);
   U88596 : NOR4_X1 port map( A1 => n114885, A2 => n114886, A3 => n114887, A4 
                           => n114888, ZN => n114869);
   U88597 : NAND4_X1 port map( A1 => n114839, A2 => n114840, A3 => n114841, A4 
                           => n114842, ZN => n5489);
   U88598 : AOI221_X1 port map( B1 => n120064, B2 => n119189, C1 => n120058, C2
                           => n118442, A => n114865, ZN => n114839);
   U88599 : AOI221_X1 port map( B1 => n120088, B2 => n118997, C1 => n120082, C2
                           => n118561, A => n114863, ZN => n114840);
   U88600 : NOR4_X1 port map( A1 => n114857, A2 => n114858, A3 => n114859, A4 
                           => n114860, ZN => n114841);
   U88601 : NAND4_X1 port map( A1 => n114811, A2 => n114812, A3 => n114813, A4 
                           => n114814, ZN => n5491);
   U88602 : AOI221_X1 port map( B1 => n120064, B2 => n119190, C1 => n120058, C2
                           => n118443, A => n114837, ZN => n114811);
   U88603 : AOI221_X1 port map( B1 => n120088, B2 => n118998, C1 => n120082, C2
                           => n118562, A => n114835, ZN => n114812);
   U88604 : NOR4_X1 port map( A1 => n114829, A2 => n114830, A3 => n114831, A4 
                           => n114832, ZN => n114813);
   U88605 : NAND4_X1 port map( A1 => n114783, A2 => n114784, A3 => n114785, A4 
                           => n114786, ZN => n5493);
   U88606 : AOI221_X1 port map( B1 => n120064, B2 => n119191, C1 => n120058, C2
                           => n118444, A => n114809, ZN => n114783);
   U88607 : AOI221_X1 port map( B1 => n120088, B2 => n118999, C1 => n120082, C2
                           => n118563, A => n114807, ZN => n114784);
   U88608 : NOR4_X1 port map( A1 => n114801, A2 => n114802, A3 => n114803, A4 
                           => n114804, ZN => n114785);
   U88609 : NAND4_X1 port map( A1 => n116435, A2 => n116436, A3 => n116437, A4 
                           => n116438, ZN => n5375);
   U88610 : AOI221_X1 port map( B1 => n120060, B2 => n119192, C1 => n120054, C2
                           => n118385, A => n116477, ZN => n116435);
   U88611 : AOI221_X1 port map( B1 => n120084, B2 => n119000, C1 => n120078, C2
                           => n118564, A => n116474, ZN => n116436);
   U88612 : NOR4_X1 port map( A1 => n116465, A2 => n116466, A3 => n116467, A4 
                           => n116468, ZN => n116437);
   U88613 : NAND4_X1 port map( A1 => n116407, A2 => n116408, A3 => n116409, A4 
                           => n116410, ZN => n5377);
   U88614 : AOI221_X1 port map( B1 => n120060, B2 => n119193, C1 => n120054, C2
                           => n118386, A => n116433, ZN => n116407);
   U88615 : AOI221_X1 port map( B1 => n120084, B2 => n119001, C1 => n120078, C2
                           => n118565, A => n116431, ZN => n116408);
   U88616 : NOR4_X1 port map( A1 => n116425, A2 => n116426, A3 => n116427, A4 
                           => n116428, ZN => n116409);
   U88617 : NAND4_X1 port map( A1 => n116379, A2 => n116380, A3 => n116381, A4 
                           => n116382, ZN => n5379);
   U88618 : AOI221_X1 port map( B1 => n120060, B2 => n119194, C1 => n120054, C2
                           => n118387, A => n116405, ZN => n116379);
   U88619 : AOI221_X1 port map( B1 => n120084, B2 => n119002, C1 => n120078, C2
                           => n118566, A => n116403, ZN => n116380);
   U88620 : NOR4_X1 port map( A1 => n116397, A2 => n116398, A3 => n116399, A4 
                           => n116400, ZN => n116381);
   U88621 : NAND4_X1 port map( A1 => n116351, A2 => n116352, A3 => n116353, A4 
                           => n116354, ZN => n5381);
   U88622 : AOI221_X1 port map( B1 => n120060, B2 => n119195, C1 => n120054, C2
                           => n118388, A => n116377, ZN => n116351);
   U88623 : AOI221_X1 port map( B1 => n120084, B2 => n119003, C1 => n120078, C2
                           => n118567, A => n116375, ZN => n116352);
   U88624 : NOR4_X1 port map( A1 => n116369, A2 => n116370, A3 => n116371, A4 
                           => n116372, ZN => n116353);
   U88625 : NAND4_X1 port map( A1 => n117781, A2 => n117782, A3 => n117783, A4 
                           => n117784, ZN => n5318);
   U88626 : AOI221_X1 port map( B1 => n119886, B2 => n118806, C1 => n119880, C2
                           => n109986, A => n117801, ZN => n117782);
   U88627 : AOI221_X1 port map( B1 => n119862, B2 => n95436, C1 => n119856, C2 
                           => n118392, A => n117802, ZN => n117781);
   U88628 : NOR4_X1 port map( A1 => n117797, A2 => n117798, A3 => n117799, A4 
                           => n117800, ZN => n117783);
   U88629 : NAND4_X1 port map( A1 => n117759, A2 => n117760, A3 => n117761, A4 
                           => n117762, ZN => n5319);
   U88630 : AOI221_X1 port map( B1 => n119886, B2 => n118807, C1 => n119880, C2
                           => n109987, A => n117779, ZN => n117760);
   U88631 : AOI221_X1 port map( B1 => n119862, B2 => n95437, C1 => n119856, C2 
                           => n118393, A => n117780, ZN => n117759);
   U88632 : NOR4_X1 port map( A1 => n117775, A2 => n117776, A3 => n117777, A4 
                           => n117778, ZN => n117761);
   U88633 : NAND4_X1 port map( A1 => n117737, A2 => n117738, A3 => n117739, A4 
                           => n117740, ZN => n5320);
   U88634 : AOI221_X1 port map( B1 => n119886, B2 => n118808, C1 => n119880, C2
                           => n109988, A => n117757, ZN => n117738);
   U88635 : AOI221_X1 port map( B1 => n119862, B2 => n95438, C1 => n119856, C2 
                           => n118394, A => n117758, ZN => n117737);
   U88636 : NOR4_X1 port map( A1 => n117753, A2 => n117754, A3 => n117755, A4 
                           => n117756, ZN => n117739);
   U88637 : NAND4_X1 port map( A1 => n117715, A2 => n117716, A3 => n117717, A4 
                           => n117718, ZN => n5321);
   U88638 : AOI221_X1 port map( B1 => n119886, B2 => n118809, C1 => n119880, C2
                           => n109989, A => n117735, ZN => n117716);
   U88639 : AOI221_X1 port map( B1 => n119862, B2 => n95439, C1 => n119856, C2 
                           => n118395, A => n117736, ZN => n117715);
   U88640 : NOR4_X1 port map( A1 => n117731, A2 => n117732, A3 => n117733, A4 
                           => n117734, ZN => n117717);
   U88641 : NAND4_X1 port map( A1 => n117935, A2 => n117936, A3 => n117937, A4 
                           => n117938, ZN => n5311);
   U88642 : AOI221_X1 port map( B1 => n119886, B2 => n118810, C1 => n119880, C2
                           => n109979, A => n117969, ZN => n117936);
   U88643 : AOI221_X1 port map( B1 => n119862, B2 => n95429, C1 => n119856, C2 
                           => n118385, A => n117972, ZN => n117935);
   U88644 : NOR4_X1 port map( A1 => n117963, A2 => n117964, A3 => n117965, A4 
                           => n117966, ZN => n117937);
   U88645 : NAND4_X1 port map( A1 => n117913, A2 => n117914, A3 => n117915, A4 
                           => n117916, ZN => n5312);
   U88646 : AOI221_X1 port map( B1 => n119886, B2 => n118811, C1 => n119880, C2
                           => n109980, A => n117933, ZN => n117914);
   U88647 : AOI221_X1 port map( B1 => n119862, B2 => n95430, C1 => n119856, C2 
                           => n118386, A => n117934, ZN => n117913);
   U88648 : NOR4_X1 port map( A1 => n117929, A2 => n117930, A3 => n117931, A4 
                           => n117932, ZN => n117915);
   U88649 : NAND4_X1 port map( A1 => n117891, A2 => n117892, A3 => n117893, A4 
                           => n117894, ZN => n5313);
   U88650 : AOI221_X1 port map( B1 => n119886, B2 => n118812, C1 => n119880, C2
                           => n109981, A => n117911, ZN => n117892);
   U88651 : AOI221_X1 port map( B1 => n119862, B2 => n95431, C1 => n119856, C2 
                           => n118387, A => n117912, ZN => n117891);
   U88652 : NOR4_X1 port map( A1 => n117907, A2 => n117908, A3 => n117909, A4 
                           => n117910, ZN => n117893);
   U88653 : NAND4_X1 port map( A1 => n117869, A2 => n117870, A3 => n117871, A4 
                           => n117872, ZN => n5314);
   U88654 : AOI221_X1 port map( B1 => n119886, B2 => n118813, C1 => n119880, C2
                           => n109982, A => n117889, ZN => n117870);
   U88655 : AOI221_X1 port map( B1 => n119862, B2 => n95432, C1 => n119856, C2 
                           => n118388, A => n117890, ZN => n117869);
   U88656 : NOR4_X1 port map( A1 => n117885, A2 => n117886, A3 => n117887, A4 
                           => n117888, ZN => n117871);
   U88657 : NAND4_X1 port map( A1 => n117847, A2 => n117848, A3 => n117849, A4 
                           => n117850, ZN => n5315);
   U88658 : AOI221_X1 port map( B1 => n119886, B2 => n118814, C1 => n119880, C2
                           => n109983, A => n117867, ZN => n117848);
   U88659 : AOI221_X1 port map( B1 => n119862, B2 => n95433, C1 => n119856, C2 
                           => n118389, A => n117868, ZN => n117847);
   U88660 : NOR4_X1 port map( A1 => n117863, A2 => n117864, A3 => n117865, A4 
                           => n117866, ZN => n117849);
   U88661 : NAND4_X1 port map( A1 => n117825, A2 => n117826, A3 => n117827, A4 
                           => n117828, ZN => n5316);
   U88662 : AOI221_X1 port map( B1 => n119886, B2 => n118815, C1 => n119880, C2
                           => n109984, A => n117845, ZN => n117826);
   U88663 : AOI221_X1 port map( B1 => n119862, B2 => n95434, C1 => n119856, C2 
                           => n118390, A => n117846, ZN => n117825);
   U88664 : NOR4_X1 port map( A1 => n117841, A2 => n117842, A3 => n117843, A4 
                           => n117844, ZN => n117827);
   U88665 : NAND4_X1 port map( A1 => n117803, A2 => n117804, A3 => n117805, A4 
                           => n117806, ZN => n5317);
   U88666 : AOI221_X1 port map( B1 => n119886, B2 => n118816, C1 => n119880, C2
                           => n109985, A => n117823, ZN => n117804);
   U88667 : AOI221_X1 port map( B1 => n119862, B2 => n95435, C1 => n119856, C2 
                           => n118391, A => n117824, ZN => n117803);
   U88668 : NOR4_X1 port map( A1 => n117819, A2 => n117820, A3 => n117821, A4 
                           => n117822, ZN => n117805);
   U88669 : NAND4_X1 port map( A1 => n116323, A2 => n116324, A3 => n116325, A4 
                           => n116326, ZN => n5383);
   U88670 : AOI221_X1 port map( B1 => n120060, B2 => n119196, C1 => n120054, C2
                           => n118389, A => n116349, ZN => n116323);
   U88671 : AOI221_X1 port map( B1 => n120084, B2 => n119004, C1 => n120078, C2
                           => n118568, A => n116347, ZN => n116324);
   U88672 : NOR4_X1 port map( A1 => n116341, A2 => n116342, A3 => n116343, A4 
                           => n116344, ZN => n116325);
   U88673 : NAND4_X1 port map( A1 => n116295, A2 => n116296, A3 => n116297, A4 
                           => n116298, ZN => n5385);
   U88674 : AOI221_X1 port map( B1 => n120060, B2 => n119197, C1 => n120054, C2
                           => n118390, A => n116321, ZN => n116295);
   U88675 : AOI221_X1 port map( B1 => n120084, B2 => n119005, C1 => n120078, C2
                           => n118569, A => n116319, ZN => n116296);
   U88676 : NOR4_X1 port map( A1 => n116313, A2 => n116314, A3 => n116315, A4 
                           => n116316, ZN => n116297);
   U88677 : NAND4_X1 port map( A1 => n116267, A2 => n116268, A3 => n116269, A4 
                           => n116270, ZN => n5387);
   U88678 : AOI221_X1 port map( B1 => n120060, B2 => n119198, C1 => n120054, C2
                           => n118391, A => n116293, ZN => n116267);
   U88679 : AOI221_X1 port map( B1 => n120084, B2 => n119006, C1 => n120078, C2
                           => n118570, A => n116291, ZN => n116268);
   U88680 : NOR4_X1 port map( A1 => n116285, A2 => n116286, A3 => n116287, A4 
                           => n116288, ZN => n116269);
   U88681 : NAND4_X1 port map( A1 => n116239, A2 => n116240, A3 => n116241, A4 
                           => n116242, ZN => n5389);
   U88682 : AOI221_X1 port map( B1 => n120060, B2 => n119199, C1 => n120054, C2
                           => n118392, A => n116265, ZN => n116239);
   U88683 : AOI221_X1 port map( B1 => n120084, B2 => n119007, C1 => n120078, C2
                           => n118571, A => n116263, ZN => n116240);
   U88684 : NOR4_X1 port map( A1 => n116257, A2 => n116258, A3 => n116259, A4 
                           => n116260, ZN => n116241);
   U88685 : NAND4_X1 port map( A1 => n116211, A2 => n116212, A3 => n116213, A4 
                           => n116214, ZN => n5391);
   U88686 : AOI221_X1 port map( B1 => n120060, B2 => n119200, C1 => n120054, C2
                           => n118393, A => n116237, ZN => n116211);
   U88687 : AOI221_X1 port map( B1 => n120084, B2 => n119008, C1 => n120078, C2
                           => n118572, A => n116235, ZN => n116212);
   U88688 : NOR4_X1 port map( A1 => n116229, A2 => n116230, A3 => n116231, A4 
                           => n116232, ZN => n116213);
   U88689 : NAND4_X1 port map( A1 => n116183, A2 => n116184, A3 => n116185, A4 
                           => n116186, ZN => n5393);
   U88690 : AOI221_X1 port map( B1 => n120060, B2 => n119201, C1 => n120054, C2
                           => n118394, A => n116209, ZN => n116183);
   U88691 : AOI221_X1 port map( B1 => n120084, B2 => n119009, C1 => n120078, C2
                           => n118573, A => n116207, ZN => n116184);
   U88692 : NOR4_X1 port map( A1 => n116201, A2 => n116202, A3 => n116203, A4 
                           => n116204, ZN => n116185);
   U88693 : NAND4_X1 port map( A1 => n116155, A2 => n116156, A3 => n116157, A4 
                           => n116158, ZN => n5395);
   U88694 : AOI221_X1 port map( B1 => n120060, B2 => n119202, C1 => n120054, C2
                           => n118395, A => n116181, ZN => n116155);
   U88695 : AOI221_X1 port map( B1 => n120084, B2 => n119010, C1 => n120078, C2
                           => n118574, A => n116179, ZN => n116156);
   U88696 : NOR4_X1 port map( A1 => n116173, A2 => n116174, A3 => n116175, A4 
                           => n116176, ZN => n116157);
   U88697 : NAND4_X1 port map( A1 => n116127, A2 => n116128, A3 => n116129, A4 
                           => n116130, ZN => n5397);
   U88698 : AOI221_X1 port map( B1 => n120060, B2 => n119203, C1 => n120054, C2
                           => n118396, A => n116153, ZN => n116127);
   U88699 : AOI221_X1 port map( B1 => n120084, B2 => n119011, C1 => n120078, C2
                           => n118575, A => n116151, ZN => n116128);
   U88700 : NOR4_X1 port map( A1 => n116145, A2 => n116146, A3 => n116147, A4 
                           => n116148, ZN => n116129);
   U88701 : NAND4_X1 port map( A1 => n116099, A2 => n116100, A3 => n116101, A4 
                           => n116102, ZN => n5399);
   U88702 : AOI221_X1 port map( B1 => n120061, B2 => n119204, C1 => n120055, C2
                           => n118397, A => n116125, ZN => n116099);
   U88703 : AOI221_X1 port map( B1 => n120085, B2 => n119012, C1 => n120079, C2
                           => n118576, A => n116123, ZN => n116100);
   U88704 : NOR4_X1 port map( A1 => n116117, A2 => n116118, A3 => n116119, A4 
                           => n116120, ZN => n116101);
   U88705 : NAND4_X1 port map( A1 => n116071, A2 => n116072, A3 => n116073, A4 
                           => n116074, ZN => n5401);
   U88706 : AOI221_X1 port map( B1 => n120061, B2 => n119205, C1 => n120055, C2
                           => n118398, A => n116097, ZN => n116071);
   U88707 : AOI221_X1 port map( B1 => n120085, B2 => n119013, C1 => n120079, C2
                           => n118577, A => n116095, ZN => n116072);
   U88708 : NOR4_X1 port map( A1 => n116089, A2 => n116090, A3 => n116091, A4 
                           => n116092, ZN => n116073);
   U88709 : NAND4_X1 port map( A1 => n116043, A2 => n116044, A3 => n116045, A4 
                           => n116046, ZN => n5403);
   U88710 : AOI221_X1 port map( B1 => n120061, B2 => n119206, C1 => n120055, C2
                           => n118399, A => n116069, ZN => n116043);
   U88711 : AOI221_X1 port map( B1 => n120085, B2 => n119014, C1 => n120079, C2
                           => n118578, A => n116067, ZN => n116044);
   U88712 : NOR4_X1 port map( A1 => n116061, A2 => n116062, A3 => n116063, A4 
                           => n116064, ZN => n116045);
   U88713 : NAND4_X1 port map( A1 => n116015, A2 => n116016, A3 => n116017, A4 
                           => n116018, ZN => n5405);
   U88714 : AOI221_X1 port map( B1 => n120061, B2 => n119207, C1 => n120055, C2
                           => n118400, A => n116041, ZN => n116015);
   U88715 : AOI221_X1 port map( B1 => n120085, B2 => n119015, C1 => n120079, C2
                           => n118579, A => n116039, ZN => n116016);
   U88716 : NOR4_X1 port map( A1 => n116033, A2 => n116034, A3 => n116035, A4 
                           => n116036, ZN => n116017);
   U88717 : NAND4_X1 port map( A1 => n115987, A2 => n115988, A3 => n115989, A4 
                           => n115990, ZN => n5407);
   U88718 : AOI221_X1 port map( B1 => n120061, B2 => n119208, C1 => n120055, C2
                           => n118401, A => n116013, ZN => n115987);
   U88719 : AOI221_X1 port map( B1 => n120085, B2 => n119016, C1 => n120079, C2
                           => n118580, A => n116011, ZN => n115988);
   U88720 : NOR4_X1 port map( A1 => n116005, A2 => n116006, A3 => n116007, A4 
                           => n116008, ZN => n115989);
   U88721 : NAND4_X1 port map( A1 => n115959, A2 => n115960, A3 => n115961, A4 
                           => n115962, ZN => n5409);
   U88722 : AOI221_X1 port map( B1 => n120061, B2 => n119209, C1 => n120055, C2
                           => n118402, A => n115985, ZN => n115959);
   U88723 : AOI221_X1 port map( B1 => n120085, B2 => n119017, C1 => n120079, C2
                           => n118581, A => n115983, ZN => n115960);
   U88724 : NOR4_X1 port map( A1 => n115977, A2 => n115978, A3 => n115979, A4 
                           => n115980, ZN => n115961);
   U88725 : NAND4_X1 port map( A1 => n115931, A2 => n115932, A3 => n115933, A4 
                           => n115934, ZN => n5411);
   U88726 : AOI221_X1 port map( B1 => n120061, B2 => n119210, C1 => n120055, C2
                           => n118403, A => n115957, ZN => n115931);
   U88727 : AOI221_X1 port map( B1 => n120085, B2 => n119018, C1 => n120079, C2
                           => n118582, A => n115955, ZN => n115932);
   U88728 : NOR4_X1 port map( A1 => n115949, A2 => n115950, A3 => n115951, A4 
                           => n115952, ZN => n115933);
   U88729 : NAND4_X1 port map( A1 => n115903, A2 => n115904, A3 => n115905, A4 
                           => n115906, ZN => n5413);
   U88730 : AOI221_X1 port map( B1 => n120061, B2 => n119211, C1 => n120055, C2
                           => n118404, A => n115929, ZN => n115903);
   U88731 : AOI221_X1 port map( B1 => n120085, B2 => n119019, C1 => n120079, C2
                           => n118583, A => n115927, ZN => n115904);
   U88732 : NOR4_X1 port map( A1 => n115921, A2 => n115922, A3 => n115923, A4 
                           => n115924, ZN => n115905);
   U88733 : NAND4_X1 port map( A1 => n115875, A2 => n115876, A3 => n115877, A4 
                           => n115878, ZN => n5415);
   U88734 : AOI221_X1 port map( B1 => n120061, B2 => n119212, C1 => n120055, C2
                           => n118405, A => n115901, ZN => n115875);
   U88735 : AOI221_X1 port map( B1 => n120085, B2 => n119020, C1 => n120079, C2
                           => n118584, A => n115899, ZN => n115876);
   U88736 : NOR4_X1 port map( A1 => n115893, A2 => n115894, A3 => n115895, A4 
                           => n115896, ZN => n115877);
   U88737 : NAND4_X1 port map( A1 => n115847, A2 => n115848, A3 => n115849, A4 
                           => n115850, ZN => n5417);
   U88738 : AOI221_X1 port map( B1 => n120061, B2 => n119213, C1 => n120055, C2
                           => n118406, A => n115873, ZN => n115847);
   U88739 : AOI221_X1 port map( B1 => n120085, B2 => n119021, C1 => n120079, C2
                           => n118585, A => n115871, ZN => n115848);
   U88740 : NOR4_X1 port map( A1 => n115865, A2 => n115866, A3 => n115867, A4 
                           => n115868, ZN => n115849);
   U88741 : NAND4_X1 port map( A1 => n115819, A2 => n115820, A3 => n115821, A4 
                           => n115822, ZN => n5419);
   U88742 : AOI221_X1 port map( B1 => n120061, B2 => n119214, C1 => n120055, C2
                           => n118407, A => n115845, ZN => n115819);
   U88743 : AOI221_X1 port map( B1 => n120085, B2 => n119022, C1 => n120079, C2
                           => n118586, A => n115843, ZN => n115820);
   U88744 : NOR4_X1 port map( A1 => n115837, A2 => n115838, A3 => n115839, A4 
                           => n115840, ZN => n115821);
   U88745 : NAND4_X1 port map( A1 => n115791, A2 => n115792, A3 => n115793, A4 
                           => n115794, ZN => n5421);
   U88746 : AOI221_X1 port map( B1 => n120061, B2 => n119215, C1 => n120055, C2
                           => n118408, A => n115817, ZN => n115791);
   U88747 : AOI221_X1 port map( B1 => n120085, B2 => n119023, C1 => n120079, C2
                           => n118587, A => n115815, ZN => n115792);
   U88748 : NOR4_X1 port map( A1 => n115809, A2 => n115810, A3 => n115811, A4 
                           => n115812, ZN => n115793);
   U88749 : NAND4_X1 port map( A1 => n115763, A2 => n115764, A3 => n115765, A4 
                           => n115766, ZN => n5423);
   U88750 : AOI221_X1 port map( B1 => n120062, B2 => n119216, C1 => n120056, C2
                           => n118409, A => n115789, ZN => n115763);
   U88751 : AOI221_X1 port map( B1 => n120086, B2 => n119024, C1 => n120080, C2
                           => n118588, A => n115787, ZN => n115764);
   U88752 : NOR4_X1 port map( A1 => n115781, A2 => n115782, A3 => n115783, A4 
                           => n115784, ZN => n115765);
   U88753 : NAND4_X1 port map( A1 => n115735, A2 => n115736, A3 => n115737, A4 
                           => n115738, ZN => n5425);
   U88754 : AOI221_X1 port map( B1 => n120062, B2 => n119217, C1 => n120056, C2
                           => n118410, A => n115761, ZN => n115735);
   U88755 : AOI221_X1 port map( B1 => n120086, B2 => n119025, C1 => n120080, C2
                           => n118589, A => n115759, ZN => n115736);
   U88756 : NOR4_X1 port map( A1 => n115753, A2 => n115754, A3 => n115755, A4 
                           => n115756, ZN => n115737);
   U88757 : NAND4_X1 port map( A1 => n115707, A2 => n115708, A3 => n115709, A4 
                           => n115710, ZN => n5427);
   U88758 : AOI221_X1 port map( B1 => n120062, B2 => n119218, C1 => n120056, C2
                           => n118411, A => n115733, ZN => n115707);
   U88759 : AOI221_X1 port map( B1 => n120086, B2 => n119026, C1 => n120080, C2
                           => n118590, A => n115731, ZN => n115708);
   U88760 : NOR4_X1 port map( A1 => n115725, A2 => n115726, A3 => n115727, A4 
                           => n115728, ZN => n115709);
   U88761 : NAND4_X1 port map( A1 => n115679, A2 => n115680, A3 => n115681, A4 
                           => n115682, ZN => n5429);
   U88762 : AOI221_X1 port map( B1 => n120062, B2 => n119219, C1 => n120056, C2
                           => n118412, A => n115705, ZN => n115679);
   U88763 : AOI221_X1 port map( B1 => n120086, B2 => n119027, C1 => n120080, C2
                           => n118591, A => n115703, ZN => n115680);
   U88764 : NOR4_X1 port map( A1 => n115697, A2 => n115698, A3 => n115699, A4 
                           => n115700, ZN => n115681);
   U88765 : NAND4_X1 port map( A1 => n115651, A2 => n115652, A3 => n115653, A4 
                           => n115654, ZN => n5431);
   U88766 : AOI221_X1 port map( B1 => n120062, B2 => n119220, C1 => n120056, C2
                           => n118413, A => n115677, ZN => n115651);
   U88767 : AOI221_X1 port map( B1 => n120086, B2 => n119028, C1 => n120080, C2
                           => n118592, A => n115675, ZN => n115652);
   U88768 : NOR4_X1 port map( A1 => n115669, A2 => n115670, A3 => n115671, A4 
                           => n115672, ZN => n115653);
   U88769 : NAND4_X1 port map( A1 => n115623, A2 => n115624, A3 => n115625, A4 
                           => n115626, ZN => n5433);
   U88770 : AOI221_X1 port map( B1 => n120062, B2 => n119221, C1 => n120056, C2
                           => n118414, A => n115649, ZN => n115623);
   U88771 : AOI221_X1 port map( B1 => n120086, B2 => n119029, C1 => n120080, C2
                           => n118593, A => n115647, ZN => n115624);
   U88772 : NOR4_X1 port map( A1 => n115641, A2 => n115642, A3 => n115643, A4 
                           => n115644, ZN => n115625);
   U88773 : NAND4_X1 port map( A1 => n115595, A2 => n115596, A3 => n115597, A4 
                           => n115598, ZN => n5435);
   U88774 : AOI221_X1 port map( B1 => n120062, B2 => n119222, C1 => n120056, C2
                           => n118415, A => n115621, ZN => n115595);
   U88775 : AOI221_X1 port map( B1 => n120086, B2 => n119030, C1 => n120080, C2
                           => n118594, A => n115619, ZN => n115596);
   U88776 : NOR4_X1 port map( A1 => n115613, A2 => n115614, A3 => n115615, A4 
                           => n115616, ZN => n115597);
   U88777 : NAND4_X1 port map( A1 => n115567, A2 => n115568, A3 => n115569, A4 
                           => n115570, ZN => n5437);
   U88778 : AOI221_X1 port map( B1 => n120062, B2 => n119223, C1 => n120056, C2
                           => n118416, A => n115593, ZN => n115567);
   U88779 : AOI221_X1 port map( B1 => n120086, B2 => n119031, C1 => n120080, C2
                           => n118595, A => n115591, ZN => n115568);
   U88780 : NOR4_X1 port map( A1 => n115585, A2 => n115586, A3 => n115587, A4 
                           => n115588, ZN => n115569);
   U88781 : NAND4_X1 port map( A1 => n115539, A2 => n115540, A3 => n115541, A4 
                           => n115542, ZN => n5439);
   U88782 : AOI221_X1 port map( B1 => n120062, B2 => n119224, C1 => n120056, C2
                           => n118417, A => n115565, ZN => n115539);
   U88783 : AOI221_X1 port map( B1 => n120086, B2 => n119032, C1 => n120080, C2
                           => n118596, A => n115563, ZN => n115540);
   U88784 : NOR4_X1 port map( A1 => n115557, A2 => n115558, A3 => n115559, A4 
                           => n115560, ZN => n115541);
   U88785 : NAND4_X1 port map( A1 => n115511, A2 => n115512, A3 => n115513, A4 
                           => n115514, ZN => n5441);
   U88786 : AOI221_X1 port map( B1 => n120062, B2 => n119225, C1 => n120056, C2
                           => n118418, A => n115537, ZN => n115511);
   U88787 : AOI221_X1 port map( B1 => n120086, B2 => n119033, C1 => n120080, C2
                           => n118597, A => n115535, ZN => n115512);
   U88788 : NOR4_X1 port map( A1 => n115529, A2 => n115530, A3 => n115531, A4 
                           => n115532, ZN => n115513);
   U88789 : NAND4_X1 port map( A1 => n115483, A2 => n115484, A3 => n115485, A4 
                           => n115486, ZN => n5443);
   U88790 : AOI221_X1 port map( B1 => n120062, B2 => n119226, C1 => n120056, C2
                           => n118419, A => n115509, ZN => n115483);
   U88791 : AOI221_X1 port map( B1 => n120086, B2 => n119034, C1 => n120080, C2
                           => n118598, A => n115507, ZN => n115484);
   U88792 : NOR4_X1 port map( A1 => n115501, A2 => n115502, A3 => n115503, A4 
                           => n115504, ZN => n115485);
   U88793 : NAND4_X1 port map( A1 => n115455, A2 => n115456, A3 => n115457, A4 
                           => n115458, ZN => n5445);
   U88794 : AOI221_X1 port map( B1 => n120062, B2 => n119227, C1 => n120056, C2
                           => n118420, A => n115481, ZN => n115455);
   U88795 : AOI221_X1 port map( B1 => n120086, B2 => n119035, C1 => n120080, C2
                           => n118599, A => n115479, ZN => n115456);
   U88796 : NOR4_X1 port map( A1 => n115473, A2 => n115474, A3 => n115475, A4 
                           => n115476, ZN => n115457);
   U88797 : NAND4_X1 port map( A1 => n115427, A2 => n115428, A3 => n115429, A4 
                           => n115430, ZN => n5447);
   U88798 : AOI221_X1 port map( B1 => n120063, B2 => n119228, C1 => n120057, C2
                           => n118421, A => n115453, ZN => n115427);
   U88799 : AOI221_X1 port map( B1 => n120087, B2 => n119036, C1 => n120081, C2
                           => n118600, A => n115451, ZN => n115428);
   U88800 : NOR4_X1 port map( A1 => n115445, A2 => n115446, A3 => n115447, A4 
                           => n115448, ZN => n115429);
   U88801 : NAND4_X1 port map( A1 => n115399, A2 => n115400, A3 => n115401, A4 
                           => n115402, ZN => n5449);
   U88802 : AOI221_X1 port map( B1 => n120063, B2 => n119229, C1 => n120057, C2
                           => n118422, A => n115425, ZN => n115399);
   U88803 : AOI221_X1 port map( B1 => n120087, B2 => n119037, C1 => n120081, C2
                           => n118601, A => n115423, ZN => n115400);
   U88804 : NOR4_X1 port map( A1 => n115417, A2 => n115418, A3 => n115419, A4 
                           => n115420, ZN => n115401);
   U88805 : NAND4_X1 port map( A1 => n115371, A2 => n115372, A3 => n115373, A4 
                           => n115374, ZN => n5451);
   U88806 : AOI221_X1 port map( B1 => n120063, B2 => n119230, C1 => n120057, C2
                           => n118423, A => n115397, ZN => n115371);
   U88807 : AOI221_X1 port map( B1 => n120087, B2 => n119038, C1 => n120081, C2
                           => n118602, A => n115395, ZN => n115372);
   U88808 : NOR4_X1 port map( A1 => n115389, A2 => n115390, A3 => n115391, A4 
                           => n115392, ZN => n115373);
   U88809 : NAND4_X1 port map( A1 => n115343, A2 => n115344, A3 => n115345, A4 
                           => n115346, ZN => n5453);
   U88810 : AOI221_X1 port map( B1 => n120063, B2 => n119231, C1 => n120057, C2
                           => n118424, A => n115369, ZN => n115343);
   U88811 : AOI221_X1 port map( B1 => n120087, B2 => n119039, C1 => n120081, C2
                           => n118603, A => n115367, ZN => n115344);
   U88812 : NOR4_X1 port map( A1 => n115361, A2 => n115362, A3 => n115363, A4 
                           => n115364, ZN => n115345);
   U88813 : NAND4_X1 port map( A1 => n115315, A2 => n115316, A3 => n115317, A4 
                           => n115318, ZN => n5455);
   U88814 : AOI221_X1 port map( B1 => n120063, B2 => n119232, C1 => n120057, C2
                           => n118425, A => n115341, ZN => n115315);
   U88815 : AOI221_X1 port map( B1 => n120087, B2 => n119040, C1 => n120081, C2
                           => n118604, A => n115339, ZN => n115316);
   U88816 : NOR4_X1 port map( A1 => n115333, A2 => n115334, A3 => n115335, A4 
                           => n115336, ZN => n115317);
   U88817 : NAND4_X1 port map( A1 => n115287, A2 => n115288, A3 => n115289, A4 
                           => n115290, ZN => n5457);
   U88818 : AOI221_X1 port map( B1 => n120063, B2 => n119233, C1 => n120057, C2
                           => n118426, A => n115313, ZN => n115287);
   U88819 : AOI221_X1 port map( B1 => n120087, B2 => n119041, C1 => n120081, C2
                           => n118605, A => n115311, ZN => n115288);
   U88820 : NOR4_X1 port map( A1 => n115305, A2 => n115306, A3 => n115307, A4 
                           => n115308, ZN => n115289);
   U88821 : NAND4_X1 port map( A1 => n115259, A2 => n115260, A3 => n115261, A4 
                           => n115262, ZN => n5459);
   U88822 : AOI221_X1 port map( B1 => n120063, B2 => n119234, C1 => n120057, C2
                           => n118427, A => n115285, ZN => n115259);
   U88823 : AOI221_X1 port map( B1 => n120087, B2 => n119042, C1 => n120081, C2
                           => n118606, A => n115283, ZN => n115260);
   U88824 : NOR4_X1 port map( A1 => n115277, A2 => n115278, A3 => n115279, A4 
                           => n115280, ZN => n115261);
   U88825 : NAND4_X1 port map( A1 => n115231, A2 => n115232, A3 => n115233, A4 
                           => n115234, ZN => n5461);
   U88826 : AOI221_X1 port map( B1 => n120063, B2 => n119235, C1 => n120057, C2
                           => n118428, A => n115257, ZN => n115231);
   U88827 : AOI221_X1 port map( B1 => n120087, B2 => n119043, C1 => n120081, C2
                           => n118607, A => n115255, ZN => n115232);
   U88828 : NOR4_X1 port map( A1 => n115249, A2 => n115250, A3 => n115251, A4 
                           => n115252, ZN => n115233);
   U88829 : NAND4_X1 port map( A1 => n115203, A2 => n115204, A3 => n115205, A4 
                           => n115206, ZN => n5463);
   U88830 : AOI221_X1 port map( B1 => n120063, B2 => n119236, C1 => n120057, C2
                           => n118429, A => n115229, ZN => n115203);
   U88831 : AOI221_X1 port map( B1 => n120087, B2 => n119044, C1 => n120081, C2
                           => n118608, A => n115227, ZN => n115204);
   U88832 : NOR4_X1 port map( A1 => n115221, A2 => n115222, A3 => n115223, A4 
                           => n115224, ZN => n115205);
   U88833 : NAND4_X1 port map( A1 => n115175, A2 => n115176, A3 => n115177, A4 
                           => n115178, ZN => n5465);
   U88834 : AOI221_X1 port map( B1 => n120063, B2 => n119237, C1 => n120057, C2
                           => n118430, A => n115201, ZN => n115175);
   U88835 : AOI221_X1 port map( B1 => n120087, B2 => n119045, C1 => n120081, C2
                           => n118609, A => n115199, ZN => n115176);
   U88836 : NOR4_X1 port map( A1 => n115193, A2 => n115194, A3 => n115195, A4 
                           => n115196, ZN => n115177);
   U88837 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n114302);
   U88838 : INV_X1 port map( A => RESET, ZN => n113892);
   U88839 : INV_X1 port map( A => DATAIN(60), ZN => n113771);
   U88840 : INV_X1 port map( A => DATAIN(61), ZN => n113770);
   U88841 : INV_X1 port map( A => DATAIN(62), ZN => n113769);
   U88842 : INV_X1 port map( A => DATAIN(63), ZN => n113768);
   U88843 : INV_X1 port map( A => DATAIN(0), ZN => n113891);
   U88844 : INV_X1 port map( A => DATAIN(1), ZN => n113889);
   U88845 : INV_X1 port map( A => DATAIN(2), ZN => n113887);
   U88846 : INV_X1 port map( A => DATAIN(3), ZN => n113885);
   U88847 : INV_X1 port map( A => DATAIN(4), ZN => n113883);
   U88848 : INV_X1 port map( A => DATAIN(5), ZN => n113881);
   U88849 : INV_X1 port map( A => DATAIN(6), ZN => n113879);
   U88850 : INV_X1 port map( A => DATAIN(7), ZN => n113877);
   U88851 : INV_X1 port map( A => DATAIN(8), ZN => n113875);
   U88852 : INV_X1 port map( A => DATAIN(9), ZN => n113873);
   U88853 : INV_X1 port map( A => DATAIN(10), ZN => n113871);
   U88854 : INV_X1 port map( A => DATAIN(11), ZN => n113869);
   U88855 : INV_X1 port map( A => DATAIN(12), ZN => n113867);
   U88856 : INV_X1 port map( A => DATAIN(13), ZN => n113865);
   U88857 : INV_X1 port map( A => DATAIN(14), ZN => n113863);
   U88858 : INV_X1 port map( A => DATAIN(15), ZN => n113861);
   U88859 : INV_X1 port map( A => DATAIN(16), ZN => n113859);
   U88860 : INV_X1 port map( A => DATAIN(17), ZN => n113857);
   U88861 : INV_X1 port map( A => DATAIN(18), ZN => n113855);
   U88862 : INV_X1 port map( A => DATAIN(19), ZN => n113853);
   U88863 : INV_X1 port map( A => DATAIN(20), ZN => n113851);
   U88864 : INV_X1 port map( A => DATAIN(21), ZN => n113849);
   U88865 : INV_X1 port map( A => DATAIN(22), ZN => n113847);
   U88866 : INV_X1 port map( A => DATAIN(23), ZN => n113845);
   U88867 : INV_X1 port map( A => DATAIN(24), ZN => n113843);
   U88868 : INV_X1 port map( A => DATAIN(25), ZN => n113841);
   U88869 : INV_X1 port map( A => DATAIN(26), ZN => n113839);
   U88870 : INV_X1 port map( A => DATAIN(27), ZN => n113837);
   U88871 : INV_X1 port map( A => DATAIN(28), ZN => n113835);
   U88872 : INV_X1 port map( A => DATAIN(29), ZN => n113833);
   U88873 : INV_X1 port map( A => DATAIN(30), ZN => n113831);
   U88874 : INV_X1 port map( A => DATAIN(31), ZN => n113829);
   U88875 : INV_X1 port map( A => DATAIN(32), ZN => n113827);
   U88876 : INV_X1 port map( A => DATAIN(33), ZN => n113825);
   U88877 : INV_X1 port map( A => DATAIN(34), ZN => n113823);
   U88878 : INV_X1 port map( A => DATAIN(35), ZN => n113821);
   U88879 : INV_X1 port map( A => DATAIN(36), ZN => n113819);
   U88880 : INV_X1 port map( A => DATAIN(37), ZN => n113817);
   U88881 : INV_X1 port map( A => DATAIN(38), ZN => n113815);
   U88882 : INV_X1 port map( A => DATAIN(39), ZN => n113813);
   U88883 : INV_X1 port map( A => DATAIN(40), ZN => n113811);
   U88884 : INV_X1 port map( A => DATAIN(41), ZN => n113809);
   U88885 : INV_X1 port map( A => DATAIN(42), ZN => n113807);
   U88886 : INV_X1 port map( A => DATAIN(43), ZN => n113805);
   U88887 : INV_X1 port map( A => DATAIN(44), ZN => n113803);
   U88888 : INV_X1 port map( A => DATAIN(45), ZN => n113801);
   U88889 : INV_X1 port map( A => DATAIN(46), ZN => n113799);
   U88890 : INV_X1 port map( A => DATAIN(47), ZN => n113797);
   U88891 : INV_X1 port map( A => DATAIN(48), ZN => n113795);
   U88892 : INV_X1 port map( A => DATAIN(49), ZN => n113793);
   U88893 : INV_X1 port map( A => DATAIN(50), ZN => n113791);
   U88894 : INV_X1 port map( A => DATAIN(51), ZN => n113789);
   U88895 : INV_X1 port map( A => DATAIN(52), ZN => n113787);
   U88896 : INV_X1 port map( A => DATAIN(53), ZN => n113785);
   U88897 : INV_X1 port map( A => DATAIN(54), ZN => n113783);
   U88898 : INV_X1 port map( A => DATAIN(55), ZN => n113781);
   U88899 : INV_X1 port map( A => DATAIN(56), ZN => n113779);
   U88900 : INV_X1 port map( A => DATAIN(57), ZN => n113777);
   U88901 : INV_X1 port map( A => DATAIN(58), ZN => n113775);
   U88902 : INV_X1 port map( A => DATAIN(59), ZN => n113773);
   U88903 : INV_X1 port map( A => ADD_WR(3), ZN => n113988);
   U88904 : INV_X1 port map( A => ADD_WR(0), ZN => n113987);
   U88905 : INV_X1 port map( A => ADD_WR(1), ZN => n114376);
   U88906 : INV_X1 port map( A => ADD_RD2(1), ZN => n117973);
   U88907 : INV_X1 port map( A => ADD_RD1(2), ZN => n116475);
   U88908 : INV_X1 port map( A => ADD_RD2(2), ZN => n117971);
   U88909 : INV_X1 port map( A => ADD_RD1(1), ZN => n116478);
   U88910 : INV_X1 port map( A => ADD_WR(2), ZN => n114375);
   U88911 : AND3_X1 port map( A1 => ENABLE, A2 => n114138, A3 => WR, ZN => 
                           n113989);
   U88912 : INV_X1 port map( A => ADD_WR(4), ZN => n114138);
   U88913 : CLKBUF_X1 port map( A => n116532, Z => n119849);
   U88914 : CLKBUF_X1 port map( A => n116531, Z => n119855);
   U88915 : CLKBUF_X1 port map( A => n116529, Z => n119861);
   U88916 : CLKBUF_X1 port map( A => n116528, Z => n119867);
   U88917 : CLKBUF_X1 port map( A => n116527, Z => n119873);
   U88918 : CLKBUF_X1 port map( A => n116526, Z => n119879);
   U88919 : CLKBUF_X1 port map( A => n116523, Z => n119885);
   U88920 : CLKBUF_X1 port map( A => n116522, Z => n119891);
   U88921 : CLKBUF_X1 port map( A => n116521, Z => n119897);
   U88922 : CLKBUF_X1 port map( A => n116520, Z => n119903);
   U88923 : CLKBUF_X1 port map( A => n116519, Z => n119909);
   U88924 : CLKBUF_X1 port map( A => n116518, Z => n119915);
   U88925 : CLKBUF_X1 port map( A => n116517, Z => n119921);
   U88926 : CLKBUF_X1 port map( A => n116516, Z => n119927);
   U88927 : CLKBUF_X1 port map( A => n116515, Z => n119933);
   U88928 : CLKBUF_X1 port map( A => n116514, Z => n119939);
   U88929 : CLKBUF_X1 port map( A => n116513, Z => n119945);
   U88930 : CLKBUF_X1 port map( A => n116508, Z => n119951);
   U88931 : CLKBUF_X1 port map( A => n116507, Z => n119957);
   U88932 : CLKBUF_X1 port map( A => n116505, Z => n119963);
   U88933 : CLKBUF_X1 port map( A => n116504, Z => n119969);
   U88934 : CLKBUF_X1 port map( A => n116503, Z => n119975);
   U88935 : CLKBUF_X1 port map( A => n116502, Z => n119981);
   U88936 : CLKBUF_X1 port map( A => n116500, Z => n119987);
   U88937 : CLKBUF_X1 port map( A => n116499, Z => n119993);
   U88938 : CLKBUF_X1 port map( A => n116497, Z => n119999);
   U88939 : CLKBUF_X1 port map( A => n116495, Z => n120005);
   U88940 : CLKBUF_X1 port map( A => n116493, Z => n120011);
   U88941 : CLKBUF_X1 port map( A => n116492, Z => n120017);
   U88942 : CLKBUF_X1 port map( A => n116491, Z => n120023);
   U88943 : CLKBUF_X1 port map( A => n116490, Z => n120029);
   U88944 : CLKBUF_X1 port map( A => n116488, Z => n120035);
   U88945 : CLKBUF_X1 port map( A => n116487, Z => n120041);
   U88946 : CLKBUF_X1 port map( A => n114703, Z => n120047);
   U88947 : CLKBUF_X1 port map( A => n114702, Z => n120053);
   U88948 : CLKBUF_X1 port map( A => n114700, Z => n120059);
   U88949 : CLKBUF_X1 port map( A => n114698, Z => n120065);
   U88950 : CLKBUF_X1 port map( A => n114697, Z => n120071);
   U88951 : CLKBUF_X1 port map( A => n114696, Z => n120077);
   U88952 : CLKBUF_X1 port map( A => n114693, Z => n120083);
   U88953 : CLKBUF_X1 port map( A => n114691, Z => n120089);
   U88954 : CLKBUF_X1 port map( A => n114690, Z => n120095);
   U88955 : CLKBUF_X1 port map( A => n114689, Z => n120101);
   U88956 : CLKBUF_X1 port map( A => n114688, Z => n120107);
   U88957 : CLKBUF_X1 port map( A => n114687, Z => n120113);
   U88958 : CLKBUF_X1 port map( A => n114686, Z => n120119);
   U88959 : CLKBUF_X1 port map( A => n114685, Z => n120125);
   U88960 : CLKBUF_X1 port map( A => n114684, Z => n120131);
   U88961 : CLKBUF_X1 port map( A => n114683, Z => n120137);
   U88962 : CLKBUF_X1 port map( A => n114682, Z => n120143);
   U88963 : CLKBUF_X1 port map( A => n114676, Z => n120149);
   U88964 : CLKBUF_X1 port map( A => n114675, Z => n120155);
   U88965 : CLKBUF_X1 port map( A => n114673, Z => n120161);
   U88966 : CLKBUF_X1 port map( A => n114672, Z => n120167);
   U88967 : CLKBUF_X1 port map( A => n114670, Z => n120173);
   U88968 : CLKBUF_X1 port map( A => n114669, Z => n120179);
   U88969 : CLKBUF_X1 port map( A => n114667, Z => n120185);
   U88970 : CLKBUF_X1 port map( A => n114666, Z => n120191);
   U88971 : CLKBUF_X1 port map( A => n114664, Z => n120197);
   U88972 : CLKBUF_X1 port map( A => n114662, Z => n120203);
   U88973 : CLKBUF_X1 port map( A => n114660, Z => n120209);
   U88974 : CLKBUF_X1 port map( A => n114659, Z => n120215);
   U88975 : CLKBUF_X1 port map( A => n114658, Z => n120221);
   U88976 : CLKBUF_X1 port map( A => n114657, Z => n120227);
   U88977 : CLKBUF_X1 port map( A => n114655, Z => n120233);
   U88978 : CLKBUF_X1 port map( A => n114654, Z => n120239);
   U88979 : CLKBUF_X1 port map( A => n114645, Z => n120245);
   U88980 : CLKBUF_X1 port map( A => n114579, Z => n120258);
   U88981 : CLKBUF_X1 port map( A => n114576, Z => n120271);
   U88982 : CLKBUF_X1 port map( A => n114575, Z => n120277);
   U88983 : CLKBUF_X1 port map( A => n114511, Z => n120283);
   U88984 : CLKBUF_X1 port map( A => n114445, Z => n120296);
   U88985 : CLKBUF_X1 port map( A => n114379, Z => n120309);
   U88986 : CLKBUF_X1 port map( A => n114373, Z => n120322);
   U88987 : CLKBUF_X1 port map( A => n114372, Z => n120328);
   U88988 : CLKBUF_X1 port map( A => n114307, Z => n120334);
   U88989 : CLKBUF_X1 port map( A => n114304, Z => n120347);
   U88990 : CLKBUF_X1 port map( A => n114303, Z => n120353);
   U88991 : CLKBUF_X1 port map( A => n114301, Z => n120359);
   U88992 : CLKBUF_X1 port map( A => n114300, Z => n120365);
   U88993 : CLKBUF_X1 port map( A => n114236, Z => n120371);
   U88994 : CLKBUF_X1 port map( A => n114214, Z => n120384);
   U88995 : CLKBUF_X1 port map( A => n114213, Z => n120390);
   U88996 : CLKBUF_X1 port map( A => n114212, Z => n120396);
   U88997 : CLKBUF_X1 port map( A => n114211, Z => n120402);
   U88998 : CLKBUF_X1 port map( A => n114147, Z => n120408);
   U88999 : CLKBUF_X1 port map( A => n114143, Z => n120421);
   U89000 : CLKBUF_X1 port map( A => n114142, Z => n120427);
   U89001 : CLKBUF_X1 port map( A => n114140, Z => n120433);
   U89002 : CLKBUF_X1 port map( A => n114139, Z => n120439);
   U89003 : CLKBUF_X1 port map( A => n114137, Z => n120445);
   U89004 : CLKBUF_X1 port map( A => n114136, Z => n120451);
   U89005 : CLKBUF_X1 port map( A => n114135, Z => n120457);
   U89006 : CLKBUF_X1 port map( A => n114134, Z => n120463);
   U89007 : CLKBUF_X1 port map( A => n114133, Z => n120469);
   U89008 : CLKBUF_X1 port map( A => n114132, Z => n120475);
   U89009 : CLKBUF_X1 port map( A => n114131, Z => n120481);
   U89010 : CLKBUF_X1 port map( A => n114130, Z => n120487);
   U89011 : CLKBUF_X1 port map( A => n114129, Z => n120493);
   U89012 : CLKBUF_X1 port map( A => n114128, Z => n120499);
   U89013 : CLKBUF_X1 port map( A => n114124, Z => n120505);
   U89014 : CLKBUF_X1 port map( A => n114122, Z => n120511);
   U89015 : CLKBUF_X1 port map( A => n114057, Z => n120517);
   U89016 : CLKBUF_X1 port map( A => n114053, Z => n120530);
   U89017 : CLKBUF_X1 port map( A => n114052, Z => n120536);
   U89018 : CLKBUF_X1 port map( A => n113991, Z => n120542);
   U89019 : CLKBUF_X1 port map( A => n113982, Z => n120555);
   U89020 : CLKBUF_X1 port map( A => n113980, Z => n120561);
   U89021 : CLKBUF_X1 port map( A => n113916, Z => n120567);
   U89022 : CLKBUF_X1 port map( A => n113912, Z => n120580);
   U89023 : CLKBUF_X1 port map( A => n113911, Z => n120586);
   U89024 : CLKBUF_X1 port map( A => n113910, Z => n120592);
   U89025 : CLKBUF_X1 port map( A => n113909, Z => n120598);
   U89026 : CLKBUF_X1 port map( A => n113904, Z => n120604);
   U89027 : CLKBUF_X1 port map( A => n113902, Z => n120610);
   U89028 : CLKBUF_X1 port map( A => n113897, Z => n120616);
   U89029 : CLKBUF_X1 port map( A => n113895, Z => n120622);
   U89030 : CLKBUF_X1 port map( A => n113892, Z => n120628);
   U89031 : CLKBUF_X1 port map( A => n113767, Z => n120826);

end SYN_behav;
