package CONSTANTS is 
   constant NumBit : integer := 32;	
end CONSTANTS;
