
module registerfile_generic_n_bit32_data_bit64 ( CLK, RESET, ENABLE, RD1, RD2, 
        WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n79527, n89493, n89496,
         n89498, n89500, n89965, n89967, n89968, n89969, n90031, n90033,
         n90034, n90035, n90036, n90037, n90038, n90039, n90040, n90041,
         n90042, n90043, n90044, n90045, n90046, n90047, n90048, n90049,
         n90050, n90051, n90052, n90053, n90054, n90055, n90056, n90057,
         n90058, n90059, n90060, n90061, n90062, n90063, n90064, n90065,
         n90066, n90067, n90068, n90069, n90070, n90071, n90072, n90073,
         n90074, n90075, n90076, n90077, n90078, n90079, n90080, n90081,
         n90082, n90083, n90084, n90085, n90086, n90087, n90088, n90089,
         n90090, n90091, n90092, n90093, n90094, n90095, n90306, n90308,
         n90309, n90310, n90311, n90312, n90313, n90314, n90315, n90316,
         n90317, n90318, n90319, n90320, n90321, n90322, n90323, n90324,
         n90325, n90326, n90327, n90328, n90329, n90330, n90331, n90332,
         n90333, n90334, n90335, n90336, n90337, n90338, n90339, n90340,
         n90341, n90342, n90343, n90344, n90345, n90346, n90347, n90348,
         n90349, n90350, n90351, n90352, n90353, n90354, n90355, n90356,
         n90357, n90358, n90359, n90360, n90361, n90362, n90363, n90364,
         n90365, n90366, n90367, n90368, n90369, n90370, n90373, n90375,
         n90376, n90377, n90378, n90379, n90380, n90381, n90382, n90383,
         n90384, n90385, n90386, n90387, n90388, n90389, n90390, n90391,
         n90392, n90393, n90394, n90395, n90396, n90397, n90398, n90399,
         n90400, n90401, n90402, n90403, n90404, n90405, n90406, n90407,
         n90408, n90409, n90410, n90411, n90412, n90413, n90414, n90415,
         n90416, n90417, n90418, n90419, n90420, n90421, n90422, n90423,
         n90424, n90425, n90426, n90427, n90428, n90429, n90430, n90431,
         n90432, n90433, n90434, n90435, n90436, n90437, n90512, n90514,
         n90515, n90516, n90517, n90518, n90519, n90520, n90521, n90522,
         n90523, n90524, n90525, n90526, n90527, n90528, n90529, n90530,
         n90531, n90532, n90533, n90534, n90535, n90536, n90537, n90538,
         n90539, n90540, n90541, n90542, n90543, n90544, n90545, n90546,
         n90547, n90548, n90549, n90550, n90551, n90552, n90553, n90554,
         n90555, n90556, n90557, n90711, n90713, n90714, n90715, n90716,
         n90717, n90718, n90719, n90720, n90721, n90722, n90723, n90724,
         n90725, n90726, n90727, n90728, n90729, n90730, n90731, n90732,
         n90733, n90734, n90735, n90736, n90737, n90738, n90739, n90740,
         n90741, n90742, n90743, n90744, n90745, n90746, n90747, n90748,
         n90749, n90750, n90751, n90752, n90753, n90754, n90755, n90756,
         n90757, n90758, n90759, n90760, n90761, n90762, n90763, n90764,
         n90765, n90766, n90767, n90768, n90769, n90770, n90771, n90772,
         n90773, n90774, n90775, n95429, n95430, n95431, n95432, n95433,
         n95434, n95435, n95436, n95437, n95438, n95439, n95440, n95441,
         n95442, n95443, n95444, n95445, n95446, n95447, n95448, n95449,
         n95450, n95451, n95452, n95453, n95454, n95455, n95456, n95457,
         n95458, n95459, n95460, n95461, n95462, n95463, n95464, n95465,
         n95466, n95467, n95468, n95469, n95470, n95471, n95472, n95473,
         n95474, n95475, n95476, n95477, n95478, n95479, n95480, n95481,
         n95482, n95483, n95484, n95485, n95486, n95487, n95488, n95525,
         n95526, n95527, n95528, n98523, n98524, n98525, n98526, n98527,
         n98528, n98529, n98530, n98531, n98532, n98533, n98534, n98535,
         n98536, n98537, n98538, n98539, n98540, n98541, n98542, n98543,
         n98544, n98545, n98546, n98547, n98548, n98549, n98550, n98551,
         n98552, n98553, n98554, n98555, n98556, n98557, n98558, n98559,
         n98560, n98561, n98562, n98563, n98564, n98565, n98566, n98567,
         n98568, n98569, n98570, n98571, n98572, n98573, n98574, n98575,
         n98576, n98577, n98578, n98579, n98580, n98581, n98582, n98586,
         n98587, n98588, n98589, n98590, n98591, n98592, n98593, n98594,
         n98595, n98596, n98597, n98598, n98599, n98600, n98601, n98602,
         n98603, n98604, n98605, n98606, n98607, n98608, n98609, n98610,
         n98611, n98612, n98613, n98614, n98615, n98616, n98617, n98618,
         n98619, n98620, n98621, n98622, n98623, n98624, n98625, n98626,
         n98627, n98628, n98629, n98630, n98631, n98632, n98633, n98634,
         n98635, n98636, n98637, n98638, n98639, n98640, n98641, n98642,
         n98643, n98644, n98645, n98648, n98650, n98651, n98652, n98653,
         n98654, n98655, n98656, n98657, n98658, n98659, n98660, n98661,
         n98662, n98663, n98664, n98665, n98666, n98667, n98668, n98669,
         n98670, n98671, n98672, n98673, n98674, n98675, n98676, n98677,
         n98678, n98679, n98680, n98681, n98682, n98683, n98684, n98685,
         n98686, n98687, n98688, n98689, n98690, n98691, n98692, n98693,
         n98694, n98695, n98696, n98697, n98698, n98699, n98700, n98701,
         n98702, n98703, n98704, n98705, n98706, n98707, n98708, n98709,
         n98710, n98711, n98712, n98714, n98716, n98717, n98718, n98719,
         n98720, n98721, n98722, n98723, n98724, n98725, n98726, n98727,
         n98728, n98729, n98730, n98731, n98732, n98733, n98734, n98735,
         n98736, n98737, n98738, n98739, n98740, n98741, n98742, n98743,
         n98744, n98745, n98746, n98747, n98748, n98749, n98750, n98751,
         n98752, n98753, n98754, n98755, n98756, n98757, n98758, n98759,
         n98760, n98761, n98762, n98763, n98764, n98765, n98766, n98767,
         n98768, n98769, n98770, n98771, n98772, n98773, n98774, n98775,
         n98776, n98777, n98778, n98848, n98849, n98850, n98851, n98852,
         n98853, n98854, n98855, n98856, n98857, n98858, n98859, n98860,
         n98861, n98862, n98863, n98864, n98865, n98866, n98867, n98868,
         n98869, n98870, n98871, n98872, n98873, n98874, n98875, n98876,
         n98877, n98878, n98879, n98880, n98881, n98882, n98883, n98884,
         n98885, n98886, n98887, n98888, n98889, n98890, n98891, n98892,
         n98893, n98894, n98895, n98896, n98897, n98898, n98899, n98900,
         n98901, n98902, n98903, n98904, n98905, n98906, n98907, n98986,
         n98987, n98988, n98989, n98990, n98991, n98992, n98993, n98994,
         n98995, n98996, n98997, n98998, n98999, n99000, n99001, n99002,
         n99003, n99004, n99005, n99006, n99007, n99008, n99009, n99010,
         n99011, n99012, n99013, n99014, n99015, n99016, n99017, n99018,
         n99019, n99020, n99021, n99022, n99023, n99024, n99025, n99026,
         n99027, n99028, n99029, n99030, n99031, n99032, n99033, n99034,
         n99035, n99036, n99037, n99038, n99039, n99040, n99041, n99042,
         n99043, n99044, n99045, n99047, n99049, n99050, n99051, n99052,
         n99053, n99054, n99055, n99056, n99057, n99058, n99059, n99060,
         n99061, n99062, n99063, n99064, n99065, n99066, n99067, n99068,
         n99069, n99070, n99071, n99072, n99073, n99074, n99075, n99076,
         n99077, n99078, n99079, n99080, n99081, n99082, n99083, n99084,
         n99085, n99086, n99087, n99088, n99089, n99090, n99091, n99092,
         n99093, n99094, n99095, n99096, n99097, n99098, n99099, n99100,
         n99101, n99102, n99103, n99104, n99105, n99106, n99107, n99108,
         n99109, n99110, n99111, n99113, n99115, n99116, n99117, n99118,
         n99119, n99120, n99121, n99122, n99123, n99124, n99125, n99126,
         n99127, n99128, n99129, n99130, n99131, n99132, n99133, n99134,
         n99135, n99136, n99137, n99138, n99139, n99140, n99141, n99142,
         n99143, n99144, n99145, n99146, n99147, n99148, n99149, n99150,
         n99151, n99152, n99153, n99154, n99155, n99156, n99157, n99158,
         n99159, n99160, n99161, n99162, n99163, n99164, n99165, n99166,
         n99167, n99168, n99169, n99170, n99171, n99172, n99173, n99174,
         n99175, n99176, n99177, n99179, n99181, n99182, n99183, n99184,
         n99185, n99186, n99187, n99188, n99189, n99190, n99191, n99192,
         n99193, n99194, n99195, n99196, n99197, n99198, n99199, n99200,
         n99201, n99202, n99203, n99204, n99205, n99206, n99207, n99208,
         n99209, n99210, n99211, n99212, n99213, n99214, n99215, n99216,
         n99217, n99218, n99219, n99220, n99221, n99222, n99223, n99224,
         n99225, n99226, n99227, n99228, n99229, n99230, n99231, n99232,
         n99233, n99234, n99235, n99236, n99237, n99238, n99239, n99240,
         n99241, n99242, n99243, n99245, n99247, n99248, n99249, n99250,
         n99251, n99252, n99253, n99254, n99255, n99256, n99257, n99258,
         n99259, n99260, n99261, n99262, n99263, n99264, n99265, n99266,
         n99267, n99268, n99269, n99270, n99271, n99272, n99273, n99274,
         n99275, n99276, n99277, n99278, n99279, n99280, n99281, n99282,
         n99283, n99284, n99285, n99286, n99287, n99288, n99289, n99290,
         n99291, n99292, n99293, n99294, n99295, n99296, n99297, n99298,
         n99299, n99300, n99301, n99302, n99303, n99304, n99305, n99306,
         n99307, n99308, n99309, n99311, n99313, n99314, n99315, n99316,
         n99317, n99318, n99319, n99320, n99321, n99322, n99323, n99324,
         n99325, n99326, n99327, n99328, n99329, n99330, n99331, n99332,
         n99333, n99334, n99335, n99336, n99337, n99338, n99339, n99340,
         n99341, n99342, n99343, n99344, n99345, n99346, n99347, n99348,
         n99349, n99350, n99351, n99352, n99353, n99354, n99355, n99356,
         n99357, n99358, n99359, n99360, n99361, n99362, n99363, n99364,
         n99365, n99366, n99367, n99368, n99369, n99370, n99371, n99372,
         n99373, n99374, n99375, n99446, n99448, n99449, n99450, n99451,
         n99452, n99453, n99454, n99455, n99456, n99457, n99458, n99459,
         n99460, n99461, n99462, n99463, n99464, n99465, n99466, n99467,
         n99468, n99469, n99470, n99471, n99472, n99473, n99474, n99475,
         n99476, n99477, n99478, n99479, n99480, n99481, n99482, n99483,
         n99484, n99485, n99486, n99487, n99488, n99489, n99490, n99491,
         n99492, n99493, n99494, n99495, n99496, n99497, n99498, n99499,
         n99500, n99501, n99502, n99503, n99504, n99505, n99506, n99507,
         n99508, n99509, n99510, n99580, n99582, n99583, n99584, n99585,
         n99586, n99587, n99588, n99589, n99590, n99591, n99592, n99593,
         n99594, n99595, n99596, n99597, n99598, n99599, n99600, n99601,
         n99602, n99603, n99604, n99605, n99606, n99607, n99608, n99609,
         n99610, n99611, n99612, n99613, n99614, n99615, n99616, n99617,
         n99618, n99619, n99620, n99621, n99622, n99623, n99624, n99625,
         n99626, n99627, n99628, n99629, n99630, n99631, n99632, n99633,
         n99634, n99635, n99636, n99637, n99638, n99639, n99640, n99641,
         n99642, n99643, n99644, n99716, n99718, n99719, n99720, n99721,
         n99722, n99723, n99724, n99725, n99726, n99727, n99728, n99729,
         n99730, n99731, n99732, n99733, n99734, n99735, n99736, n99737,
         n99738, n99739, n99740, n99741, n99742, n99743, n99744, n99745,
         n99746, n99747, n99748, n99749, n99750, n99751, n99752, n99753,
         n99754, n99755, n99756, n99757, n99758, n99759, n99760, n99761,
         n99762, n99763, n99764, n99765, n99766, n99767, n99768, n99769,
         n99770, n99771, n99772, n99773, n99774, n99775, n99776, n99777,
         n99778, n99779, n99780, n99914, n99916, n99917, n99918, n99919,
         n99920, n99921, n99922, n99923, n99924, n99925, n99926, n99927,
         n99928, n99929, n99930, n99931, n99932, n99933, n99934, n99935,
         n99936, n99937, n99938, n99939, n99940, n99941, n99942, n99943,
         n99944, n99945, n99946, n99947, n99948, n99949, n99950, n99951,
         n99952, n99953, n99954, n99955, n99956, n99957, n99958, n99959,
         n99960, n99961, n99962, n99963, n99964, n99965, n99966, n99967,
         n99968, n99969, n99970, n99971, n99972, n99973, n99974, n99975,
         n99976, n99977, n99978, n109895, n109896, n109897, n109898, n109903,
         n109904, n109905, n109906, n109979, n109980, n109981, n109982,
         n109983, n109984, n109985, n109986, n109987, n109988, n109989,
         n109990, n109991, n109992, n109993, n109994, n109995, n109996,
         n109997, n110107, n110108, n110109, n110110, n110171, n110172,
         n110173, n110174, n110175, n110176, n110177, n110178, n110179,
         n110180, n110181, n110182, n110183, n110184, n110185, n110186,
         n110187, n110188, n110189, n110190, n110191, n110192, n110193,
         n110194, n110195, n110196, n110197, n110198, n110199, n110200,
         n110201, n110202, n110203, n110204, n110205, n110206, n110207,
         n110208, n110209, n110210, n110211, n110212, n110213, n110214,
         n110215, n110216, n110217, n110218, n110219, n110220, n110221,
         n110222, n110223, n110224, n110225, n110226, n110227, n110228,
         n110229, n110230, n110231, n110232, n110233, n110234, n110363,
         n110364, n110365, n110366, n110431, n110432, n110433, n110434,
         n110435, n110436, n110437, n110438, n110439, n110440, n110441,
         n110442, n110443, n110444, n110445, n110446, n110447, n110448,
         n110449, n110450, n110451, n110452, n110453, n110454, n110455,
         n110456, n110457, n110458, n110459, n110460, n110461, n110462,
         n110463, n110464, n110465, n110466, n110467, n110468, n110469,
         n110470, n110471, n110472, n110473, n110474, n110475, n110476,
         n110477, n110478, n110479, n110480, n110481, n110482, n110483,
         n110484, n110485, n110486, n110487, n110488, n110489, n110490,
         n110491, n110492, n110493, n110494, n110495, n110496, n110497,
         n110498, n110499, n110500, n110501, n110502, n110503, n110504,
         n110505, n110506, n110507, n110508, n110509, n110510, n110511,
         n110512, n110513, n110514, n110515, n110516, n110517, n110518,
         n110519, n110520, n110521, n110522, n110523, n110524, n110525,
         n110526, n110527, n110528, n110529, n110530, n110531, n110532,
         n110533, n110534, n110535, n110536, n110537, n110538, n110539,
         n110540, n110541, n110542, n110543, n110544, n110545, n110546,
         n110547, n110548, n110549, n110550, n110551, n110552, n110553,
         n110554, n110555, n110556, n110557, n110558, n110559, n110560,
         n110561, n110562, n110563, n110564, n110565, n110566, n110567,
         n110568, n110569, n110570, n110571, n110572, n110573, n110574,
         n110575, n110576, n110577, n110578, n110579, n110580, n110581,
         n110582, n110583, n110584, n110585, n110586, n110587, n110588,
         n110589, n110590, n110591, n110592, n110593, n110594, n110595,
         n110596, n110597, n110598, n110599, n110600, n110601, n110602,
         n110603, n110604, n110605, n110606, n110607, n110608, n110609,
         n110610, n110611, n110612, n110613, n110614, n110615, n110616,
         n110617, n110618, n110619, n110620, n110621, n110622, n110811,
         n110812, n110813, n110814, n110815, n110816, n110817, n110818,
         n110819, n110820, n110821, n110822, n110823, n110824, n110825,
         n110826, n110827, n110828, n110829, n110830, n110831, n110832,
         n110833, n110834, n110835, n110836, n110837, n110838, n110839,
         n110840, n110841, n110842, n110843, n110844, n110845, n110846,
         n110847, n110848, n110849, n110850, n110851, n110852, n110853,
         n110854, n110855, n110856, n110857, n110858, n110859, n110860,
         n110861, n110862, n110863, n110864, n110865, n110866, n110867,
         n110868, n110869, n110870, n110871, n110872, n110873, n110874,
         n110996, n110997, n110998, n110999, n111000, n111001, n111002,
         n111003, n111004, n111005, n111006, n111007, n111008, n111009,
         n111010, n111011, n111012, n111013, n111014, n111015, n111016,
         n111017, n111018, n111019, n111020, n111021, n111022, n111023,
         n111024, n111025, n111026, n111027, n111028, n111029, n111030,
         n111031, n111032, n111033, n111034, n111035, n111036, n111037,
         n111038, n111039, n111040, n111041, n111042, n111043, n111044,
         n111045, n111046, n111047, n111048, n113766, n113767, n113768,
         n113769, n113770, n113771, n113772, n113773, n113774, n113775,
         n113776, n113777, n113778, n113779, n113780, n113781, n113782,
         n113783, n113784, n113785, n113786, n113787, n113788, n113789,
         n113790, n113791, n113792, n113793, n113794, n113795, n113796,
         n113797, n113798, n113799, n113800, n113801, n113802, n113803,
         n113804, n113805, n113806, n113807, n113808, n113809, n113810,
         n113811, n113812, n113813, n113814, n113815, n113816, n113817,
         n113818, n113819, n113820, n113821, n113822, n113823, n113824,
         n113825, n113826, n113827, n113828, n113829, n113830, n113831,
         n113832, n113833, n113834, n113835, n113836, n113837, n113838,
         n113839, n113840, n113841, n113842, n113843, n113844, n113845,
         n113846, n113847, n113848, n113849, n113850, n113851, n113852,
         n113853, n113854, n113855, n113856, n113857, n113858, n113859,
         n113860, n113861, n113862, n113863, n113864, n113865, n113866,
         n113867, n113868, n113869, n113870, n113871, n113872, n113873,
         n113874, n113875, n113876, n113877, n113878, n113879, n113880,
         n113881, n113882, n113883, n113884, n113885, n113886, n113887,
         n113888, n113889, n113890, n113891, n113892, n113893, n113894,
         n113895, n113896, n113897, n113898, n113899, n113900, n113901,
         n113902, n113903, n113904, n113905, n113906, n113907, n113908,
         n113909, n113910, n113911, n113912, n113913, n113914, n113915,
         n113916, n113917, n113918, n113919, n113920, n113921, n113922,
         n113923, n113924, n113925, n113926, n113927, n113928, n113929,
         n113930, n113931, n113932, n113933, n113934, n113935, n113936,
         n113937, n113938, n113939, n113940, n113941, n113942, n113943,
         n113944, n113945, n113946, n113947, n113948, n113949, n113950,
         n113951, n113952, n113953, n113954, n113955, n113956, n113957,
         n113958, n113959, n113960, n113961, n113962, n113963, n113964,
         n113965, n113966, n113967, n113968, n113969, n113970, n113971,
         n113972, n113973, n113974, n113975, n113976, n113977, n113978,
         n113979, n113980, n113981, n113982, n113983, n113984, n113985,
         n113986, n113987, n113988, n113989, n113990, n113991, n113992,
         n113993, n113994, n113995, n113996, n113997, n113998, n113999,
         n114000, n114001, n114002, n114003, n114004, n114005, n114006,
         n114007, n114008, n114009, n114010, n114011, n114012, n114013,
         n114014, n114015, n114016, n114017, n114018, n114019, n114020,
         n114021, n114022, n114023, n114024, n114025, n114026, n114027,
         n114028, n114029, n114030, n114031, n114032, n114033, n114034,
         n114035, n114036, n114037, n114038, n114039, n114040, n114041,
         n114042, n114043, n114044, n114045, n114046, n114047, n114048,
         n114049, n114050, n114051, n114052, n114053, n114054, n114055,
         n114056, n114057, n114058, n114059, n114060, n114061, n114062,
         n114063, n114064, n114065, n114066, n114067, n114068, n114069,
         n114070, n114071, n114072, n114073, n114074, n114075, n114076,
         n114077, n114078, n114079, n114080, n114081, n114082, n114083,
         n114084, n114085, n114086, n114087, n114088, n114089, n114090,
         n114091, n114092, n114093, n114094, n114095, n114096, n114097,
         n114098, n114099, n114100, n114101, n114102, n114103, n114104,
         n114105, n114106, n114107, n114108, n114109, n114110, n114111,
         n114112, n114113, n114114, n114115, n114116, n114117, n114118,
         n114119, n114120, n114121, n114122, n114123, n114124, n114125,
         n114126, n114127, n114128, n114129, n114130, n114131, n114132,
         n114133, n114134, n114135, n114136, n114137, n114138, n114139,
         n114140, n114141, n114142, n114143, n114144, n114145, n114146,
         n114147, n114148, n114149, n114150, n114151, n114152, n114153,
         n114154, n114155, n114156, n114157, n114158, n114159, n114160,
         n114161, n114162, n114163, n114164, n114165, n114166, n114167,
         n114168, n114169, n114170, n114171, n114172, n114173, n114174,
         n114175, n114176, n114177, n114178, n114179, n114180, n114181,
         n114182, n114183, n114184, n114185, n114186, n114187, n114188,
         n114189, n114190, n114191, n114192, n114193, n114194, n114195,
         n114196, n114197, n114198, n114199, n114200, n114201, n114202,
         n114203, n114204, n114205, n114206, n114207, n114208, n114209,
         n114210, n114211, n114212, n114213, n114214, n114215, n114216,
         n114217, n114218, n114219, n114220, n114221, n114222, n114223,
         n114224, n114225, n114226, n114227, n114228, n114229, n114230,
         n114231, n114232, n114233, n114234, n114235, n114236, n114237,
         n114238, n114239, n114240, n114241, n114242, n114243, n114244,
         n114245, n114246, n114247, n114248, n114249, n114250, n114251,
         n114252, n114253, n114254, n114255, n114256, n114257, n114258,
         n114259, n114260, n114261, n114262, n114263, n114264, n114265,
         n114266, n114267, n114268, n114269, n114270, n114271, n114272,
         n114273, n114274, n114275, n114276, n114277, n114278, n114279,
         n114280, n114281, n114282, n114283, n114284, n114285, n114286,
         n114287, n114288, n114289, n114290, n114291, n114292, n114293,
         n114294, n114295, n114296, n114297, n114298, n114299, n114300,
         n114301, n114302, n114303, n114304, n114305, n114306, n114307,
         n114308, n114309, n114310, n114311, n114312, n114313, n114314,
         n114315, n114316, n114317, n114318, n114319, n114320, n114321,
         n114322, n114323, n114324, n114325, n114326, n114327, n114328,
         n114329, n114330, n114331, n114332, n114333, n114334, n114335,
         n114336, n114337, n114338, n114339, n114340, n114341, n114342,
         n114343, n114344, n114345, n114346, n114347, n114348, n114349,
         n114350, n114351, n114352, n114353, n114354, n114355, n114356,
         n114357, n114358, n114359, n114360, n114361, n114362, n114363,
         n114364, n114365, n114366, n114367, n114368, n114369, n114370,
         n114371, n114372, n114373, n114374, n114375, n114376, n114377,
         n114378, n114379, n114380, n114381, n114382, n114383, n114384,
         n114385, n114386, n114387, n114388, n114389, n114390, n114391,
         n114392, n114393, n114394, n114395, n114396, n114397, n114398,
         n114399, n114400, n114401, n114402, n114403, n114404, n114405,
         n114406, n114407, n114408, n114409, n114410, n114411, n114412,
         n114413, n114414, n114415, n114416, n114417, n114418, n114419,
         n114420, n114421, n114422, n114423, n114424, n114425, n114426,
         n114427, n114428, n114429, n114430, n114431, n114432, n114433,
         n114434, n114435, n114436, n114437, n114438, n114439, n114440,
         n114441, n114442, n114443, n114444, n114445, n114446, n114447,
         n114448, n114449, n114450, n114451, n114452, n114453, n114454,
         n114455, n114456, n114457, n114458, n114459, n114460, n114461,
         n114462, n114463, n114464, n114465, n114466, n114467, n114468,
         n114469, n114470, n114471, n114472, n114473, n114474, n114475,
         n114476, n114477, n114478, n114479, n114480, n114481, n114482,
         n114483, n114484, n114485, n114486, n114487, n114488, n114489,
         n114490, n114491, n114492, n114493, n114494, n114495, n114496,
         n114497, n114498, n114499, n114500, n114501, n114502, n114503,
         n114504, n114505, n114506, n114507, n114508, n114509, n114510,
         n114511, n114512, n114513, n114514, n114515, n114516, n114517,
         n114518, n114519, n114520, n114521, n114522, n114523, n114524,
         n114525, n114526, n114527, n114528, n114529, n114530, n114531,
         n114532, n114533, n114534, n114535, n114536, n114537, n114538,
         n114539, n114540, n114541, n114542, n114543, n114544, n114545,
         n114546, n114547, n114548, n114549, n114550, n114551, n114552,
         n114553, n114554, n114555, n114556, n114557, n114558, n114559,
         n114560, n114561, n114562, n114563, n114564, n114565, n114566,
         n114567, n114568, n114569, n114570, n114571, n114572, n114573,
         n114574, n114575, n114576, n114577, n114578, n114579, n114580,
         n114581, n114582, n114583, n114584, n114585, n114586, n114587,
         n114588, n114589, n114590, n114591, n114592, n114593, n114594,
         n114595, n114596, n114597, n114598, n114599, n114600, n114601,
         n114602, n114603, n114604, n114605, n114606, n114607, n114608,
         n114609, n114610, n114611, n114612, n114613, n114614, n114615,
         n114616, n114617, n114618, n114619, n114620, n114621, n114622,
         n114623, n114624, n114625, n114626, n114627, n114628, n114629,
         n114630, n114631, n114632, n114633, n114634, n114635, n114636,
         n114637, n114638, n114639, n114640, n114641, n114642, n114643,
         n114644, n114645, n114646, n114647, n114648, n114649, n114650,
         n114651, n114652, n114653, n114654, n114655, n114656, n114657,
         n114658, n114659, n114660, n114661, n114662, n114664, n114666,
         n114667, n114668, n114669, n114670, n114672, n114673, n114674,
         n114675, n114676, n114678, n114679, n114680, n114681, n114682,
         n114683, n114684, n114685, n114686, n114687, n114688, n114689,
         n114690, n114691, n114693, n114695, n114696, n114697, n114698,
         n114700, n114701, n114702, n114703, n114704, n114705, n114706,
         n114707, n114708, n114709, n114710, n114711, n114712, n114713,
         n114714, n114717, n114719, n114721, n114722, n114723, n114724,
         n114727, n114729, n114730, n114731, n114732, n114733, n114734,
         n114735, n114736, n114737, n114738, n114739, n114740, n114743,
         n114745, n114747, n114748, n114749, n114750, n114753, n114755,
         n114756, n114757, n114758, n114759, n114760, n114761, n114762,
         n114763, n114764, n114765, n114766, n114769, n114771, n114773,
         n114774, n114775, n114776, n114779, n114781, n114782, n114783,
         n114784, n114785, n114786, n114787, n114788, n114789, n114790,
         n114791, n114793, n114796, n114798, n114801, n114802, n114803,
         n114804, n114807, n114809, n114810, n114811, n114812, n114813,
         n114814, n114815, n114816, n114817, n114818, n114819, n114821,
         n114824, n114826, n114829, n114830, n114831, n114832, n114835,
         n114837, n114838, n114839, n114840, n114841, n114842, n114843,
         n114844, n114845, n114846, n114847, n114849, n114852, n114854,
         n114857, n114858, n114859, n114860, n114863, n114865, n114866,
         n114867, n114868, n114869, n114870, n114871, n114872, n114873,
         n114874, n114875, n114877, n114880, n114882, n114885, n114886,
         n114887, n114888, n114891, n114893, n114894, n114895, n114896,
         n114897, n114898, n114899, n114900, n114901, n114902, n114903,
         n114905, n114908, n114910, n114913, n114914, n114915, n114916,
         n114919, n114921, n114922, n114923, n114924, n114925, n114926,
         n114927, n114928, n114929, n114930, n114931, n114933, n114936,
         n114938, n114941, n114942, n114943, n114944, n114947, n114949,
         n114950, n114951, n114952, n114953, n114954, n114955, n114956,
         n114957, n114958, n114959, n114961, n114964, n114966, n114969,
         n114970, n114971, n114972, n114975, n114977, n114978, n114979,
         n114980, n114981, n114982, n114983, n114984, n114985, n114986,
         n114987, n114989, n114992, n114994, n114997, n114998, n114999,
         n115000, n115003, n115005, n115006, n115007, n115008, n115009,
         n115010, n115011, n115012, n115013, n115014, n115015, n115017,
         n115020, n115022, n115025, n115026, n115027, n115028, n115031,
         n115033, n115034, n115035, n115036, n115037, n115038, n115039,
         n115040, n115041, n115042, n115043, n115045, n115048, n115050,
         n115053, n115054, n115055, n115056, n115059, n115061, n115062,
         n115063, n115064, n115065, n115066, n115067, n115068, n115069,
         n115070, n115071, n115073, n115076, n115078, n115081, n115082,
         n115083, n115084, n115087, n115089, n115090, n115091, n115092,
         n115093, n115094, n115095, n115096, n115097, n115098, n115099,
         n115101, n115104, n115106, n115109, n115110, n115111, n115112,
         n115115, n115117, n115118, n115119, n115120, n115121, n115122,
         n115123, n115124, n115125, n115126, n115127, n115129, n115132,
         n115134, n115137, n115138, n115139, n115140, n115143, n115145,
         n115146, n115147, n115148, n115149, n115150, n115151, n115152,
         n115153, n115154, n115155, n115157, n115160, n115162, n115165,
         n115166, n115167, n115168, n115171, n115173, n115174, n115175,
         n115176, n115177, n115178, n115179, n115180, n115181, n115182,
         n115183, n115185, n115188, n115190, n115193, n115194, n115195,
         n115196, n115199, n115201, n115202, n115203, n115204, n115205,
         n115206, n115207, n115208, n115209, n115210, n115211, n115213,
         n115216, n115218, n115221, n115222, n115223, n115224, n115227,
         n115229, n115230, n115231, n115232, n115233, n115234, n115235,
         n115236, n115237, n115238, n115239, n115241, n115244, n115246,
         n115249, n115250, n115251, n115252, n115255, n115257, n115258,
         n115259, n115260, n115261, n115262, n115263, n115264, n115265,
         n115266, n115267, n115269, n115272, n115274, n115277, n115278,
         n115279, n115280, n115283, n115285, n115286, n115287, n115288,
         n115289, n115290, n115291, n115292, n115293, n115294, n115295,
         n115297, n115300, n115302, n115305, n115306, n115307, n115308,
         n115311, n115313, n115314, n115315, n115316, n115317, n115318,
         n115319, n115320, n115321, n115322, n115323, n115325, n115328,
         n115330, n115333, n115334, n115335, n115336, n115339, n115341,
         n115342, n115343, n115344, n115345, n115346, n115347, n115348,
         n115349, n115350, n115351, n115353, n115356, n115358, n115361,
         n115362, n115363, n115364, n115367, n115369, n115370, n115371,
         n115372, n115373, n115374, n115375, n115376, n115377, n115378,
         n115379, n115381, n115384, n115386, n115389, n115390, n115391,
         n115392, n115395, n115397, n115398, n115399, n115400, n115401,
         n115402, n115403, n115404, n115405, n115406, n115407, n115409,
         n115412, n115414, n115417, n115418, n115419, n115420, n115423,
         n115425, n115426, n115427, n115428, n115429, n115430, n115431,
         n115432, n115433, n115434, n115435, n115437, n115440, n115442,
         n115445, n115446, n115447, n115448, n115451, n115453, n115454,
         n115455, n115456, n115457, n115458, n115459, n115460, n115461,
         n115462, n115463, n115465, n115468, n115470, n115473, n115474,
         n115475, n115476, n115479, n115481, n115482, n115483, n115484,
         n115485, n115486, n115487, n115488, n115489, n115490, n115491,
         n115493, n115496, n115498, n115501, n115502, n115503, n115504,
         n115507, n115509, n115510, n115511, n115512, n115513, n115514,
         n115515, n115516, n115517, n115518, n115519, n115521, n115524,
         n115526, n115529, n115530, n115531, n115532, n115535, n115537,
         n115538, n115539, n115540, n115541, n115542, n115543, n115544,
         n115545, n115546, n115547, n115549, n115552, n115554, n115557,
         n115558, n115559, n115560, n115563, n115565, n115566, n115567,
         n115568, n115569, n115570, n115571, n115572, n115573, n115574,
         n115575, n115577, n115580, n115582, n115585, n115586, n115587,
         n115588, n115591, n115593, n115594, n115595, n115596, n115597,
         n115598, n115599, n115600, n115601, n115602, n115603, n115605,
         n115608, n115610, n115613, n115614, n115615, n115616, n115619,
         n115621, n115622, n115623, n115624, n115625, n115626, n115627,
         n115628, n115629, n115630, n115631, n115633, n115636, n115638,
         n115641, n115642, n115643, n115644, n115647, n115649, n115650,
         n115651, n115652, n115653, n115654, n115655, n115656, n115657,
         n115658, n115659, n115661, n115664, n115666, n115669, n115670,
         n115671, n115672, n115675, n115677, n115678, n115679, n115680,
         n115681, n115682, n115683, n115684, n115685, n115686, n115687,
         n115689, n115692, n115694, n115697, n115698, n115699, n115700,
         n115703, n115705, n115706, n115707, n115708, n115709, n115710,
         n115711, n115712, n115713, n115714, n115715, n115717, n115720,
         n115722, n115725, n115726, n115727, n115728, n115731, n115733,
         n115734, n115735, n115736, n115737, n115738, n115739, n115740,
         n115741, n115742, n115743, n115745, n115748, n115750, n115753,
         n115754, n115755, n115756, n115759, n115761, n115762, n115763,
         n115764, n115765, n115766, n115767, n115768, n115769, n115770,
         n115771, n115773, n115776, n115778, n115781, n115782, n115783,
         n115784, n115787, n115789, n115790, n115791, n115792, n115793,
         n115794, n115795, n115796, n115797, n115798, n115799, n115801,
         n115804, n115806, n115809, n115810, n115811, n115812, n115815,
         n115817, n115818, n115819, n115820, n115821, n115822, n115823,
         n115824, n115825, n115826, n115827, n115829, n115832, n115834,
         n115837, n115838, n115839, n115840, n115843, n115845, n115846,
         n115847, n115848, n115849, n115850, n115851, n115852, n115853,
         n115854, n115855, n115857, n115860, n115862, n115865, n115866,
         n115867, n115868, n115871, n115873, n115874, n115875, n115876,
         n115877, n115878, n115879, n115880, n115881, n115882, n115883,
         n115885, n115888, n115890, n115893, n115894, n115895, n115896,
         n115899, n115901, n115902, n115903, n115904, n115905, n115906,
         n115907, n115908, n115909, n115910, n115911, n115913, n115916,
         n115918, n115921, n115922, n115923, n115924, n115927, n115929,
         n115930, n115931, n115932, n115933, n115934, n115935, n115936,
         n115937, n115938, n115939, n115941, n115944, n115946, n115949,
         n115950, n115951, n115952, n115955, n115957, n115958, n115959,
         n115960, n115961, n115962, n115963, n115964, n115965, n115966,
         n115967, n115969, n115972, n115974, n115977, n115978, n115979,
         n115980, n115983, n115985, n115986, n115987, n115988, n115989,
         n115990, n115991, n115992, n115993, n115994, n115995, n115997,
         n116000, n116002, n116005, n116006, n116007, n116008, n116011,
         n116013, n116014, n116015, n116016, n116017, n116018, n116019,
         n116020, n116021, n116022, n116023, n116025, n116028, n116030,
         n116033, n116034, n116035, n116036, n116039, n116041, n116042,
         n116043, n116044, n116045, n116046, n116047, n116048, n116049,
         n116050, n116051, n116053, n116056, n116058, n116061, n116062,
         n116063, n116064, n116067, n116069, n116070, n116071, n116072,
         n116073, n116074, n116075, n116076, n116077, n116078, n116079,
         n116081, n116084, n116086, n116089, n116090, n116091, n116092,
         n116095, n116097, n116098, n116099, n116100, n116101, n116102,
         n116103, n116104, n116105, n116106, n116107, n116109, n116112,
         n116114, n116117, n116118, n116119, n116120, n116123, n116125,
         n116126, n116127, n116128, n116129, n116130, n116131, n116132,
         n116133, n116134, n116135, n116137, n116140, n116142, n116145,
         n116146, n116147, n116148, n116151, n116153, n116154, n116155,
         n116156, n116157, n116158, n116159, n116160, n116161, n116162,
         n116163, n116165, n116168, n116170, n116173, n116174, n116175,
         n116176, n116179, n116181, n116182, n116183, n116184, n116185,
         n116186, n116187, n116188, n116189, n116190, n116191, n116193,
         n116196, n116198, n116201, n116202, n116203, n116204, n116207,
         n116209, n116210, n116211, n116212, n116213, n116214, n116215,
         n116216, n116217, n116218, n116219, n116221, n116224, n116226,
         n116229, n116230, n116231, n116232, n116235, n116237, n116238,
         n116239, n116240, n116241, n116242, n116243, n116244, n116245,
         n116246, n116247, n116249, n116252, n116254, n116257, n116258,
         n116259, n116260, n116263, n116265, n116266, n116267, n116268,
         n116269, n116270, n116271, n116272, n116273, n116274, n116275,
         n116277, n116280, n116282, n116285, n116286, n116287, n116288,
         n116291, n116293, n116294, n116295, n116296, n116297, n116298,
         n116299, n116300, n116301, n116302, n116303, n116305, n116308,
         n116310, n116313, n116314, n116315, n116316, n116319, n116321,
         n116322, n116323, n116324, n116325, n116326, n116327, n116328,
         n116329, n116330, n116331, n116333, n116336, n116338, n116341,
         n116342, n116343, n116344, n116347, n116349, n116350, n116351,
         n116352, n116353, n116354, n116355, n116356, n116357, n116358,
         n116359, n116361, n116364, n116366, n116369, n116370, n116371,
         n116372, n116375, n116377, n116378, n116379, n116380, n116381,
         n116382, n116383, n116384, n116385, n116386, n116387, n116389,
         n116392, n116394, n116397, n116398, n116399, n116400, n116403,
         n116405, n116406, n116407, n116408, n116409, n116410, n116411,
         n116412, n116413, n116414, n116415, n116417, n116420, n116422,
         n116425, n116426, n116427, n116428, n116431, n116433, n116434,
         n116435, n116436, n116437, n116438, n116439, n116440, n116441,
         n116442, n116443, n116445, n116446, n116447, n116448, n116449,
         n116452, n116453, n116454, n116455, n116457, n116458, n116459,
         n116460, n116463, n116464, n116465, n116466, n116467, n116468,
         n116469, n116470, n116471, n116474, n116475, n116477, n116478,
         n116479, n116480, n116481, n116482, n116483, n116484, n116485,
         n116486, n116487, n116488, n116489, n116490, n116491, n116492,
         n116493, n116494, n116495, n116497, n116499, n116500, n116501,
         n116502, n116503, n116504, n116505, n116506, n116507, n116508,
         n116509, n116510, n116511, n116512, n116513, n116514, n116515,
         n116516, n116517, n116518, n116519, n116520, n116521, n116522,
         n116523, n116525, n116526, n116527, n116528, n116529, n116530,
         n116531, n116532, n116533, n116534, n116535, n116536, n116537,
         n116538, n116539, n116540, n116541, n116542, n116545, n116546,
         n116547, n116548, n116549, n116550, n116552, n116553, n116554,
         n116555, n116556, n116557, n116558, n116559, n116560, n116561,
         n116562, n116563, n116566, n116567, n116568, n116569, n116570,
         n116571, n116573, n116574, n116575, n116576, n116577, n116578,
         n116579, n116580, n116581, n116582, n116583, n116584, n116587,
         n116588, n116589, n116590, n116591, n116592, n116594, n116595,
         n116596, n116597, n116598, n116599, n116600, n116601, n116602,
         n116603, n116604, n116606, n116609, n116611, n116612, n116613,
         n116614, n116615, n116617, n116618, n116619, n116620, n116621,
         n116622, n116623, n116624, n116625, n116626, n116627, n116629,
         n116632, n116634, n116635, n116636, n116637, n116638, n116640,
         n116641, n116642, n116643, n116644, n116645, n116646, n116647,
         n116648, n116649, n116650, n116652, n116655, n116657, n116658,
         n116659, n116660, n116661, n116663, n116664, n116665, n116666,
         n116667, n116668, n116669, n116670, n116671, n116672, n116673,
         n116675, n116678, n116680, n116681, n116682, n116683, n116684,
         n116686, n116687, n116688, n116689, n116690, n116691, n116692,
         n116693, n116694, n116695, n116696, n116698, n116701, n116703,
         n116704, n116705, n116706, n116707, n116709, n116710, n116711,
         n116712, n116713, n116714, n116715, n116716, n116717, n116718,
         n116719, n116721, n116724, n116726, n116727, n116728, n116729,
         n116730, n116732, n116733, n116734, n116735, n116736, n116737,
         n116738, n116739, n116740, n116741, n116742, n116744, n116747,
         n116749, n116750, n116751, n116752, n116753, n116755, n116756,
         n116757, n116758, n116759, n116760, n116761, n116762, n116763,
         n116764, n116765, n116767, n116770, n116772, n116773, n116774,
         n116775, n116776, n116778, n116779, n116780, n116781, n116782,
         n116783, n116784, n116785, n116786, n116787, n116788, n116790,
         n116793, n116795, n116796, n116797, n116798, n116799, n116801,
         n116802, n116803, n116804, n116805, n116806, n116807, n116808,
         n116809, n116810, n116811, n116813, n116816, n116818, n116819,
         n116820, n116821, n116822, n116824, n116825, n116826, n116827,
         n116828, n116829, n116830, n116831, n116832, n116833, n116834,
         n116836, n116839, n116841, n116842, n116843, n116844, n116845,
         n116847, n116848, n116849, n116850, n116851, n116852, n116853,
         n116854, n116855, n116856, n116857, n116859, n116862, n116864,
         n116865, n116866, n116867, n116868, n116870, n116871, n116872,
         n116873, n116874, n116875, n116876, n116877, n116878, n116879,
         n116880, n116882, n116885, n116887, n116888, n116889, n116890,
         n116891, n116893, n116894, n116895, n116896, n116897, n116898,
         n116899, n116900, n116901, n116902, n116903, n116905, n116908,
         n116910, n116911, n116912, n116913, n116914, n116916, n116917,
         n116918, n116919, n116920, n116921, n116922, n116923, n116924,
         n116925, n116926, n116928, n116931, n116933, n116934, n116935,
         n116936, n116937, n116939, n116940, n116941, n116942, n116943,
         n116944, n116945, n116946, n116947, n116948, n116949, n116951,
         n116954, n116956, n116957, n116958, n116959, n116960, n116962,
         n116963, n116964, n116965, n116966, n116967, n116968, n116969,
         n116970, n116971, n116972, n116974, n116977, n116979, n116980,
         n116981, n116982, n116983, n116985, n116986, n116987, n116988,
         n116989, n116990, n116991, n116992, n116993, n116994, n116995,
         n116997, n117000, n117002, n117003, n117004, n117005, n117006,
         n117008, n117009, n117010, n117011, n117012, n117013, n117014,
         n117015, n117016, n117017, n117018, n117020, n117023, n117025,
         n117026, n117027, n117028, n117029, n117031, n117032, n117033,
         n117034, n117035, n117036, n117037, n117038, n117039, n117040,
         n117041, n117043, n117046, n117048, n117049, n117050, n117051,
         n117052, n117054, n117055, n117056, n117057, n117058, n117059,
         n117060, n117061, n117062, n117063, n117064, n117066, n117069,
         n117071, n117072, n117073, n117074, n117075, n117077, n117078,
         n117079, n117080, n117081, n117082, n117083, n117084, n117085,
         n117086, n117087, n117089, n117092, n117094, n117095, n117096,
         n117097, n117098, n117100, n117101, n117102, n117103, n117104,
         n117105, n117106, n117107, n117108, n117109, n117110, n117112,
         n117115, n117117, n117118, n117119, n117120, n117121, n117123,
         n117124, n117125, n117126, n117127, n117128, n117129, n117130,
         n117131, n117132, n117133, n117135, n117138, n117140, n117141,
         n117142, n117143, n117144, n117146, n117147, n117148, n117149,
         n117150, n117151, n117152, n117153, n117154, n117155, n117156,
         n117158, n117161, n117163, n117164, n117165, n117166, n117167,
         n117169, n117170, n117171, n117172, n117173, n117174, n117175,
         n117176, n117177, n117178, n117179, n117181, n117184, n117186,
         n117187, n117188, n117189, n117190, n117192, n117193, n117194,
         n117195, n117196, n117197, n117198, n117199, n117200, n117201,
         n117202, n117204, n117207, n117209, n117210, n117211, n117212,
         n117213, n117215, n117216, n117217, n117218, n117219, n117220,
         n117221, n117222, n117223, n117224, n117225, n117227, n117230,
         n117232, n117233, n117234, n117235, n117236, n117238, n117239,
         n117240, n117241, n117242, n117243, n117244, n117245, n117246,
         n117247, n117248, n117250, n117253, n117255, n117256, n117257,
         n117258, n117259, n117261, n117262, n117263, n117264, n117265,
         n117266, n117267, n117268, n117269, n117270, n117271, n117273,
         n117276, n117278, n117279, n117280, n117281, n117282, n117284,
         n117285, n117286, n117287, n117288, n117289, n117290, n117291,
         n117292, n117293, n117294, n117296, n117299, n117301, n117302,
         n117303, n117304, n117305, n117307, n117308, n117309, n117310,
         n117311, n117312, n117313, n117314, n117315, n117316, n117317,
         n117319, n117322, n117324, n117325, n117326, n117327, n117328,
         n117330, n117331, n117332, n117333, n117334, n117335, n117336,
         n117337, n117338, n117339, n117340, n117342, n117345, n117347,
         n117348, n117349, n117350, n117351, n117353, n117354, n117355,
         n117356, n117357, n117358, n117359, n117360, n117361, n117362,
         n117363, n117365, n117368, n117370, n117371, n117372, n117373,
         n117374, n117376, n117377, n117378, n117379, n117380, n117381,
         n117382, n117383, n117384, n117385, n117386, n117388, n117391,
         n117393, n117394, n117395, n117396, n117397, n117399, n117400,
         n117401, n117402, n117403, n117404, n117405, n117406, n117407,
         n117408, n117409, n117411, n117414, n117416, n117417, n117418,
         n117419, n117420, n117422, n117423, n117424, n117425, n117426,
         n117427, n117428, n117429, n117430, n117431, n117432, n117434,
         n117437, n117439, n117440, n117441, n117442, n117443, n117445,
         n117446, n117447, n117448, n117449, n117450, n117451, n117452,
         n117453, n117454, n117455, n117457, n117460, n117462, n117463,
         n117464, n117465, n117466, n117468, n117469, n117470, n117471,
         n117472, n117473, n117474, n117475, n117476, n117477, n117478,
         n117480, n117483, n117485, n117486, n117487, n117488, n117489,
         n117491, n117492, n117493, n117494, n117495, n117496, n117497,
         n117498, n117499, n117500, n117501, n117503, n117506, n117508,
         n117509, n117510, n117511, n117512, n117514, n117515, n117516,
         n117517, n117518, n117519, n117520, n117521, n117522, n117523,
         n117524, n117526, n117529, n117531, n117532, n117533, n117534,
         n117535, n117537, n117538, n117539, n117540, n117541, n117542,
         n117543, n117544, n117545, n117546, n117547, n117549, n117552,
         n117554, n117555, n117556, n117557, n117558, n117559, n117560,
         n117561, n117562, n117563, n117564, n117565, n117566, n117567,
         n117568, n117569, n117571, n117574, n117576, n117577, n117578,
         n117579, n117580, n117581, n117582, n117583, n117584, n117585,
         n117586, n117587, n117588, n117589, n117590, n117591, n117593,
         n117596, n117598, n117599, n117600, n117601, n117602, n117603,
         n117604, n117605, n117606, n117607, n117608, n117609, n117610,
         n117611, n117612, n117613, n117615, n117618, n117620, n117621,
         n117622, n117623, n117624, n117625, n117626, n117627, n117628,
         n117629, n117630, n117631, n117632, n117633, n117634, n117635,
         n117637, n117640, n117642, n117643, n117644, n117645, n117646,
         n117647, n117648, n117649, n117650, n117651, n117652, n117653,
         n117654, n117655, n117656, n117657, n117659, n117662, n117664,
         n117665, n117666, n117667, n117668, n117669, n117670, n117671,
         n117672, n117673, n117674, n117675, n117676, n117677, n117678,
         n117679, n117681, n117684, n117686, n117687, n117688, n117689,
         n117690, n117691, n117692, n117693, n117694, n117695, n117696,
         n117697, n117698, n117699, n117700, n117701, n117703, n117706,
         n117708, n117709, n117710, n117711, n117712, n117713, n117714,
         n117715, n117716, n117717, n117718, n117719, n117720, n117721,
         n117722, n117723, n117725, n117728, n117730, n117731, n117732,
         n117733, n117734, n117735, n117736, n117737, n117738, n117739,
         n117740, n117741, n117742, n117743, n117744, n117745, n117747,
         n117750, n117752, n117753, n117754, n117755, n117756, n117757,
         n117758, n117759, n117760, n117761, n117762, n117763, n117764,
         n117765, n117766, n117767, n117769, n117772, n117774, n117775,
         n117776, n117777, n117778, n117779, n117780, n117781, n117782,
         n117783, n117784, n117785, n117786, n117787, n117788, n117789,
         n117791, n117794, n117796, n117797, n117798, n117799, n117800,
         n117801, n117802, n117803, n117804, n117805, n117806, n117807,
         n117808, n117809, n117810, n117811, n117813, n117816, n117818,
         n117819, n117820, n117821, n117822, n117823, n117824, n117825,
         n117826, n117827, n117828, n117829, n117830, n117831, n117832,
         n117833, n117835, n117838, n117840, n117841, n117842, n117843,
         n117844, n117845, n117846, n117847, n117848, n117849, n117850,
         n117851, n117852, n117853, n117854, n117855, n117857, n117860,
         n117862, n117863, n117864, n117865, n117866, n117867, n117868,
         n117869, n117870, n117871, n117872, n117873, n117874, n117875,
         n117876, n117877, n117879, n117882, n117884, n117885, n117886,
         n117887, n117888, n117889, n117890, n117891, n117892, n117893,
         n117894, n117895, n117896, n117897, n117898, n117899, n117901,
         n117904, n117906, n117907, n117908, n117909, n117910, n117911,
         n117912, n117913, n117914, n117915, n117916, n117917, n117918,
         n117919, n117920, n117921, n117923, n117926, n117928, n117929,
         n117930, n117931, n117932, n117933, n117934, n117935, n117936,
         n117937, n117938, n117939, n117940, n117941, n117942, n117943,
         n117945, n117946, n117947, n117948, n117949, n117950, n117953,
         n117954, n117955, n117956, n117958, n117959, n117960, n117961,
         n117962, n117963, n117964, n117965, n117966, n117967, n117968,
         n117969, n117970, n117971, n117972, n117973, n117974, n117975,
         n117976, n117977, n117981, n117982, n117983, n117984, n117985,
         n117986, n117987, n117988, n117993, n117994, n117995, n117996,
         n118070, n118071, n118072, n118073, n118074, n118075, n118076,
         n118077, n118078, n118079, n118080, n118081, n118082, n118083,
         n118084, n118205, n118206, n118207, n118208, n118209, n118210,
         n118211, n118212, n118213, n118214, n118215, n118216, n118217,
         n118218, n118219, n118220, n118221, n118222, n118223, n118224,
         n118225, n118226, n118227, n118228, n118229, n118230, n118231,
         n118232, n118233, n118234, n118235, n118236, n118237, n118238,
         n118239, n118240, n118241, n118242, n118243, n118244, n118245,
         n118246, n118247, n118248, n118249, n118250, n118251, n118252,
         n118253, n118254, n118255, n118256, n118257, n118258, n118259,
         n118260, n118261, n118262, n118263, n118264, n118325, n118326,
         n118327, n118328, n118329, n118330, n118331, n118332, n118333,
         n118334, n118335, n118336, n118337, n118338, n118339, n118340,
         n118341, n118342, n118343, n118344, n118345, n118346, n118347,
         n118348, n118349, n118350, n118351, n118352, n118353, n118354,
         n118355, n118356, n118357, n118358, n118359, n118360, n118361,
         n118362, n118363, n118364, n118365, n118366, n118367, n118368,
         n118369, n118370, n118371, n118372, n118373, n118374, n118375,
         n118376, n118377, n118378, n118379, n118380, n118381, n118382,
         n118383, n118384, n118385, n118386, n118387, n118388, n118389,
         n118390, n118391, n118392, n118393, n118394, n118395, n118396,
         n118397, n118398, n118399, n118400, n118401, n118402, n118403,
         n118404, n118405, n118406, n118407, n118408, n118409, n118410,
         n118411, n118412, n118413, n118414, n118415, n118416, n118417,
         n118418, n118419, n118420, n118421, n118422, n118423, n118424,
         n118425, n118426, n118427, n118428, n118429, n118430, n118431,
         n118432, n118433, n118434, n118435, n118436, n118437, n118438,
         n118439, n118440, n118441, n118442, n118443, n118444, n118505,
         n118506, n118507, n118508, n118509, n118510, n118511, n118512,
         n118513, n118514, n118515, n118516, n118517, n118518, n118519,
         n118520, n118521, n118522, n118523, n118524, n118525, n118526,
         n118527, n118528, n118529, n118530, n118531, n118532, n118533,
         n118534, n118535, n118536, n118537, n118538, n118539, n118540,
         n118541, n118542, n118543, n118544, n118545, n118546, n118547,
         n118548, n118549, n118550, n118551, n118552, n118553, n118554,
         n118555, n118556, n118557, n118558, n118559, n118560, n118561,
         n118562, n118563, n118564, n118565, n118566, n118567, n118568,
         n118569, n118570, n118571, n118572, n118573, n118574, n118575,
         n118576, n118577, n118578, n118579, n118580, n118581, n118582,
         n118583, n118584, n118585, n118586, n118587, n118588, n118589,
         n118590, n118591, n118592, n118593, n118594, n118595, n118596,
         n118597, n118598, n118599, n118600, n118601, n118602, n118603,
         n118604, n118605, n118606, n118607, n118608, n118609, n118610,
         n118611, n118612, n118613, n118614, n118615, n118616, n118617,
         n118618, n118619, n118620, n118621, n118622, n118623, n118624,
         n118625, n118626, n118627, n118628, n118629, n118630, n118631,
         n118632, n118633, n118634, n118635, n118636, n118637, n118638,
         n118639, n118640, n118641, n118642, n118643, n118644, n118645,
         n118646, n118647, n118648, n118649, n118650, n118651, n118652,
         n118653, n118654, n118655, n118656, n118657, n118658, n118659,
         n118660, n118661, n118662, n118663, n118664, n118665, n118666,
         n118667, n118668, n118669, n118670, n118671, n118672, n118673,
         n118674, n118675, n118676, n118677, n118678, n118679, n118680,
         n118681, n118682, n118683, n118684, n118685, n118686, n118687,
         n118688, n118689, n118690, n118691, n118692, n118693, n118694,
         n118695, n118696, n118697, n118698, n118699, n118700, n118701,
         n118702, n118703, n118704, n118705, n118706, n118707, n118708,
         n118709, n118710, n118711, n118712, n118713, n118714, n118715,
         n118716, n118717, n118718, n118719, n118720, n118721, n118722,
         n118723, n118724, n118725, n118726, n118727, n118728, n118729,
         n118730, n118731, n118732, n118733, n118734, n118735, n118736,
         n118737, n118738, n118739, n118740, n118741, n118742, n118743,
         n118744, n118745, n118746, n118747, n118748, n118749, n118750,
         n118751, n118752, n118753, n118754, n118755, n118756, n118757,
         n118758, n118759, n118760, n118761, n118762, n118763, n118764,
         n118765, n118766, n118767, n118768, n118769, n118770, n118771,
         n118772, n118773, n118774, n118775, n118776, n118777, n118778,
         n118779, n118780, n118781, n118782, n118783, n118784, n118785,
         n118786, n118787, n118788, n118789, n118790, n118791, n118792,
         n118793, n118794, n118795, n118796, n118797, n118798, n118799,
         n118800, n118801, n118802, n118803, n118804, n118805, n118806,
         n118807, n118808, n118809, n118810, n118811, n118812, n118813,
         n118814, n118815, n118816, n118817, n118818, n118819, n118820,
         n118821, n118822, n118823, n118824, n118825, n118826, n118827,
         n118828, n118829, n118830, n118831, n118832, n118833, n118834,
         n118835, n118836, n118837, n118838, n118839, n118840, n118841,
         n118842, n118843, n118844, n118845, n118846, n118847, n118848,
         n118849, n118850, n118851, n118852, n118853, n118854, n118855,
         n118856, n118857, n118858, n118859, n118860, n118861, n118862,
         n118863, n118864, n118865, n118866, n118867, n118868, n118869,
         n118870, n118871, n118872, n118873, n118874, n118875, n118876,
         n118877, n118878, n118879, n118880, n118881, n118882, n118883,
         n118884, n118885, n118886, n118887, n118888, n118889, n118890,
         n118891, n118892, n118893, n118894, n118895, n118896, n118897,
         n118898, n118899, n118900, n118901, n118902, n118903, n118904,
         n118905, n118906, n118907, n118908, n118909, n118910, n118911,
         n118912, n118913, n118914, n118915, n118916, n118917, n118918,
         n118919, n118920, n118921, n118922, n118923, n118924, n118925,
         n118926, n118927, n118928, n118929, n118930, n118931, n118932,
         n118933, n118934, n118935, n118936, n118937, n118938, n118939,
         n118940, n118941, n118942, n118943, n118944, n118945, n118946,
         n118947, n118948, n118949, n118950, n118951, n118952, n118953,
         n118954, n118955, n118956, n118957, n118958, n118959, n118960,
         n118961, n118962, n118963, n118964, n118965, n118966, n118967,
         n118968, n118969, n118970, n118971, n118972, n118973, n118974,
         n118975, n118976, n118977, n118978, n118979, n118980, n118981,
         n118982, n118983, n118984, n118985, n118986, n118987, n118988,
         n118989, n118990, n118991, n118992, n118993, n118994, n118995,
         n118996, n118997, n118998, n118999, n119000, n119001, n119002,
         n119003, n119004, n119005, n119006, n119007, n119008, n119009,
         n119010, n119011, n119012, n119013, n119014, n119015, n119016,
         n119017, n119018, n119019, n119020, n119021, n119022, n119023,
         n119024, n119025, n119026, n119027, n119028, n119029, n119030,
         n119031, n119032, n119033, n119034, n119035, n119036, n119037,
         n119038, n119039, n119040, n119041, n119042, n119043, n119044,
         n119045, n119046, n119047, n119048, n119049, n119050, n119051,
         n119052, n119053, n119054, n119055, n119056, n119057, n119058,
         n119059, n119060, n119061, n119062, n119063, n119064, n119065,
         n119066, n119067, n119068, n119069, n119070, n119071, n119072,
         n119073, n119074, n119075, n119076, n119077, n119078, n119079,
         n119080, n119081, n119082, n119083, n119084, n119085, n119086,
         n119087, n119088, n119089, n119090, n119091, n119092, n119093,
         n119094, n119095, n119096, n119097, n119098, n119099, n119100,
         n119101, n119102, n119103, n119104, n119105, n119106, n119107,
         n119108, n119109, n119110, n119111, n119112, n119113, n119114,
         n119115, n119116, n119117, n119118, n119119, n119120, n119121,
         n119122, n119123, n119124, n119125, n119126, n119127, n119128,
         n119129, n119130, n119131, n119132, n119133, n119134, n119135,
         n119136, n119137, n119138, n119139, n119140, n119141, n119142,
         n119143, n119144, n119145, n119146, n119147, n119148, n119149,
         n119150, n119151, n119152, n119153, n119154, n119155, n119156,
         n119157, n119158, n119159, n119160, n119161, n119162, n119163,
         n119164, n119165, n119166, n119167, n119168, n119169, n119170,
         n119171, n119172, n119173, n119174, n119175, n119176, n119177,
         n119178, n119179, n119180, n119181, n119182, n119183, n119184,
         n119185, n119186, n119187, n119188, n119189, n119190, n119191,
         n119192, n119193, n119194, n119195, n119196, n119197, n119198,
         n119199, n119200, n119201, n119202, n119203, n119204, n119205,
         n119206, n119207, n119208, n119209, n119210, n119211, n119212,
         n119213, n119214, n119215, n119216, n119217, n119218, n119219,
         n119220, n119221, n119222, n119223, n119224, n119225, n119226,
         n119227, n119228, n119229, n119230, n119231, n119232, n119233,
         n119234, n119235, n119236, n119237, n119238, n119239, n119240,
         n119241, n119242, n119243, n119244, n119245, n119246, n119247,
         n119248, n119249, n119250, n119251, n119252, n119253, n119254,
         n119255, n119256, n119257, n119258, n119259, n119260, n119261,
         n119262, n119263, n119264, n119265, n119266, n119267, n119268,
         n119269, n119270, n119271, n119272, n119273, n119274, n119275,
         n119276, n119277, n119278, n119279, n119280, n119281, n119282,
         n119283, n119284, n119285, n119286, n119287, n119288, n119289,
         n119290, n119291, n119292, n119293, n119294, n119295, n119296,
         n119297, n119298, n119299, n119300, n119301, n119302, n119303,
         n119304, n119305, n119306, n119307, n119308, n119309, n119310,
         n119311, n119312, n119313, n119314, n119315, n119316, n119317,
         n119318, n119319, n119320, n119321, n119322, n119323, n119324,
         n119325, n119326, n119327, n119328, n119329, n119330, n119331,
         n119332, n119333, n119334, n119335, n119336, n119337, n119338,
         n119339, n119340, n119341, n119342, n119343, n119344, n119345,
         n119346, n119347, n119348, n119349, n119350, n119351, n119352,
         n119353, n119354, n119355, n119356, n119357, n119358, n119359,
         n119360, n119361, n119362, n119363, n119364, n119365, n119844,
         n119845, n119846, n119847, n119848, n119849, n119850, n119851,
         n119852, n119853, n119854, n119855, n119856, n119857, n119858,
         n119859, n119860, n119861, n119862, n119863, n119864, n119865,
         n119866, n119867, n119868, n119869, n119870, n119871, n119872,
         n119873, n119874, n119875, n119876, n119877, n119878, n119879,
         n119880, n119881, n119882, n119883, n119884, n119885, n119886,
         n119887, n119888, n119889, n119890, n119891, n119892, n119893,
         n119894, n119895, n119896, n119897, n119898, n119899, n119900,
         n119901, n119902, n119903, n119904, n119905, n119906, n119907,
         n119908, n119909, n119910, n119911, n119912, n119913, n119914,
         n119915, n119916, n119917, n119918, n119919, n119920, n119921,
         n119922, n119923, n119924, n119925, n119926, n119927, n119928,
         n119929, n119930, n119931, n119932, n119933, n119934, n119935,
         n119936, n119937, n119938, n119939, n119940, n119941, n119942,
         n119943, n119944, n119945, n119946, n119947, n119948, n119949,
         n119950, n119951, n119952, n119953, n119954, n119955, n119956,
         n119957, n119958, n119959, n119960, n119961, n119962, n119963,
         n119964, n119965, n119966, n119967, n119968, n119969, n119970,
         n119971, n119972, n119973, n119974, n119975, n119976, n119977,
         n119978, n119979, n119980, n119981, n119982, n119983, n119984,
         n119985, n119986, n119987, n119988, n119989, n119990, n119991,
         n119992, n119993, n119994, n119995, n119996, n119997, n119998,
         n119999, n120000, n120001, n120002, n120003, n120004, n120005,
         n120006, n120007, n120008, n120009, n120010, n120011, n120012,
         n120013, n120014, n120015, n120016, n120017, n120018, n120019,
         n120020, n120021, n120022, n120023, n120024, n120025, n120026,
         n120027, n120028, n120029, n120030, n120031, n120032, n120033,
         n120034, n120035, n120036, n120037, n120038, n120039, n120040,
         n120041, n120042, n120043, n120044, n120045, n120046, n120047,
         n120048, n120049, n120050, n120051, n120052, n120053, n120054,
         n120055, n120056, n120057, n120058, n120059, n120060, n120061,
         n120062, n120063, n120064, n120065, n120066, n120067, n120068,
         n120069, n120070, n120071, n120072, n120073, n120074, n120075,
         n120076, n120077, n120078, n120079, n120080, n120081, n120082,
         n120083, n120084, n120085, n120086, n120087, n120088, n120089,
         n120090, n120091, n120092, n120093, n120094, n120095, n120096,
         n120097, n120098, n120099, n120100, n120101, n120102, n120103,
         n120104, n120105, n120106, n120107, n120108, n120109, n120110,
         n120111, n120112, n120113, n120114, n120115, n120116, n120117,
         n120118, n120119, n120120, n120121, n120122, n120123, n120124,
         n120125, n120126, n120127, n120128, n120129, n120130, n120131,
         n120132, n120133, n120134, n120135, n120136, n120137, n120138,
         n120139, n120140, n120141, n120142, n120143, n120144, n120145,
         n120146, n120147, n120148, n120149, n120150, n120151, n120152,
         n120153, n120154, n120155, n120156, n120157, n120158, n120159,
         n120160, n120161, n120162, n120163, n120164, n120165, n120166,
         n120167, n120168, n120169, n120170, n120171, n120172, n120173,
         n120174, n120175, n120176, n120177, n120178, n120179, n120180,
         n120181, n120182, n120183, n120184, n120185, n120186, n120187,
         n120188, n120189, n120190, n120191, n120192, n120193, n120194,
         n120195, n120196, n120197, n120198, n120199, n120200, n120201,
         n120202, n120203, n120204, n120205, n120206, n120207, n120208,
         n120209, n120210, n120211, n120212, n120213, n120214, n120215,
         n120216, n120217, n120218, n120219, n120220, n120221, n120222,
         n120223, n120224, n120225, n120226, n120227, n120228, n120229,
         n120230, n120231, n120232, n120233, n120234, n120235, n120236,
         n120237, n120238, n120239, n120240, n120241, n120242, n120243,
         n120244, n120245, n120246, n120247, n120248, n120249, n120250,
         n120251, n120252, n120253, n120254, n120255, n120256, n120257,
         n120258, n120259, n120260, n120261, n120262, n120263, n120264,
         n120265, n120266, n120267, n120268, n120269, n120270, n120271,
         n120272, n120273, n120274, n120275, n120276, n120277, n120278,
         n120279, n120280, n120281, n120282, n120283, n120284, n120285,
         n120286, n120287, n120288, n120289, n120290, n120291, n120292,
         n120293, n120294, n120295, n120296, n120297, n120298, n120299,
         n120300, n120301, n120302, n120303, n120304, n120305, n120306,
         n120307, n120308, n120309, n120310, n120311, n120312, n120313,
         n120314, n120315, n120316, n120317, n120318, n120319, n120320,
         n120321, n120322, n120323, n120324, n120325, n120326, n120327,
         n120328, n120329, n120330, n120331, n120332, n120333, n120334,
         n120335, n120336, n120337, n120338, n120339, n120340, n120341,
         n120342, n120343, n120344, n120345, n120346, n120347, n120348,
         n120349, n120350, n120351, n120352, n120353, n120354, n120355,
         n120356, n120357, n120358, n120359, n120360, n120361, n120362,
         n120363, n120364, n120365, n120366, n120367, n120368, n120369,
         n120370, n120371, n120372, n120373, n120374, n120375, n120376,
         n120377, n120378, n120379, n120380, n120381, n120382, n120383,
         n120384, n120385, n120386, n120387, n120388, n120389, n120390,
         n120391, n120392, n120393, n120394, n120395, n120396, n120397,
         n120398, n120399, n120400, n120401, n120402, n120403, n120404,
         n120405, n120406, n120407, n120408, n120409, n120410, n120411,
         n120412, n120413, n120414, n120415, n120416, n120417, n120418,
         n120419, n120420, n120421, n120422, n120423, n120424, n120425,
         n120426, n120427, n120428, n120429, n120430, n120431, n120432,
         n120433, n120434, n120435, n120436, n120437, n120438, n120439,
         n120440, n120441, n120442, n120443, n120444, n120445, n120446,
         n120447, n120448, n120449, n120450, n120451, n120452, n120453,
         n120454, n120455, n120456, n120457, n120458, n120459, n120460,
         n120461, n120462, n120463, n120464, n120465, n120466, n120467,
         n120468, n120469, n120470, n120471, n120472, n120473, n120474,
         n120475, n120476, n120477, n120478, n120479, n120480, n120481,
         n120482, n120483, n120484, n120485, n120486, n120487, n120488,
         n120489, n120490, n120491, n120492, n120493, n120494, n120495,
         n120496, n120497, n120498, n120499, n120500, n120501, n120502,
         n120503, n120504, n120505, n120506, n120507, n120508, n120509,
         n120510, n120511, n120512, n120513, n120514, n120515, n120516,
         n120517, n120518, n120519, n120520, n120521, n120522, n120523,
         n120524, n120525, n120526, n120527, n120528, n120529, n120530,
         n120531, n120532, n120533, n120534, n120535, n120536, n120537,
         n120538, n120539, n120540, n120541, n120542, n120543, n120544,
         n120545, n120546, n120547, n120548, n120549, n120550, n120551,
         n120552, n120553, n120554, n120555, n120556, n120557, n120558,
         n120559, n120560, n120561, n120562, n120563, n120564, n120565,
         n120566, n120567, n120568, n120569, n120570, n120571, n120572,
         n120573, n120574, n120575, n120576, n120577, n120578, n120579,
         n120580, n120581, n120582, n120583, n120584, n120585, n120586,
         n120587, n120588, n120589, n120590, n120591, n120592, n120593,
         n120594, n120595, n120596, n120597, n120598, n120599, n120600,
         n120601, n120602, n120603, n120604, n120605, n120606, n120607,
         n120608, n120609, n120610, n120611, n120612, n120613, n120614,
         n120615, n120616, n120617, n120618, n120619, n120620, n120621,
         n120622, n120623, n120624, n120625, n120626, n120627, n120628,
         n120629, n120630, n120631, n120632, n120633, n120634, n120635,
         n120636, n120637, n120638, n120639, n120640, n120641, n120642,
         n120643, n120644, n120645, n120646, n120647, n120648, n120649,
         n120650, n120651, n120652, n120653, n120654, n120655, n120656,
         n120657, n120658, n120659, n120660, n120661, n120662, n120663,
         n120664, n120665, n120666, n120667, n120668, n120669, n120670,
         n120671, n120672, n120673, n120674, n120675, n120676, n120677,
         n120678, n120679, n120680, n120681, n120682, n120683, n120684,
         n120685, n120686, n120687, n120688, n120689, n120690, n120691,
         n120692, n120693, n120694, n120695, n120696, n120697, n120698,
         n120699, n120700, n120701, n120702, n120703, n120704, n120705,
         n120706, n120707, n120708, n120709, n120710, n120711, n120712,
         n120713, n120714, n120715, n120716, n120717, n120718, n120719,
         n120720, n120721, n120722, n120723, n120724, n120725, n120726,
         n120727, n120728, n120729, n120730, n120731, n120732, n120733,
         n120734, n120735, n120736, n120737, n120738, n120739, n120740,
         n120741, n120742, n120743, n120744, n120745, n120746, n120747,
         n120748, n120749, n120750, n120751, n120752, n120753, n120754,
         n120755, n120756, n120757, n120758, n120759, n120760, n120761,
         n120762, n120763, n120764, n120765, n120766, n120767, n120768,
         n120769, n120770, n120771, n120772, n120773, n120774, n120775,
         n120776, n120777, n120778, n120779, n120780, n120781, n120782,
         n120783, n120784, n120785, n120786, n120787, n120788, n120789,
         n120790, n120791, n120792, n120793, n120794, n120795, n120796,
         n120797, n120798, n120799, n120800, n120801, n120802, n120803,
         n120804, n120805, n120806, n120807, n120808, n120809, n120810,
         n120811, n120812, n120813, n120814, n120815, n120816, n120817,
         n120818, n120819, n120820, n120821, n120822, n120823, n120824,
         n120825, n120826, n120827, n120828, n120829, n120830, n120831,
         n120832, n120833;
  assign n79527 = CLK;

  DFF_X1 \OUT1_reg[45]  ( .D(n5465), .CK(n79527), .Q(OUT1[45]) );
  DFF_X1 \OUT1_reg[44]  ( .D(n5463), .CK(n79527), .Q(OUT1[44]) );
  DFF_X1 \OUT1_reg[43]  ( .D(n5461), .CK(n79527), .Q(OUT1[43]) );
  DFF_X1 \OUT1_reg[42]  ( .D(n5459), .CK(n79527), .Q(OUT1[42]) );
  DFF_X1 \OUT1_reg[41]  ( .D(n5457), .CK(n79527), .Q(OUT1[41]) );
  DFF_X1 \OUT1_reg[40]  ( .D(n5455), .CK(n79527), .Q(OUT1[40]) );
  DFF_X1 \OUT1_reg[39]  ( .D(n5453), .CK(n79527), .Q(OUT1[39]) );
  DFF_X1 \OUT1_reg[38]  ( .D(n5451), .CK(n79527), .Q(OUT1[38]) );
  DFF_X1 \OUT1_reg[37]  ( .D(n5449), .CK(n79527), .Q(OUT1[37]) );
  DFF_X1 \OUT1_reg[36]  ( .D(n5447), .CK(n79527), .Q(OUT1[36]) );
  DFF_X1 \OUT1_reg[35]  ( .D(n5445), .CK(n79527), .Q(OUT1[35]) );
  DFF_X1 \OUT1_reg[34]  ( .D(n5443), .CK(n79527), .Q(OUT1[34]) );
  DFF_X1 \OUT1_reg[33]  ( .D(n5441), .CK(n79527), .Q(OUT1[33]) );
  DFF_X1 \OUT1_reg[32]  ( .D(n5439), .CK(n79527), .Q(OUT1[32]) );
  DFF_X1 \OUT1_reg[31]  ( .D(n5437), .CK(n79527), .Q(OUT1[31]) );
  DFF_X1 \OUT1_reg[30]  ( .D(n5435), .CK(n79527), .Q(OUT1[30]) );
  DFF_X1 \OUT1_reg[29]  ( .D(n5433), .CK(n79527), .Q(OUT1[29]) );
  DFF_X1 \OUT1_reg[28]  ( .D(n5431), .CK(n79527), .Q(OUT1[28]) );
  DFF_X1 \OUT1_reg[27]  ( .D(n5429), .CK(n79527), .Q(OUT1[27]) );
  DFF_X1 \OUT1_reg[26]  ( .D(n5427), .CK(n79527), .Q(OUT1[26]) );
  DFF_X1 \OUT1_reg[25]  ( .D(n5425), .CK(n79527), .Q(OUT1[25]) );
  DFF_X1 \OUT1_reg[24]  ( .D(n5423), .CK(n79527), .Q(OUT1[24]) );
  DFF_X1 \OUT1_reg[23]  ( .D(n5421), .CK(n79527), .Q(OUT1[23]) );
  DFF_X1 \OUT1_reg[22]  ( .D(n5419), .CK(n79527), .Q(OUT1[22]) );
  DFF_X1 \OUT1_reg[21]  ( .D(n5417), .CK(n79527), .Q(OUT1[21]) );
  DFF_X1 \OUT1_reg[20]  ( .D(n5415), .CK(n79527), .Q(OUT1[20]) );
  DFF_X1 \OUT1_reg[19]  ( .D(n5413), .CK(n79527), .Q(OUT1[19]) );
  DFF_X1 \OUT1_reg[18]  ( .D(n5411), .CK(n79527), .Q(OUT1[18]) );
  DFF_X1 \OUT1_reg[17]  ( .D(n5409), .CK(n79527), .Q(OUT1[17]) );
  DFF_X1 \OUT1_reg[16]  ( .D(n5407), .CK(n79527), .Q(OUT1[16]) );
  DFF_X1 \OUT1_reg[15]  ( .D(n5405), .CK(n79527), .Q(OUT1[15]) );
  DFF_X1 \OUT1_reg[14]  ( .D(n5403), .CK(n79527), .Q(OUT1[14]) );
  DFF_X1 \OUT1_reg[13]  ( .D(n5401), .CK(n79527), .Q(OUT1[13]) );
  DFF_X1 \OUT1_reg[12]  ( .D(n5399), .CK(n79527), .Q(OUT1[12]) );
  DFF_X1 \OUT1_reg[11]  ( .D(n5397), .CK(n79527), .Q(OUT1[11]) );
  DFF_X1 \OUT1_reg[10]  ( .D(n5395), .CK(n79527), .Q(OUT1[10]) );
  DFF_X1 \OUT1_reg[9]  ( .D(n5393), .CK(n79527), .Q(OUT1[9]) );
  DFF_X1 \OUT1_reg[8]  ( .D(n5391), .CK(n79527), .Q(OUT1[8]) );
  DFF_X1 \OUT1_reg[7]  ( .D(n5389), .CK(n79527), .Q(OUT1[7]) );
  DFF_X1 \OUT1_reg[6]  ( .D(n5387), .CK(n79527), .Q(OUT1[6]) );
  DFF_X1 \OUT1_reg[5]  ( .D(n5385), .CK(n79527), .Q(OUT1[5]) );
  DFF_X1 \OUT1_reg[4]  ( .D(n5383), .CK(n79527), .Q(OUT1[4]) );
  DFF_X1 \OUT2_reg[6]  ( .D(n5317), .CK(n79527), .Q(OUT2[6]) );
  DFF_X1 \OUT2_reg[5]  ( .D(n5316), .CK(n79527), .Q(OUT2[5]) );
  DFF_X1 \OUT2_reg[4]  ( .D(n5315), .CK(n79527), .Q(OUT2[4]) );
  DFF_X1 \OUT2_reg[3]  ( .D(n5314), .CK(n79527), .Q(OUT2[3]) );
  DFF_X1 \OUT2_reg[2]  ( .D(n5313), .CK(n79527), .Q(OUT2[2]) );
  DFF_X1 \OUT2_reg[1]  ( .D(n5312), .CK(n79527), .Q(OUT2[1]) );
  DFF_X1 \OUT2_reg[0]  ( .D(n5311), .CK(n79527), .Q(OUT2[0]) );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n6970), .CK(n79527), .Q(n118718), .QN(
        n90036) );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n6969), .CK(n79527), .Q(n118717), .QN(
        n90037) );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n6968), .CK(n79527), .Q(n118716), .QN(
        n90038) );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n6967), .CK(n79527), .Q(n118715), .QN(
        n90039) );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n6966), .CK(n79527), .Q(n118714), .QN(
        n90040) );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n6965), .CK(n79527), .Q(n118713), .QN(
        n90041) );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n6964), .CK(n79527), .Q(n118712), .QN(
        n90042) );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n6963), .CK(n79527), .Q(n118711), .QN(
        n90043) );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n6962), .CK(n79527), .Q(n118710), .QN(
        n90044) );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n6961), .CK(n79527), .Q(n118709), .QN(
        n90045) );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n6960), .CK(n79527), .Q(n118708), .QN(
        n90046) );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n6959), .CK(n79527), .Q(n118707), .QN(
        n90047) );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n6958), .CK(n79527), .Q(n118706), .QN(
        n90048) );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n6957), .CK(n79527), .Q(n118705), .QN(
        n90049) );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n6956), .CK(n79527), .Q(n118704), .QN(
        n90050) );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n6955), .CK(n79527), .Q(n118703), .QN(
        n90051) );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n6954), .CK(n79527), .Q(n118702), .QN(
        n90052) );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n6953), .CK(n79527), .Q(n118701), .QN(
        n90053) );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n6952), .CK(n79527), .Q(n118700), .QN(
        n90054) );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n6951), .CK(n79527), .Q(n118699), .QN(
        n90055) );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n6950), .CK(n79527), .Q(n118698), .QN(
        n90056) );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n6949), .CK(n79527), .Q(n118697), .QN(
        n90057) );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n6948), .CK(n79527), .Q(n118696), .QN(
        n90058) );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n6947), .CK(n79527), .Q(n118695), .QN(
        n90059) );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n6946), .CK(n79527), .Q(n118694), .QN(
        n90060) );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n6945), .CK(n79527), .Q(n118693), .QN(
        n90061) );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n6944), .CK(n79527), .Q(n118692), .QN(
        n90062) );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n6943), .CK(n79527), .Q(n118691), .QN(
        n90063) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n6942), .CK(n79527), .Q(n118690), .QN(
        n90064) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n6941), .CK(n79527), .Q(n118689), .QN(
        n90065) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n6940), .CK(n79527), .Q(n118688), .QN(
        n90066) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n6939), .CK(n79527), .Q(n118687), .QN(
        n90067) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n6938), .CK(n79527), .Q(n118686), .QN(
        n90068) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n6937), .CK(n79527), .Q(n118685), .QN(
        n90069) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n6936), .CK(n79527), .Q(n118684), .QN(
        n90070) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n6935), .CK(n79527), .Q(n118683), .QN(
        n90071) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n6934), .CK(n79527), .Q(n118682), .QN(
        n90072) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n6933), .CK(n79527), .Q(n118681), .QN(
        n90073) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n6932), .CK(n79527), .Q(n118680), .QN(
        n90074) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n6931), .CK(n79527), .Q(n118679), .QN(
        n90075) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n6930), .CK(n79527), .Q(n118678), .QN(
        n90076) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n6929), .CK(n79527), .Q(n118677), .QN(
        n90077) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n6928), .CK(n79527), .Q(n118676), .QN(
        n90078) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n6927), .CK(n79527), .Q(n118675), .QN(
        n90079) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n6926), .CK(n79527), .Q(n118674), .QN(
        n90080) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n6925), .CK(n79527), .Q(n118673), .QN(
        n90081) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n6924), .CK(n79527), .Q(n118672), .QN(
        n90082) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n6923), .CK(n79527), .Q(n118671), .QN(
        n90083) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n6922), .CK(n79527), .Q(n118670), .QN(
        n90084) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n6921), .CK(n79527), .Q(n118730), .QN(
        n90085) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n6920), .CK(n79527), .Q(n118729), .QN(
        n90086) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n6919), .CK(n79527), .Q(n118728), .QN(
        n90087) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n6918), .CK(n79527), .Q(n118727), .QN(
        n90088) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n6917), .CK(n79527), .Q(n118737), .QN(
        n90089) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n6916), .CK(n79527), .Q(n118736), .QN(
        n90090) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n6915), .CK(n79527), .Q(n118735), .QN(
        n90091) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n6914), .CK(n79527), .Q(n118734), .QN(
        n90092) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n6913), .CK(n79527), .Q(n118733), .QN(
        n90093) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n6912), .CK(n79527), .Q(n118732), .QN(
        n90094) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n6911), .CK(n79527), .Q(n118731), .QN(
        n90095) );
  DFF_X1 \OUT2_reg[10]  ( .D(n5321), .CK(n79527), .Q(OUT2[10]) );
  DFF_X1 \OUT2_reg[9]  ( .D(n5320), .CK(n79527), .Q(OUT2[9]) );
  DFF_X1 \OUT2_reg[8]  ( .D(n5319), .CK(n79527), .Q(OUT2[8]) );
  DFF_X1 \OUT2_reg[7]  ( .D(n5318), .CK(n79527), .Q(OUT2[7]) );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n6014), .CK(n79527), .Q(n118985), .QN(
        n90711) );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n6013), .CK(n79527), .Q(n118984), .QN(
        n90713) );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n6012), .CK(n79527), .Q(n118983), .QN(
        n90714) );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n6011), .CK(n79527), .Q(n118982), .QN(
        n90715) );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n6398), .CK(n79527), .Q(n118549), .QN(
        n90373) );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n6397), .CK(n79527), .Q(n118548), .QN(
        n90375) );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n6396), .CK(n79527), .Q(n118547), .QN(
        n90376) );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n6395), .CK(n79527), .Q(n118546), .QN(
        n90377) );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n6462), .CK(n79527), .Q(n110482), .QN(
        n90306) );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n6461), .CK(n79527), .Q(n110481), .QN(
        n90308) );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n6460), .CK(n79527), .Q(n110480), .QN(
        n90309) );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n6459), .CK(n79527), .Q(n110479), .QN(
        n90310) );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n6206), .CK(n79527), .Q(n118861), .QN(
        n90512) );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n6205), .CK(n79527), .Q(n118860), .QN(
        n90514) );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n6204), .CK(n79527), .Q(n118859), .QN(
        n90515) );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n6203), .CK(n79527), .Q(n118858), .QN(
        n90516) );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n7486), .CK(n79527), .Q(n110110), .QN(
        n89493) );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n7485), .CK(n79527), .Q(n110109), .QN(
        n89496) );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n7484), .CK(n79527), .Q(n110108), .QN(
        n89498) );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n7483), .CK(n79527), .Q(n110107), .QN(
        n89500) );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n7038), .CK(n79527), .Q(n110366), .QN(
        n89965) );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n7037), .CK(n79527), .Q(n110365), .QN(
        n89967) );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n7036), .CK(n79527), .Q(n110364), .QN(
        n89968) );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n7035), .CK(n79527), .Q(n110363), .QN(
        n89969) );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n6974), .CK(n79527), .Q(n118726), .QN(
        n90031) );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n6973), .CK(n79527), .Q(n118725), .QN(
        n90033) );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n6972), .CK(n79527), .Q(n118724), .QN(
        n90034) );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n6971), .CK(n79527), .Q(n118723), .QN(
        n90035) );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n6010), .CK(n79527), .Q(n118999), .QN(
        n90716) );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n6009), .CK(n79527), .Q(n118998), .QN(
        n90717) );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n6008), .CK(n79527), .Q(n118997), .QN(
        n90718) );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n6007), .CK(n79527), .Q(n118996), .QN(
        n90719) );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n6006), .CK(n79527), .Q(n118995), .QN(
        n90720) );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n6005), .CK(n79527), .Q(n118994), .QN(
        n90721) );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n6004), .CK(n79527), .Q(n118993), .QN(
        n90722) );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n6003), .CK(n79527), .Q(n118992), .QN(
        n90723) );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n6002), .CK(n79527), .Q(n118991), .QN(
        n90724) );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n6001), .CK(n79527), .Q(n118990), .QN(
        n90725) );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n6000), .CK(n79527), .Q(n118989), .QN(
        n90726) );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n5999), .CK(n79527), .Q(n118988), .QN(
        n90727) );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n5998), .CK(n79527), .Q(n118987), .QN(
        n90728) );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n5997), .CK(n79527), .Q(n118986), .QN(
        n90729) );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n5996), .CK(n79527), .Q(n119045), .QN(
        n90730) );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n5995), .CK(n79527), .Q(n119044), .QN(
        n90731) );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n5994), .CK(n79527), .Q(n119043), .QN(
        n90732) );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n5993), .CK(n79527), .Q(n119042), .QN(
        n90733) );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n5992), .CK(n79527), .Q(n119041), .QN(
        n90734) );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n5991), .CK(n79527), .Q(n119040), .QN(
        n90735) );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n5990), .CK(n79527), .Q(n119039), .QN(
        n90736) );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n5989), .CK(n79527), .Q(n119038), .QN(
        n90737) );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n5988), .CK(n79527), .Q(n119037), .QN(
        n90738) );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n5987), .CK(n79527), .Q(n119036), .QN(
        n90739) );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n5986), .CK(n79527), .Q(n119035), .QN(
        n90740) );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n5985), .CK(n79527), .Q(n119034), .QN(
        n90741) );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n5984), .CK(n79527), .Q(n119033), .QN(
        n90742) );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n5983), .CK(n79527), .Q(n119032), .QN(
        n90743) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n5982), .CK(n79527), .Q(n119031), .QN(
        n90744) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5981), .CK(n79527), .Q(n119030), .QN(
        n90745) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5980), .CK(n79527), .Q(n119029), .QN(
        n90746) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5979), .CK(n79527), .Q(n119028), .QN(
        n90747) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n5978), .CK(n79527), .Q(n119027), .QN(
        n90748) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n5977), .CK(n79527), .Q(n119026), .QN(
        n90749) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n5976), .CK(n79527), .Q(n119025), .QN(
        n90750) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n5975), .CK(n79527), .Q(n119024), .QN(
        n90751) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n5974), .CK(n79527), .Q(n119023), .QN(
        n90752) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n5973), .CK(n79527), .Q(n119022), .QN(
        n90753) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n5972), .CK(n79527), .Q(n119021), .QN(
        n90754) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n5971), .CK(n79527), .Q(n119020), .QN(
        n90755) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n5970), .CK(n79527), .Q(n119019), .QN(
        n90756) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n5969), .CK(n79527), .Q(n119018), .QN(
        n90757) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n5968), .CK(n79527), .Q(n119017), .QN(
        n90758) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n5967), .CK(n79527), .Q(n119016), .QN(
        n90759) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n5966), .CK(n79527), .Q(n119015), .QN(
        n90760) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n5965), .CK(n79527), .Q(n119014), .QN(
        n90761) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n5964), .CK(n79527), .Q(n119013), .QN(
        n90762) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n5963), .CK(n79527), .Q(n119012), .QN(
        n90763) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n5962), .CK(n79527), .Q(n119011), .QN(
        n90764) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n5961), .CK(n79527), .Q(n119010), .QN(
        n90765) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n5960), .CK(n79527), .Q(n119009), .QN(
        n90766) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n5959), .CK(n79527), .Q(n119008), .QN(
        n90767) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n5958), .CK(n79527), .Q(n119007), .QN(
        n90768) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n5957), .CK(n79527), .Q(n119006), .QN(
        n90769) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n5956), .CK(n79527), .Q(n119005), .QN(
        n90770) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n5955), .CK(n79527), .Q(n119004), .QN(
        n90771) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n5954), .CK(n79527), .Q(n119003), .QN(
        n90772) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n5953), .CK(n79527), .Q(n119002), .QN(
        n90773) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n5952), .CK(n79527), .Q(n119001), .QN(
        n90774) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n5951), .CK(n79527), .Q(n119000), .QN(
        n90775) );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n6394), .CK(n79527), .Q(n118563), .QN(
        n90378) );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n6393), .CK(n79527), .Q(n118562), .QN(
        n90379) );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n6392), .CK(n79527), .Q(n118561), .QN(
        n90380) );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n6391), .CK(n79527), .Q(n118560), .QN(
        n90381) );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n6390), .CK(n79527), .Q(n118559), .QN(
        n90382) );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n6389), .CK(n79527), .Q(n118558), .QN(
        n90383) );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n6388), .CK(n79527), .Q(n118557), .QN(
        n90384) );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n6387), .CK(n79527), .Q(n118556), .QN(
        n90385) );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n6386), .CK(n79527), .Q(n118555), .QN(
        n90386) );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n6385), .CK(n79527), .Q(n118554), .QN(
        n90387) );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n6384), .CK(n79527), .Q(n118553), .QN(
        n90388) );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n6383), .CK(n79527), .Q(n118552), .QN(
        n90389) );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n6382), .CK(n79527), .Q(n118551), .QN(
        n90390) );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n6381), .CK(n79527), .Q(n118550), .QN(
        n90391) );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n6380), .CK(n79527), .Q(n118609), .QN(
        n90392) );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n6379), .CK(n79527), .Q(n118608), .QN(
        n90393) );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n6378), .CK(n79527), .Q(n118607), .QN(
        n90394) );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n6377), .CK(n79527), .Q(n118606), .QN(
        n90395) );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n6376), .CK(n79527), .Q(n118605), .QN(
        n90396) );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n6375), .CK(n79527), .Q(n118604), .QN(
        n90397) );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n6374), .CK(n79527), .Q(n118603), .QN(
        n90398) );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n6373), .CK(n79527), .Q(n118602), .QN(
        n90399) );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n6372), .CK(n79527), .Q(n118601), .QN(
        n90400) );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n6371), .CK(n79527), .Q(n118600), .QN(
        n90401) );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n6370), .CK(n79527), .Q(n118599), .QN(
        n90402) );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n6369), .CK(n79527), .Q(n118598), .QN(
        n90403) );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n6368), .CK(n79527), .Q(n118597), .QN(
        n90404) );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n6367), .CK(n79527), .Q(n118596), .QN(
        n90405) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n6366), .CK(n79527), .Q(n118595), .QN(
        n90406) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n6365), .CK(n79527), .Q(n118594), .QN(
        n90407) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n6364), .CK(n79527), .Q(n118593), .QN(
        n90408) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n6363), .CK(n79527), .Q(n118592), .QN(
        n90409) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n6362), .CK(n79527), .Q(n118591), .QN(
        n90410) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n6361), .CK(n79527), .Q(n118590), .QN(
        n90411) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n6360), .CK(n79527), .Q(n118589), .QN(
        n90412) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n6359), .CK(n79527), .Q(n118588), .QN(
        n90413) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n6358), .CK(n79527), .Q(n118587), .QN(
        n90414) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n6357), .CK(n79527), .Q(n118586), .QN(
        n90415) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n6356), .CK(n79527), .Q(n118585), .QN(
        n90416) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n6355), .CK(n79527), .Q(n118584), .QN(
        n90417) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n6354), .CK(n79527), .Q(n118583), .QN(
        n90418) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n6353), .CK(n79527), .Q(n118582), .QN(
        n90419) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n6352), .CK(n79527), .Q(n118581), .QN(
        n90420) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n6351), .CK(n79527), .Q(n118580), .QN(
        n90421) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n6350), .CK(n79527), .Q(n118579), .QN(
        n90422) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n6349), .CK(n79527), .Q(n118578), .QN(
        n90423) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n6348), .CK(n79527), .Q(n118577), .QN(
        n90424) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n6347), .CK(n79527), .Q(n118576), .QN(
        n90425) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n6346), .CK(n79527), .Q(n118575), .QN(
        n90426) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n6345), .CK(n79527), .Q(n118574), .QN(
        n90427) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n6344), .CK(n79527), .Q(n118573), .QN(
        n90428) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n6343), .CK(n79527), .Q(n118572), .QN(
        n90429) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n6342), .CK(n79527), .Q(n118571), .QN(
        n90430) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n6341), .CK(n79527), .Q(n118570), .QN(
        n90431) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n6340), .CK(n79527), .Q(n118569), .QN(
        n90432) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n6339), .CK(n79527), .Q(n118568), .QN(
        n90433) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n6338), .CK(n79527), .Q(n118567), .QN(
        n90434) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n6337), .CK(n79527), .Q(n118566), .QN(
        n90435) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n6336), .CK(n79527), .Q(n118565), .QN(
        n90436) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n6335), .CK(n79527), .Q(n118564), .QN(
        n90437) );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n6458), .CK(n79527), .Q(n110478), .QN(
        n90311) );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n6457), .CK(n79527), .Q(n110477), .QN(
        n90312) );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n6456), .CK(n79527), .Q(n110476), .QN(
        n90313) );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n6455), .CK(n79527), .Q(n110475), .QN(
        n90314) );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n6454), .CK(n79527), .Q(n110474), .QN(
        n90315) );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n6453), .CK(n79527), .Q(n110473), .QN(
        n90316) );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n6452), .CK(n79527), .Q(n110472), .QN(
        n90317) );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n6451), .CK(n79527), .Q(n110471), .QN(
        n90318) );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n6450), .CK(n79527), .Q(n110470), .QN(
        n90319) );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n6449), .CK(n79527), .Q(n110469), .QN(
        n90320) );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n6448), .CK(n79527), .Q(n110468), .QN(
        n90321) );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n6447), .CK(n79527), .Q(n110467), .QN(
        n90322) );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n6446), .CK(n79527), .Q(n110466), .QN(
        n90323) );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n6445), .CK(n79527), .Q(n110465), .QN(
        n90324) );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n6444), .CK(n79527), .Q(n110464), .QN(
        n90325) );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n6443), .CK(n79527), .Q(n110463), .QN(
        n90326) );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n6442), .CK(n79527), .Q(n110462), .QN(
        n90327) );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n6441), .CK(n79527), .Q(n110461), .QN(
        n90328) );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n6440), .CK(n79527), .Q(n110460), .QN(
        n90329) );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n6439), .CK(n79527), .Q(n110459), .QN(
        n90330) );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n6438), .CK(n79527), .Q(n110458), .QN(
        n90331) );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n6437), .CK(n79527), .Q(n110457), .QN(
        n90332) );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n6436), .CK(n79527), .Q(n110456), .QN(
        n90333) );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n6435), .CK(n79527), .Q(n110455), .QN(
        n90334) );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n6434), .CK(n79527), .Q(n110454), .QN(
        n90335) );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n6433), .CK(n79527), .Q(n110453), .QN(
        n90336) );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n6432), .CK(n79527), .Q(n110452), .QN(
        n90337) );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n6431), .CK(n79527), .Q(n110451), .QN(
        n90338) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n6430), .CK(n79527), .Q(n110450), .QN(
        n90339) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n6429), .CK(n79527), .Q(n110449), .QN(
        n90340) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n6428), .CK(n79527), .Q(n110448), .QN(
        n90341) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n6427), .CK(n79527), .Q(n110447), .QN(
        n90342) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n6426), .CK(n79527), .Q(n110446), .QN(
        n90343) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n6425), .CK(n79527), .Q(n110445), .QN(
        n90344) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n6424), .CK(n79527), .Q(n110444), .QN(
        n90345) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n6423), .CK(n79527), .Q(n110443), .QN(
        n90346) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n6422), .CK(n79527), .Q(n110442), .QN(
        n90347) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n6421), .CK(n79527), .Q(n110441), .QN(
        n90348) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n6420), .CK(n79527), .Q(n110440), .QN(
        n90349) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n6419), .CK(n79527), .Q(n110439), .QN(
        n90350) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n6418), .CK(n79527), .Q(n110438), .QN(
        n90351) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n6417), .CK(n79527), .Q(n110437), .QN(
        n90352) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n6416), .CK(n79527), .Q(n110436), .QN(
        n90353) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n6415), .CK(n79527), .Q(n110435), .QN(
        n90354) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n6414), .CK(n79527), .Q(n110434), .QN(
        n90355) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n6413), .CK(n79527), .Q(n110433), .QN(
        n90356) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n6412), .CK(n79527), .Q(n110432), .QN(
        n90357) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n6411), .CK(n79527), .Q(n110431), .QN(
        n90358) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n6410), .CK(n79527), .Q(n110491), .QN(
        n90359) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n6409), .CK(n79527), .Q(n110490), .QN(
        n90360) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n6408), .CK(n79527), .Q(n110489), .QN(
        n90361) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n6407), .CK(n79527), .Q(n110488), .QN(
        n90362) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n6406), .CK(n79527), .Q(n110487), .QN(
        n90363) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n6405), .CK(n79527), .Q(n110546), .QN(
        n90364) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n6404), .CK(n79527), .Q(n110545), .QN(
        n90365) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n6403), .CK(n79527), .Q(n110544), .QN(
        n90366) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n6402), .CK(n79527), .Q(n110543), .QN(
        n90367) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n6401), .CK(n79527), .Q(n110542), .QN(
        n90368) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n6400), .CK(n79527), .Q(n110541), .QN(
        n90369) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n6399), .CK(n79527), .Q(n110540), .QN(
        n90370) );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n6202), .CK(n79527), .Q(n118857), .QN(
        n90517) );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n6201), .CK(n79527), .Q(n118856), .QN(
        n90518) );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n6200), .CK(n79527), .Q(n118855), .QN(
        n90519) );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n6199), .CK(n79527), .Q(n118854), .QN(
        n90520) );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n6198), .CK(n79527), .Q(n118853), .QN(
        n90521) );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n6197), .CK(n79527), .Q(n118852), .QN(
        n90522) );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n6196), .CK(n79527), .Q(n118851), .QN(
        n90523) );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n6195), .CK(n79527), .Q(n118850), .QN(
        n90524) );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n6194), .CK(n79527), .Q(n118849), .QN(
        n90525) );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n6193), .CK(n79527), .Q(n118848), .QN(
        n90526) );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n6192), .CK(n79527), .Q(n118847), .QN(
        n90527) );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n6191), .CK(n79527), .Q(n118846), .QN(
        n90528) );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n6190), .CK(n79527), .Q(n118845), .QN(
        n90529) );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n6189), .CK(n79527), .Q(n118844), .QN(
        n90530) );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n6188), .CK(n79527), .Q(n118843), .QN(
        n90531) );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n6187), .CK(n79527), .Q(n118842), .QN(
        n90532) );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n6186), .CK(n79527), .Q(n118841), .QN(
        n90533) );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n6185), .CK(n79527), .Q(n118840), .QN(
        n90534) );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n6184), .CK(n79527), .Q(n118839), .QN(
        n90535) );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n6183), .CK(n79527), .Q(n118838), .QN(
        n90536) );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n6182), .CK(n79527), .Q(n118837), .QN(
        n90537) );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n6181), .CK(n79527), .Q(n118836), .QN(
        n90538) );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n6180), .CK(n79527), .Q(n118835), .QN(
        n90539) );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n6179), .CK(n79527), .Q(n118834), .QN(
        n90540) );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n6178), .CK(n79527), .Q(n118833), .QN(
        n90541) );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n6177), .CK(n79527), .Q(n118832), .QN(
        n90542) );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n6176), .CK(n79527), .Q(n118831), .QN(
        n90543) );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n6175), .CK(n79527), .Q(n118830), .QN(
        n90544) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n6174), .CK(n79527), .Q(n118829), .QN(
        n90545) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n6173), .CK(n79527), .Q(n118828), .QN(
        n90546) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n6172), .CK(n79527), .Q(n118827), .QN(
        n90547) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n6171), .CK(n79527), .Q(n118826), .QN(
        n90548) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n6170), .CK(n79527), .Q(n118825), .QN(
        n90549) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n6169), .CK(n79527), .Q(n118824), .QN(
        n90550) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n6168), .CK(n79527), .Q(n118823), .QN(
        n90551) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n6167), .CK(n79527), .Q(n118822), .QN(
        n90552) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n6166), .CK(n79527), .Q(n118821), .QN(
        n90553) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n6165), .CK(n79527), .Q(n118820), .QN(
        n90554) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n6164), .CK(n79527), .Q(n118819), .QN(
        n90555) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n6163), .CK(n79527), .Q(n118818), .QN(
        n90556) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n6162), .CK(n79527), .Q(n118817), .QN(
        n90557) );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n5630), .CK(n79527), .Q(n110874), .QN(
        n99914) );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n5629), .CK(n79527), .Q(n110873), .QN(
        n99916) );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n5628), .CK(n79527), .Q(n110872), .QN(
        n99917) );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n5627), .CK(n79527), .Q(n110871), .QN(
        n99918) );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n5886), .CK(n79527), .Q(n119049), .QN(
        n99716) );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n5885), .CK(n79527), .Q(n119048), .QN(
        n99718) );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n5884), .CK(n79527), .Q(n119047), .QN(
        n99719) );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n5883), .CK(n79527), .Q(n119046), .QN(
        n99720) );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n6270), .CK(n79527), .Q(n118722), .QN(
        n99446) );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n6269), .CK(n79527), .Q(n118721), .QN(
        n99448) );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n6268), .CK(n79527), .Q(n118720), .QN(
        n99449) );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n6267), .CK(n79527), .Q(n118719), .QN(
        n99450) );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n6078), .CK(n79527), .QN(n99580) );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n6077), .CK(n79527), .QN(n99582) );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n6076), .CK(n79527), .QN(n99583) );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n6075), .CK(n79527), .QN(n99584) );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n7294), .CK(n79527), .Q(n110192), .QN(
        n98648) );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n7293), .CK(n79527), .Q(n110191), .QN(
        n98650) );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n7292), .CK(n79527), .Q(n110190), .QN(
        n98651) );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n7291), .CK(n79527), .Q(n110189), .QN(
        n98652) );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n7230), .CK(n79527), .Q(n110486), .QN(
        n98714) );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n7229), .CK(n79527), .Q(n110485), .QN(
        n98716) );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n7228), .CK(n79527), .Q(n110484), .QN(
        n98717) );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n7227), .CK(n79527), .Q(n110483), .QN(
        n98718) );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n6590), .CK(n79527), .Q(n119177), .QN(
        n99245) );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n6589), .CK(n79527), .Q(n119176), .QN(
        n99247) );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n6588), .CK(n79527), .Q(n119175), .QN(
        n99248) );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n6587), .CK(n79527), .Q(n119174), .QN(
        n99249) );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n6718), .CK(n79527), .Q(n119354), .QN(
        n99113) );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n6717), .CK(n79527), .Q(n119353), .QN(
        n99115) );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n6716), .CK(n79527), .Q(n119352), .QN(
        n99116) );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n6715), .CK(n79527), .Q(n119351), .QN(
        n99117) );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n5626), .CK(n79527), .Q(n110863), .QN(
        n99919) );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n5625), .CK(n79527), .Q(n110862), .QN(
        n99920) );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n5624), .CK(n79527), .Q(n110861), .QN(
        n99921) );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n5623), .CK(n79527), .Q(n110860), .QN(
        n99922) );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n5622), .CK(n79527), .Q(n110859), .QN(
        n99923) );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n5621), .CK(n79527), .Q(n110858), .QN(
        n99924) );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n5620), .CK(n79527), .Q(n110857), .QN(
        n99925) );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n5619), .CK(n79527), .Q(n110856), .QN(
        n99926) );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n5618), .CK(n79527), .Q(n110855), .QN(
        n99927) );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n5617), .CK(n79527), .Q(n110854), .QN(
        n99928) );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n5616), .CK(n79527), .Q(n110853), .QN(
        n99929) );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n5615), .CK(n79527), .Q(n110852), .QN(
        n99930) );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n5614), .CK(n79527), .Q(n110851), .QN(
        n99931) );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n5613), .CK(n79527), .Q(n110850), .QN(
        n99932) );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n5612), .CK(n79527), .Q(n110849), .QN(
        n99933) );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n5611), .CK(n79527), .Q(n110848), .QN(
        n99934) );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n5610), .CK(n79527), .Q(n110847), .QN(
        n99935) );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n5609), .CK(n79527), .Q(n110846), .QN(
        n99936) );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n5608), .CK(n79527), .Q(n110845), .QN(
        n99937) );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n5607), .CK(n79527), .Q(n110844), .QN(
        n99938) );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n5606), .CK(n79527), .Q(n110843), .QN(
        n99939) );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n5605), .CK(n79527), .Q(n110842), .QN(
        n99940) );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n5604), .CK(n79527), .Q(n110841), .QN(
        n99941) );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n5603), .CK(n79527), .Q(n110840), .QN(
        n99942) );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n5602), .CK(n79527), .Q(n110839), .QN(
        n99943) );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n5601), .CK(n79527), .Q(n110838), .QN(
        n99944) );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n5600), .CK(n79527), .Q(n110837), .QN(
        n99945) );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n5599), .CK(n79527), .Q(n110836), .QN(
        n99946) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n5598), .CK(n79527), .Q(n110835), .QN(
        n99947) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5597), .CK(n79527), .Q(n110834), .QN(
        n99948) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5596), .CK(n79527), .Q(n110833), .QN(
        n99949) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5595), .CK(n79527), .Q(n110832), .QN(
        n99950) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n5594), .CK(n79527), .Q(n110831), .QN(
        n99951) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n5593), .CK(n79527), .Q(n110830), .QN(
        n99952) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n5592), .CK(n79527), .Q(n110829), .QN(
        n99953) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n5591), .CK(n79527), .Q(n110828), .QN(
        n99954) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n5590), .CK(n79527), .Q(n110827), .QN(
        n99955) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n5589), .CK(n79527), .Q(n110826), .QN(
        n99956) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n5588), .CK(n79527), .Q(n110825), .QN(
        n99957) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n5587), .CK(n79527), .Q(n110824), .QN(
        n99958) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n5586), .CK(n79527), .Q(n110823), .QN(
        n99959) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n5585), .CK(n79527), .Q(n110822), .QN(
        n99960) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n5584), .CK(n79527), .Q(n110821), .QN(
        n99961) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n5583), .CK(n79527), .Q(n110820), .QN(
        n99962) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n5582), .CK(n79527), .Q(n110819), .QN(
        n99963) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n5581), .CK(n79527), .Q(n110818), .QN(
        n99964) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n5580), .CK(n79527), .Q(n110817), .QN(
        n99965) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n5579), .CK(n79527), .Q(n110816), .QN(
        n99966) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n5578), .CK(n79527), .Q(n110815), .QN(
        n99967) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n5577), .CK(n79527), .Q(n110814), .QN(
        n99968) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n5576), .CK(n79527), .Q(n110813), .QN(
        n99969) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n5575), .CK(n79527), .Q(n110812), .QN(
        n99970) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n5574), .CK(n79527), .Q(n110811), .QN(
        n99971) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n5573), .CK(n79527), .Q(n110870), .QN(
        n99972) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n5572), .CK(n79527), .Q(n110869), .QN(
        n99973) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n5571), .CK(n79527), .Q(n110868), .QN(
        n99974) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n5570), .CK(n79527), .Q(n110867), .QN(
        n99975) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n5569), .CK(n79527), .Q(n110866), .QN(
        n99976) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n5568), .CK(n79527), .Q(n110865), .QN(
        n99977) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n5567), .CK(n79527), .Q(n110864), .QN(
        n99978) );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n5882), .CK(n79527), .Q(n119063), .QN(
        n99721) );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n5881), .CK(n79527), .Q(n119062), .QN(
        n99722) );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n5880), .CK(n79527), .Q(n119061), .QN(
        n99723) );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n5879), .CK(n79527), .Q(n119060), .QN(
        n99724) );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n5878), .CK(n79527), .Q(n119059), .QN(
        n99725) );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n5877), .CK(n79527), .Q(n119058), .QN(
        n99726) );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n5876), .CK(n79527), .Q(n119057), .QN(
        n99727) );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n5875), .CK(n79527), .Q(n119056), .QN(
        n99728) );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n5874), .CK(n79527), .Q(n119055), .QN(
        n99729) );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n5873), .CK(n79527), .Q(n119054), .QN(
        n99730) );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n5872), .CK(n79527), .Q(n119053), .QN(
        n99731) );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n5871), .CK(n79527), .Q(n119052), .QN(
        n99732) );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n5870), .CK(n79527), .Q(n119051), .QN(
        n99733) );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n5869), .CK(n79527), .Q(n119050), .QN(
        n99734) );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n5868), .CK(n79527), .Q(n119109), .QN(
        n99735) );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n5867), .CK(n79527), .Q(n119108), .QN(
        n99736) );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n5866), .CK(n79527), .Q(n119107), .QN(
        n99737) );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n5865), .CK(n79527), .Q(n119106), .QN(
        n99738) );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n5864), .CK(n79527), .Q(n119105), .QN(
        n99739) );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n5863), .CK(n79527), .Q(n119104), .QN(
        n99740) );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n5862), .CK(n79527), .Q(n119103), .QN(
        n99741) );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n5861), .CK(n79527), .Q(n119102), .QN(
        n99742) );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n5860), .CK(n79527), .Q(n119101), .QN(
        n99743) );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n5859), .CK(n79527), .Q(n119100), .QN(
        n99744) );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n5858), .CK(n79527), .Q(n119099), .QN(
        n99745) );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n5857), .CK(n79527), .Q(n119098), .QN(
        n99746) );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n5856), .CK(n79527), .Q(n119097), .QN(
        n99747) );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n5855), .CK(n79527), .Q(n119096), .QN(
        n99748) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n5854), .CK(n79527), .Q(n119095), .QN(
        n99749) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5853), .CK(n79527), .Q(n119094), .QN(
        n99750) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5852), .CK(n79527), .Q(n119093), .QN(
        n99751) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5851), .CK(n79527), .Q(n119092), .QN(
        n99752) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n5850), .CK(n79527), .Q(n119091), .QN(
        n99753) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n5849), .CK(n79527), .Q(n119090), .QN(
        n99754) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n5848), .CK(n79527), .Q(n119089), .QN(
        n99755) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n5847), .CK(n79527), .Q(n119088), .QN(
        n99756) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n5846), .CK(n79527), .Q(n119087), .QN(
        n99757) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n5845), .CK(n79527), .Q(n119086), .QN(
        n99758) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n5844), .CK(n79527), .Q(n119085), .QN(
        n99759) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n5843), .CK(n79527), .Q(n119084), .QN(
        n99760) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n5842), .CK(n79527), .Q(n119083), .QN(
        n99761) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n5841), .CK(n79527), .Q(n119082), .QN(
        n99762) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n5840), .CK(n79527), .Q(n119081), .QN(
        n99763) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n5839), .CK(n79527), .Q(n119080), .QN(
        n99764) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n5838), .CK(n79527), .Q(n119079), .QN(
        n99765) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n5837), .CK(n79527), .Q(n119078), .QN(
        n99766) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n5836), .CK(n79527), .Q(n119077), .QN(
        n99767) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n5835), .CK(n79527), .Q(n119076), .QN(
        n99768) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n5834), .CK(n79527), .Q(n119075), .QN(
        n99769) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n5833), .CK(n79527), .Q(n119074), .QN(
        n99770) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n5832), .CK(n79527), .Q(n119073), .QN(
        n99771) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n5831), .CK(n79527), .Q(n119072), .QN(
        n99772) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n5830), .CK(n79527), .Q(n119071), .QN(
        n99773) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n5829), .CK(n79527), .Q(n119070), .QN(
        n99774) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n5828), .CK(n79527), .Q(n119069), .QN(
        n99775) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n5827), .CK(n79527), .Q(n119068), .QN(
        n99776) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n5826), .CK(n79527), .Q(n119067), .QN(
        n99777) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n5825), .CK(n79527), .Q(n119066), .QN(
        n99778) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n5824), .CK(n79527), .Q(n119065), .QN(
        n99779) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n5823), .CK(n79527), .Q(n119064), .QN(
        n99780) );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n6266), .CK(n79527), .Q(n118623), .QN(
        n99451) );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n6265), .CK(n79527), .Q(n118622), .QN(
        n99452) );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n6264), .CK(n79527), .Q(n118621), .QN(
        n99453) );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n6263), .CK(n79527), .Q(n118620), .QN(
        n99454) );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n6262), .CK(n79527), .Q(n118619), .QN(
        n99455) );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n6261), .CK(n79527), .Q(n118618), .QN(
        n99456) );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n6260), .CK(n79527), .Q(n118617), .QN(
        n99457) );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n6259), .CK(n79527), .Q(n118616), .QN(
        n99458) );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n6258), .CK(n79527), .Q(n118615), .QN(
        n99459) );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n6257), .CK(n79527), .Q(n118614), .QN(
        n99460) );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n6256), .CK(n79527), .Q(n118613), .QN(
        n99461) );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n6255), .CK(n79527), .Q(n118612), .QN(
        n99462) );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n6254), .CK(n79527), .Q(n118611), .QN(
        n99463) );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n6253), .CK(n79527), .Q(n118610), .QN(
        n99464) );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n6252), .CK(n79527), .Q(n118657), .QN(
        n99465) );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n6251), .CK(n79527), .Q(n118656), .QN(
        n99466) );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n6250), .CK(n79527), .Q(n118655), .QN(
        n99467) );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n6249), .CK(n79527), .Q(n118654), .QN(
        n99468) );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n6248), .CK(n79527), .Q(n118653), .QN(
        n99469) );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n6247), .CK(n79527), .Q(n118652), .QN(
        n99470) );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n6246), .CK(n79527), .Q(n118651), .QN(
        n99471) );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n6245), .CK(n79527), .Q(n118650), .QN(
        n99472) );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n6244), .CK(n79527), .Q(n118649), .QN(
        n99473) );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n6243), .CK(n79527), .Q(n118648), .QN(
        n99474) );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n6242), .CK(n79527), .Q(n118647), .QN(
        n99475) );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n6241), .CK(n79527), .Q(n118646), .QN(
        n99476) );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n6240), .CK(n79527), .Q(n118645), .QN(
        n99477) );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n6239), .CK(n79527), .Q(n118644), .QN(
        n99478) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n6238), .CK(n79527), .Q(n118643), .QN(
        n99479) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n6237), .CK(n79527), .Q(n118642), .QN(
        n99480) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n6236), .CK(n79527), .Q(n118641), .QN(
        n99481) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n6235), .CK(n79527), .Q(n118640), .QN(
        n99482) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n6234), .CK(n79527), .Q(n118639), .QN(
        n99483) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n6233), .CK(n79527), .Q(n118638), .QN(
        n99484) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n6232), .CK(n79527), .Q(n118637), .QN(
        n99485) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n6231), .CK(n79527), .Q(n118636), .QN(
        n99486) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n6230), .CK(n79527), .Q(n118635), .QN(
        n99487) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n6229), .CK(n79527), .Q(n118634), .QN(
        n99488) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n6228), .CK(n79527), .Q(n118633), .QN(
        n99489) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n6227), .CK(n79527), .Q(n118632), .QN(
        n99490) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n6226), .CK(n79527), .Q(n118631), .QN(
        n99491) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n6225), .CK(n79527), .Q(n118630), .QN(
        n99492) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n6224), .CK(n79527), .Q(n118629), .QN(
        n99493) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n6223), .CK(n79527), .Q(n118628), .QN(
        n99494) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n6222), .CK(n79527), .Q(n118627), .QN(
        n99495) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n6221), .CK(n79527), .Q(n118626), .QN(
        n99496) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n6220), .CK(n79527), .Q(n118625), .QN(
        n99497) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n6219), .CK(n79527), .Q(n118624), .QN(
        n99498) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n6218), .CK(n79527), .Q(n118669), .QN(
        n99499) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n6217), .CK(n79527), .Q(n118668), .QN(
        n99500) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n6216), .CK(n79527), .Q(n118667), .QN(
        n99501) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n6215), .CK(n79527), .Q(n118666), .QN(
        n99502) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n6214), .CK(n79527), .Q(n118665), .QN(
        n99503) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n6213), .CK(n79527), .Q(n118664), .QN(
        n99504) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n6212), .CK(n79527), .Q(n118663), .QN(
        n99505) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n6211), .CK(n79527), .Q(n118662), .QN(
        n99506) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n6210), .CK(n79527), .Q(n118661), .QN(
        n99507) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n6209), .CK(n79527), .Q(n118660), .QN(
        n99508) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n6208), .CK(n79527), .Q(n118659), .QN(
        n99509) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n6207), .CK(n79527), .Q(n118658), .QN(
        n99510) );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n6074), .CK(n79527), .QN(n99585) );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n6073), .CK(n79527), .QN(n99586) );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n6072), .CK(n79527), .QN(n99587) );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n6071), .CK(n79527), .QN(n99588) );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n6070), .CK(n79527), .QN(n99589) );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n6069), .CK(n79527), .QN(n99590) );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n6068), .CK(n79527), .QN(n99591) );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n6067), .CK(n79527), .QN(n99592) );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n6066), .CK(n79527), .QN(n99593) );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n6065), .CK(n79527), .QN(n99594) );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n6064), .CK(n79527), .QN(n99595) );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n6063), .CK(n79527), .QN(n99596) );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n6062), .CK(n79527), .QN(n99597) );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n6061), .CK(n79527), .QN(n99598) );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n6060), .CK(n79527), .QN(n99599) );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n6059), .CK(n79527), .QN(n99600) );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n6058), .CK(n79527), .QN(n99601) );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n6057), .CK(n79527), .QN(n99602) );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n6056), .CK(n79527), .QN(n99603) );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n6055), .CK(n79527), .QN(n99604) );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n6054), .CK(n79527), .QN(n99605) );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n6053), .CK(n79527), .QN(n99606) );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n6052), .CK(n79527), .QN(n99607) );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n6051), .CK(n79527), .QN(n99608) );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n6050), .CK(n79527), .QN(n99609) );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n6049), .CK(n79527), .QN(n99610) );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n6048), .CK(n79527), .QN(n99611) );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n6047), .CK(n79527), .QN(n99612) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n6046), .CK(n79527), .QN(n99613) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n6045), .CK(n79527), .QN(n99614) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n6044), .CK(n79527), .QN(n99615) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n6043), .CK(n79527), .QN(n99616) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n6042), .CK(n79527), .QN(n99617) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n6041), .CK(n79527), .QN(n99618) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n6040), .CK(n79527), .QN(n99619) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n6039), .CK(n79527), .QN(n99620) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n6038), .CK(n79527), .QN(n99621) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n6037), .CK(n79527), .QN(n99622) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n6036), .CK(n79527), .QN(n99623) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n6035), .CK(n79527), .QN(n99624) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n6034), .CK(n79527), .QN(n99625) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n6033), .CK(n79527), .QN(n99626) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n6032), .CK(n79527), .QN(n99627) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n6031), .CK(n79527), .QN(n99628) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n6030), .CK(n79527), .QN(n99629) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n6029), .CK(n79527), .QN(n99630) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n6028), .CK(n79527), .QN(n99631) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n6027), .CK(n79527), .QN(n99632) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n6026), .CK(n79527), .QN(n99633) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n6025), .CK(n79527), .QN(n99634) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n6024), .CK(n79527), .QN(n99635) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n6023), .CK(n79527), .QN(n99636) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n6022), .CK(n79527), .QN(n99637) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n6021), .CK(n79527), .QN(n99638) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n6020), .CK(n79527), .QN(n99639) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n6019), .CK(n79527), .QN(n99640) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n6018), .CK(n79527), .QN(n99641) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n6017), .CK(n79527), .QN(n99642) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n6016), .CK(n79527), .QN(n99643) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n6015), .CK(n79527), .QN(n99644) );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n6782), .CK(n79527), .Q(n110580), .QN(
        n99047) );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n6781), .CK(n79527), .Q(n110579), .QN(
        n99049) );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n6780), .CK(n79527), .Q(n110578), .QN(
        n99050) );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n6779), .CK(n79527), .Q(n110577), .QN(
        n99051) );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n6526), .CK(n79527), .Q(n119301), .QN(
        n99311) );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n6525), .CK(n79527), .Q(n119300), .QN(
        n99313) );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n6524), .CK(n79527), .Q(n119299), .QN(
        n99314) );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n6523), .CK(n79527), .Q(n119298), .QN(
        n99315) );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n6654), .CK(n79527), .Q(n119113), .QN(
        n99179) );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n6653), .CK(n79527), .Q(n119112), .QN(
        n99181) );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n6652), .CK(n79527), .Q(n119111), .QN(
        n99182) );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n6651), .CK(n79527), .Q(n119110), .QN(
        n99183) );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n7354), .CK(n79527), .Q(n118910), .QN(
        n98586) );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n7353), .CK(n79527), .Q(n118909), .QN(
        n98587) );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n7352), .CK(n79527), .Q(n118908), .QN(
        n98588) );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n7351), .CK(n79527), .Q(n118907), .QN(
        n98589) );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n7350), .CK(n79527), .Q(n118906), .QN(
        n98590) );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n7349), .CK(n79527), .Q(n118905), .QN(
        n98591) );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n7348), .CK(n79527), .Q(n118904), .QN(
        n98592) );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n7347), .CK(n79527), .Q(n118903), .QN(
        n98593) );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n7346), .CK(n79527), .Q(n118902), .QN(
        n98594) );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n7345), .CK(n79527), .Q(n118901), .QN(
        n98595) );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n7344), .CK(n79527), .Q(n118900), .QN(
        n98596) );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n7343), .CK(n79527), .Q(n118899), .QN(
        n98597) );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n7342), .CK(n79527), .Q(n118898), .QN(
        n98598) );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n7341), .CK(n79527), .Q(n118897), .QN(
        n98599) );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n7340), .CK(n79527), .Q(n118896), .QN(
        n98600) );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n7339), .CK(n79527), .Q(n118895), .QN(
        n98601) );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n7338), .CK(n79527), .Q(n118894), .QN(
        n98602) );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n7337), .CK(n79527), .Q(n118893), .QN(
        n98603) );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n7336), .CK(n79527), .Q(n118892), .QN(
        n98604) );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n7335), .CK(n79527), .Q(n118891), .QN(
        n98605) );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n7334), .CK(n79527), .Q(n118890), .QN(
        n98606) );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n7333), .CK(n79527), .Q(n118889), .QN(
        n98607) );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n7332), .CK(n79527), .Q(n118888), .QN(
        n98608) );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n7331), .CK(n79527), .Q(n118887), .QN(
        n98609) );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n7330), .CK(n79527), .Q(n118886), .QN(
        n98610) );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n7329), .CK(n79527), .Q(n118885), .QN(
        n98611) );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n7328), .CK(n79527), .Q(n118884), .QN(
        n98612) );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n7327), .CK(n79527), .Q(n118883), .QN(
        n98613) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n7326), .CK(n79527), .Q(n118882), .QN(
        n98614) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n7325), .CK(n79527), .Q(n118881), .QN(
        n98615) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n7324), .CK(n79527), .Q(n118880), .QN(
        n98616) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n7323), .CK(n79527), .Q(n118879), .QN(
        n98617) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n7322), .CK(n79527), .Q(n118878), .QN(
        n98618) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n7321), .CK(n79527), .Q(n118877), .QN(
        n98619) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n7320), .CK(n79527), .Q(n118876), .QN(
        n98620) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n7319), .CK(n79527), .Q(n118875), .QN(
        n98621) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n7318), .CK(n79527), .Q(n118874), .QN(
        n98622) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n7317), .CK(n79527), .Q(n118873), .QN(
        n98623) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n7316), .CK(n79527), .Q(n118872), .QN(
        n98624) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n7315), .CK(n79527), .Q(n118871), .QN(
        n98625) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n7314), .CK(n79527), .Q(n118870), .QN(
        n98626) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n7313), .CK(n79527), .Q(n118869), .QN(
        n98627) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n7312), .CK(n79527), .Q(n118868), .QN(
        n98628) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n7311), .CK(n79527), .Q(n118867), .QN(
        n98629) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n7310), .CK(n79527), .Q(n118866), .QN(
        n98630) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n7309), .CK(n79527), .Q(n118865), .QN(
        n98631) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n7308), .CK(n79527), .Q(n118864), .QN(
        n98632) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n7307), .CK(n79527), .Q(n118863), .QN(
        n98633) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n7306), .CK(n79527), .Q(n118862), .QN(
        n98634) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n7305), .CK(n79527), .Q(n118914), .QN(
        n98635) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n7304), .CK(n79527), .Q(n118913), .QN(
        n98636) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n7303), .CK(n79527), .Q(n118912), .QN(
        n98637) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n7302), .CK(n79527), .Q(n118911), .QN(
        n98638) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n7301), .CK(n79527), .Q(n118921), .QN(
        n98639) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n7300), .CK(n79527), .Q(n118920), .QN(
        n98640) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n7299), .CK(n79527), .Q(n118919), .QN(
        n98641) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n7298), .CK(n79527), .Q(n118918), .QN(
        n98642) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n7297), .CK(n79527), .Q(n118917), .QN(
        n98643) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n7296), .CK(n79527), .Q(n118916), .QN(
        n98644) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n7295), .CK(n79527), .Q(n118915), .QN(
        n98645) );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n7290), .CK(n79527), .Q(n110184), .QN(
        n98653) );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n7289), .CK(n79527), .Q(n110183), .QN(
        n98654) );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n7288), .CK(n79527), .Q(n110182), .QN(
        n98655) );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n7287), .CK(n79527), .Q(n110181), .QN(
        n98656) );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n7286), .CK(n79527), .Q(n110180), .QN(
        n98657) );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n7285), .CK(n79527), .Q(n110179), .QN(
        n98658) );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n7284), .CK(n79527), .Q(n110178), .QN(
        n98659) );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n7283), .CK(n79527), .Q(n110177), .QN(
        n98660) );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n7282), .CK(n79527), .Q(n110176), .QN(
        n98661) );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n7281), .CK(n79527), .Q(n110175), .QN(
        n98662) );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n7280), .CK(n79527), .Q(n110174), .QN(
        n98663) );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n7279), .CK(n79527), .Q(n110173), .QN(
        n98664) );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n7278), .CK(n79527), .Q(n110172), .QN(
        n98665) );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n7277), .CK(n79527), .Q(n110171), .QN(
        n98666) );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n7276), .CK(n79527), .Q(n110234), .QN(
        n98667) );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n7275), .CK(n79527), .Q(n110233), .QN(
        n98668) );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n7274), .CK(n79527), .Q(n110232), .QN(
        n98669) );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n7273), .CK(n79527), .Q(n110231), .QN(
        n98670) );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n7272), .CK(n79527), .Q(n110230), .QN(
        n98671) );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n7271), .CK(n79527), .Q(n110229), .QN(
        n98672) );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n7270), .CK(n79527), .Q(n110228), .QN(
        n98673) );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n7269), .CK(n79527), .Q(n110227), .QN(
        n98674) );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n7268), .CK(n79527), .Q(n110226), .QN(
        n98675) );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n7267), .CK(n79527), .Q(n110225), .QN(
        n98676) );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n7266), .CK(n79527), .Q(n110224), .QN(
        n98677) );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n7265), .CK(n79527), .Q(n110223), .QN(
        n98678) );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n7264), .CK(n79527), .Q(n110222), .QN(
        n98679) );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n7263), .CK(n79527), .Q(n110221), .QN(
        n98680) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n7262), .CK(n79527), .Q(n110220), .QN(
        n98681) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n7261), .CK(n79527), .Q(n110219), .QN(
        n98682) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n7260), .CK(n79527), .Q(n110218), .QN(
        n98683) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n7259), .CK(n79527), .Q(n110217), .QN(
        n98684) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n7258), .CK(n79527), .Q(n110216), .QN(
        n98685) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n7257), .CK(n79527), .Q(n110215), .QN(
        n98686) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n7256), .CK(n79527), .Q(n110214), .QN(
        n98687) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n7255), .CK(n79527), .Q(n110213), .QN(
        n98688) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n7254), .CK(n79527), .Q(n110212), .QN(
        n98689) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n7253), .CK(n79527), .Q(n110211), .QN(
        n98690) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n7252), .CK(n79527), .Q(n110210), .QN(
        n98691) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n7251), .CK(n79527), .Q(n110209), .QN(
        n98692) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n7250), .CK(n79527), .Q(n110208), .QN(
        n98693) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n7249), .CK(n79527), .Q(n110207), .QN(
        n98694) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n7248), .CK(n79527), .Q(n110206), .QN(
        n98695) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n7247), .CK(n79527), .Q(n110205), .QN(
        n98696) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n7246), .CK(n79527), .Q(n110204), .QN(
        n98697) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n7245), .CK(n79527), .Q(n110203), .QN(
        n98698) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n7244), .CK(n79527), .Q(n110202), .QN(
        n98699) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n7243), .CK(n79527), .Q(n110201), .QN(
        n98700) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n7242), .CK(n79527), .Q(n110200), .QN(
        n98701) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n7241), .CK(n79527), .Q(n110199), .QN(
        n98702) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n7240), .CK(n79527), .Q(n110198), .QN(
        n98703) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n7239), .CK(n79527), .Q(n110197), .QN(
        n98704) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n7238), .CK(n79527), .Q(n110196), .QN(
        n98705) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n7237), .CK(n79527), .Q(n110195), .QN(
        n98706) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n7236), .CK(n79527), .Q(n110194), .QN(
        n98707) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n7235), .CK(n79527), .Q(n110193), .QN(
        n98708) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n7234), .CK(n79527), .Q(n110188), .QN(
        n98709) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n7233), .CK(n79527), .Q(n110187), .QN(
        n98710) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n7232), .CK(n79527), .Q(n110186), .QN(
        n98711) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n7231), .CK(n79527), .Q(n110185), .QN(
        n98712) );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n7418), .CK(n79527), .Q(n118545), .QN(
        n98523) );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n7417), .CK(n79527), .Q(n118544), .QN(
        n98524) );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n7416), .CK(n79527), .Q(n118543), .QN(
        n98525) );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n7415), .CK(n79527), .Q(n118542), .QN(
        n98526) );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n7414), .CK(n79527), .Q(n118541), .QN(
        n98527) );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n7413), .CK(n79527), .Q(n118540), .QN(
        n98528) );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n7412), .CK(n79527), .Q(n118539), .QN(
        n98529) );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n7411), .CK(n79527), .Q(n118538), .QN(
        n98530) );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n7410), .CK(n79527), .Q(n118537), .QN(
        n98531) );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n7409), .CK(n79527), .Q(n118536), .QN(
        n98532) );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n7408), .CK(n79527), .Q(n118535), .QN(
        n98533) );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n7407), .CK(n79527), .Q(n118534), .QN(
        n98534) );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n7406), .CK(n79527), .Q(n118533), .QN(
        n98535) );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n7405), .CK(n79527), .Q(n118532), .QN(
        n98536) );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n7404), .CK(n79527), .Q(n118531), .QN(
        n98537) );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n7403), .CK(n79527), .Q(n118530), .QN(
        n98538) );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n7402), .CK(n79527), .Q(n118529), .QN(
        n98539) );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n7401), .CK(n79527), .Q(n118528), .QN(
        n98540) );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n7400), .CK(n79527), .Q(n118527), .QN(
        n98541) );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n7399), .CK(n79527), .Q(n118526), .QN(
        n98542) );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n7398), .CK(n79527), .Q(n118525), .QN(
        n98543) );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n7397), .CK(n79527), .Q(n118524), .QN(
        n98544) );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n7396), .CK(n79527), .Q(n118523), .QN(
        n98545) );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n7395), .CK(n79527), .Q(n118522), .QN(
        n98546) );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n7394), .CK(n79527), .Q(n118521), .QN(
        n98547) );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n7393), .CK(n79527), .Q(n118520), .QN(
        n98548) );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n7392), .CK(n79527), .Q(n118519), .QN(
        n98549) );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n7391), .CK(n79527), .Q(n118518), .QN(
        n98550) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n7390), .CK(n79527), .Q(n118517), .QN(
        n98551) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n7389), .CK(n79527), .Q(n118516), .QN(
        n98552) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n7388), .CK(n79527), .Q(n118515), .QN(
        n98553) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n7387), .CK(n79527), .Q(n118514), .QN(
        n98554) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n7386), .CK(n79527), .Q(n118513), .QN(
        n98555) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n7385), .CK(n79527), .Q(n118512), .QN(
        n98556) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n7384), .CK(n79527), .Q(n118511), .QN(
        n98557) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n7383), .CK(n79527), .Q(n118510), .QN(
        n98558) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n7382), .CK(n79527), .Q(n118509), .QN(
        n98559) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n7381), .CK(n79527), .Q(n118508), .QN(
        n98560) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n7380), .CK(n79527), .Q(n118507), .QN(
        n98561) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n7379), .CK(n79527), .Q(n118506), .QN(
        n98562) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n7378), .CK(n79527), .Q(n118505), .QN(
        n98563) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n7377), .CK(n79527), .Q(n118805), .QN(
        n98564) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n7376), .CK(n79527), .Q(n118804), .QN(
        n98565) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n7375), .CK(n79527), .Q(n118803), .QN(
        n98566) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n7374), .CK(n79527), .Q(n118802), .QN(
        n98567) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n7373), .CK(n79527), .Q(n118801), .QN(
        n98568) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n7372), .CK(n79527), .Q(n118800), .QN(
        n98569) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n7371), .CK(n79527), .Q(n118799), .QN(
        n98570) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n7370), .CK(n79527), .Q(n118798), .QN(
        n98571) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n7369), .CK(n79527), .Q(n118809), .QN(
        n98572) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n7368), .CK(n79527), .Q(n118808), .QN(
        n98573) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n7367), .CK(n79527), .Q(n118807), .QN(
        n98574) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n7366), .CK(n79527), .Q(n118806), .QN(
        n98575) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n7365), .CK(n79527), .Q(n118816), .QN(
        n98576) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n7364), .CK(n79527), .Q(n118815), .QN(
        n98577) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n7363), .CK(n79527), .Q(n118814), .QN(
        n98578) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n7362), .CK(n79527), .Q(n118813), .QN(
        n98579) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n7361), .CK(n79527), .Q(n118812), .QN(
        n98580) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n7360), .CK(n79527), .Q(n118811), .QN(
        n98581) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n7359), .CK(n79527), .Q(n118810), .QN(
        n98582) );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n7098), .CK(n79527), .Q(n118751), .QN(
        n98848) );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n7097), .CK(n79527), .Q(n118750), .QN(
        n98849) );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n7096), .CK(n79527), .Q(n118749), .QN(
        n98850) );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n7095), .CK(n79527), .Q(n118748), .QN(
        n98851) );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n7094), .CK(n79527), .Q(n118747), .QN(
        n98852) );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n7093), .CK(n79527), .Q(n118746), .QN(
        n98853) );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n7092), .CK(n79527), .Q(n118745), .QN(
        n98854) );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n7091), .CK(n79527), .Q(n118744), .QN(
        n98855) );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n7090), .CK(n79527), .Q(n118743), .QN(
        n98856) );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n7089), .CK(n79527), .Q(n118742), .QN(
        n98857) );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n7088), .CK(n79527), .Q(n118741), .QN(
        n98858) );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n7087), .CK(n79527), .Q(n118740), .QN(
        n98859) );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n7086), .CK(n79527), .Q(n118739), .QN(
        n98860) );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n7085), .CK(n79527), .Q(n118738), .QN(
        n98861) );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n7084), .CK(n79527), .Q(n118797), .QN(
        n98862) );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n7083), .CK(n79527), .Q(n118796), .QN(
        n98863) );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n7082), .CK(n79527), .Q(n118795), .QN(
        n98864) );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n7081), .CK(n79527), .Q(n118794), .QN(
        n98865) );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n7080), .CK(n79527), .Q(n118793), .QN(
        n98866) );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n7079), .CK(n79527), .Q(n118792), .QN(
        n98867) );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n7078), .CK(n79527), .Q(n118791), .QN(
        n98868) );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n7077), .CK(n79527), .Q(n118790), .QN(
        n98869) );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n7076), .CK(n79527), .Q(n118789), .QN(
        n98870) );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n7075), .CK(n79527), .Q(n118788), .QN(
        n98871) );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n7074), .CK(n79527), .Q(n118787), .QN(
        n98872) );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n7073), .CK(n79527), .Q(n118786), .QN(
        n98873) );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n7072), .CK(n79527), .Q(n118785), .QN(
        n98874) );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n7071), .CK(n79527), .Q(n118784), .QN(
        n98875) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n7070), .CK(n79527), .Q(n118783), .QN(
        n98876) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n7069), .CK(n79527), .Q(n118782), .QN(
        n98877) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n7068), .CK(n79527), .Q(n118781), .QN(
        n98878) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n7067), .CK(n79527), .Q(n118780), .QN(
        n98879) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n7066), .CK(n79527), .Q(n118779), .QN(
        n98880) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n7065), .CK(n79527), .Q(n118778), .QN(
        n98881) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n7064), .CK(n79527), .Q(n118777), .QN(
        n98882) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n7063), .CK(n79527), .Q(n118776), .QN(
        n98883) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n7062), .CK(n79527), .Q(n118775), .QN(
        n98884) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n7061), .CK(n79527), .Q(n118774), .QN(
        n98885) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n7060), .CK(n79527), .Q(n118773), .QN(
        n98886) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n7059), .CK(n79527), .Q(n118772), .QN(
        n98887) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n7058), .CK(n79527), .Q(n118771), .QN(
        n98888) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n7057), .CK(n79527), .Q(n118770), .QN(
        n98889) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n7056), .CK(n79527), .Q(n118769), .QN(
        n98890) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n7055), .CK(n79527), .Q(n118768), .QN(
        n98891) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n7054), .CK(n79527), .Q(n118767), .QN(
        n98892) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n7053), .CK(n79527), .Q(n118766), .QN(
        n98893) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n7052), .CK(n79527), .Q(n118765), .QN(
        n98894) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n7051), .CK(n79527), .Q(n118764), .QN(
        n98895) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n7050), .CK(n79527), .Q(n118763), .QN(
        n98896) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n7049), .CK(n79527), .Q(n118762), .QN(
        n98897) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n7048), .CK(n79527), .Q(n118761), .QN(
        n98898) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n7047), .CK(n79527), .Q(n118760), .QN(
        n98899) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n7046), .CK(n79527), .Q(n118759), .QN(
        n98900) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n7045), .CK(n79527), .Q(n118758), .QN(
        n98901) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n7044), .CK(n79527), .Q(n118757), .QN(
        n98902) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n7043), .CK(n79527), .Q(n118756), .QN(
        n98903) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n7042), .CK(n79527), .Q(n118755), .QN(
        n98904) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n7041), .CK(n79527), .Q(n118754), .QN(
        n98905) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n7040), .CK(n79527), .Q(n118753), .QN(
        n98906) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n7039), .CK(n79527), .Q(n118752), .QN(
        n98907) );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n6842), .CK(n79527), .Q(n118970), .QN(
        n98986) );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n6841), .CK(n79527), .Q(n118969), .QN(
        n98987) );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n6840), .CK(n79527), .Q(n118968), .QN(
        n98988) );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n6839), .CK(n79527), .Q(n118967), .QN(
        n98989) );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n6838), .CK(n79527), .Q(n118966), .QN(
        n98990) );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n6837), .CK(n79527), .Q(n118965), .QN(
        n98991) );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n6836), .CK(n79527), .Q(n118964), .QN(
        n98992) );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n6835), .CK(n79527), .Q(n118963), .QN(
        n98993) );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n6834), .CK(n79527), .Q(n118962), .QN(
        n98994) );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n6833), .CK(n79527), .Q(n118961), .QN(
        n98995) );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n6832), .CK(n79527), .Q(n118960), .QN(
        n98996) );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n6831), .CK(n79527), .Q(n118959), .QN(
        n98997) );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n6830), .CK(n79527), .Q(n118958), .QN(
        n98998) );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n6829), .CK(n79527), .Q(n118957), .QN(
        n98999) );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n6828), .CK(n79527), .Q(n118956), .QN(
        n99000) );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n6827), .CK(n79527), .Q(n118955), .QN(
        n99001) );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n6826), .CK(n79527), .Q(n118954), .QN(
        n99002) );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n6825), .CK(n79527), .Q(n118953), .QN(
        n99003) );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n6824), .CK(n79527), .Q(n118952), .QN(
        n99004) );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n6823), .CK(n79527), .Q(n118951), .QN(
        n99005) );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n6822), .CK(n79527), .Q(n118950), .QN(
        n99006) );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n6821), .CK(n79527), .Q(n118949), .QN(
        n99007) );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n6820), .CK(n79527), .Q(n118948), .QN(
        n99008) );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n6819), .CK(n79527), .Q(n118947), .QN(
        n99009) );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n6818), .CK(n79527), .Q(n118946), .QN(
        n99010) );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n6817), .CK(n79527), .Q(n118945), .QN(
        n99011) );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n6816), .CK(n79527), .Q(n118944), .QN(
        n99012) );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n6815), .CK(n79527), .Q(n118943), .QN(
        n99013) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n6814), .CK(n79527), .Q(n118942), .QN(
        n99014) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n6813), .CK(n79527), .Q(n118941), .QN(
        n99015) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n6812), .CK(n79527), .Q(n118940), .QN(
        n99016) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n6811), .CK(n79527), .Q(n118939), .QN(
        n99017) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n6810), .CK(n79527), .Q(n118938), .QN(
        n99018) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n6809), .CK(n79527), .Q(n118937), .QN(
        n99019) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n6808), .CK(n79527), .Q(n118936), .QN(
        n99020) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n6807), .CK(n79527), .Q(n118935), .QN(
        n99021) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n6806), .CK(n79527), .Q(n118934), .QN(
        n99022) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n6805), .CK(n79527), .Q(n118933), .QN(
        n99023) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n6804), .CK(n79527), .Q(n118932), .QN(
        n99024) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n6803), .CK(n79527), .Q(n118931), .QN(
        n99025) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n6802), .CK(n79527), .Q(n118930), .QN(
        n99026) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n6801), .CK(n79527), .Q(n118929), .QN(
        n99027) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n6800), .CK(n79527), .Q(n118928), .QN(
        n99028) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n6799), .CK(n79527), .Q(n118927), .QN(
        n99029) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n6798), .CK(n79527), .Q(n118926), .QN(
        n99030) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n6797), .CK(n79527), .Q(n118925), .QN(
        n99031) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n6796), .CK(n79527), .Q(n118924), .QN(
        n99032) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n6795), .CK(n79527), .Q(n118923), .QN(
        n99033) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n6794), .CK(n79527), .Q(n118922), .QN(
        n99034) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n6793), .CK(n79527), .Q(n118974), .QN(
        n99035) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n6792), .CK(n79527), .Q(n118973), .QN(
        n99036) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n6791), .CK(n79527), .Q(n118972), .QN(
        n99037) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n6790), .CK(n79527), .Q(n118971), .QN(
        n99038) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n6789), .CK(n79527), .Q(n118981), .QN(
        n99039) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n6788), .CK(n79527), .Q(n118980), .QN(
        n99040) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n6787), .CK(n79527), .Q(n118979), .QN(
        n99041) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n6786), .CK(n79527), .Q(n118978), .QN(
        n99042) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n6785), .CK(n79527), .Q(n118977), .QN(
        n99043) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n6784), .CK(n79527), .Q(n118976), .QN(
        n99044) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n6783), .CK(n79527), .Q(n118975), .QN(
        n99045) );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n7226), .CK(n79527), .Q(n110539), .QN(
        n98719) );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n7225), .CK(n79527), .Q(n110538), .QN(
        n98720) );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n7224), .CK(n79527), .Q(n110537), .QN(
        n98721) );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n7223), .CK(n79527), .Q(n110536), .QN(
        n98722) );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n7222), .CK(n79527), .Q(n110535), .QN(
        n98723) );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n7221), .CK(n79527), .Q(n110534), .QN(
        n98724) );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n7220), .CK(n79527), .Q(n110533), .QN(
        n98725) );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n7219), .CK(n79527), .Q(n110532), .QN(
        n98726) );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n7218), .CK(n79527), .Q(n110531), .QN(
        n98727) );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n7217), .CK(n79527), .Q(n110530), .QN(
        n98728) );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n7216), .CK(n79527), .Q(n110529), .QN(
        n98729) );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n7215), .CK(n79527), .Q(n110528), .QN(
        n98730) );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n7214), .CK(n79527), .Q(n110527), .QN(
        n98731) );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n7213), .CK(n79527), .Q(n110526), .QN(
        n98732) );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n7212), .CK(n79527), .Q(n110525), .QN(
        n98733) );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n7211), .CK(n79527), .Q(n110524), .QN(
        n98734) );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n7210), .CK(n79527), .Q(n110523), .QN(
        n98735) );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n7209), .CK(n79527), .Q(n110522), .QN(
        n98736) );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n7208), .CK(n79527), .Q(n110521), .QN(
        n98737) );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n7207), .CK(n79527), .Q(n110520), .QN(
        n98738) );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n7206), .CK(n79527), .Q(n110519), .QN(
        n98739) );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n7205), .CK(n79527), .Q(n110518), .QN(
        n98740) );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n7204), .CK(n79527), .Q(n110517), .QN(
        n98741) );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n7203), .CK(n79527), .Q(n110516), .QN(
        n98742) );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n7202), .CK(n79527), .Q(n110515), .QN(
        n98743) );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n7201), .CK(n79527), .Q(n110514), .QN(
        n98744) );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n7200), .CK(n79527), .Q(n110513), .QN(
        n98745) );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n7199), .CK(n79527), .Q(n110512), .QN(
        n98746) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n7198), .CK(n79527), .Q(n110511), .QN(
        n98747) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n7197), .CK(n79527), .Q(n110510), .QN(
        n98748) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n7196), .CK(n79527), .Q(n110509), .QN(
        n98749) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n7195), .CK(n79527), .Q(n110508), .QN(
        n98750) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n7194), .CK(n79527), .Q(n110507), .QN(
        n98751) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n7193), .CK(n79527), .Q(n110506), .QN(
        n98752) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n7192), .CK(n79527), .Q(n110505), .QN(
        n98753) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n7191), .CK(n79527), .Q(n110504), .QN(
        n98754) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n7190), .CK(n79527), .Q(n110503), .QN(
        n98755) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n7189), .CK(n79527), .Q(n110502), .QN(
        n98756) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n7188), .CK(n79527), .Q(n110501), .QN(
        n98757) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n7187), .CK(n79527), .Q(n110500), .QN(
        n98758) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n7186), .CK(n79527), .Q(n110499), .QN(
        n98759) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n7185), .CK(n79527), .Q(n110498), .QN(
        n98760) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n7184), .CK(n79527), .Q(n110497), .QN(
        n98761) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n7183), .CK(n79527), .Q(n110496), .QN(
        n98762) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n7182), .CK(n79527), .Q(n110495), .QN(
        n98763) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n7181), .CK(n79527), .Q(n110494), .QN(
        n98764) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n7180), .CK(n79527), .Q(n110493), .QN(
        n98765) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n7179), .CK(n79527), .Q(n110492), .QN(
        n98766) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n7178), .CK(n79527), .Q(n110551), .QN(
        n98767) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n7177), .CK(n79527), .Q(n110550), .QN(
        n98768) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n7176), .CK(n79527), .Q(n110549), .QN(
        n98769) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n7175), .CK(n79527), .Q(n110548), .QN(
        n98770) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n7174), .CK(n79527), .Q(n110547), .QN(
        n98771) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n7173), .CK(n79527), .Q(n110558), .QN(
        n98772) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n7172), .CK(n79527), .Q(n110557), .QN(
        n98773) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n7171), .CK(n79527), .Q(n110556), .QN(
        n98774) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n7170), .CK(n79527), .Q(n110555), .QN(
        n98775) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n7169), .CK(n79527), .Q(n110554), .QN(
        n98776) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n7168), .CK(n79527), .Q(n110553), .QN(
        n98777) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n7167), .CK(n79527), .Q(n110552), .QN(
        n98778) );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n6586), .CK(n79527), .Q(n119191), .QN(
        n99250) );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n6585), .CK(n79527), .Q(n119190), .QN(
        n99251) );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n6584), .CK(n79527), .Q(n119189), .QN(
        n99252) );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n6583), .CK(n79527), .Q(n119188), .QN(
        n99253) );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n6582), .CK(n79527), .Q(n119187), .QN(
        n99254) );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n6581), .CK(n79527), .Q(n119186), .QN(
        n99255) );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n6580), .CK(n79527), .Q(n119185), .QN(
        n99256) );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n6579), .CK(n79527), .Q(n119184), .QN(
        n99257) );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n6578), .CK(n79527), .Q(n119183), .QN(
        n99258) );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n6577), .CK(n79527), .Q(n119182), .QN(
        n99259) );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n6576), .CK(n79527), .Q(n119181), .QN(
        n99260) );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n6575), .CK(n79527), .Q(n119180), .QN(
        n99261) );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n6574), .CK(n79527), .Q(n119179), .QN(
        n99262) );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n6573), .CK(n79527), .Q(n119178), .QN(
        n99263) );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n6572), .CK(n79527), .Q(n119237), .QN(
        n99264) );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n6571), .CK(n79527), .Q(n119236), .QN(
        n99265) );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n6570), .CK(n79527), .Q(n119235), .QN(
        n99266) );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n6569), .CK(n79527), .Q(n119234), .QN(
        n99267) );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n6568), .CK(n79527), .Q(n119233), .QN(
        n99268) );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n6567), .CK(n79527), .Q(n119232), .QN(
        n99269) );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n6566), .CK(n79527), .Q(n119231), .QN(
        n99270) );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n6565), .CK(n79527), .Q(n119230), .QN(
        n99271) );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n6564), .CK(n79527), .Q(n119229), .QN(
        n99272) );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n6563), .CK(n79527), .Q(n119228), .QN(
        n99273) );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n6562), .CK(n79527), .Q(n119227), .QN(
        n99274) );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n6561), .CK(n79527), .Q(n119226), .QN(
        n99275) );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n6560), .CK(n79527), .Q(n119225), .QN(
        n99276) );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n6559), .CK(n79527), .Q(n119224), .QN(
        n99277) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n6558), .CK(n79527), .Q(n119223), .QN(
        n99278) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n6557), .CK(n79527), .Q(n119222), .QN(
        n99279) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n6556), .CK(n79527), .Q(n119221), .QN(
        n99280) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n6555), .CK(n79527), .Q(n119220), .QN(
        n99281) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n6554), .CK(n79527), .Q(n119219), .QN(
        n99282) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n6553), .CK(n79527), .Q(n119218), .QN(
        n99283) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n6552), .CK(n79527), .Q(n119217), .QN(
        n99284) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n6551), .CK(n79527), .Q(n119216), .QN(
        n99285) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n6550), .CK(n79527), .Q(n119215), .QN(
        n99286) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n6549), .CK(n79527), .Q(n119214), .QN(
        n99287) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n6548), .CK(n79527), .Q(n119213), .QN(
        n99288) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n6547), .CK(n79527), .Q(n119212), .QN(
        n99289) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n6546), .CK(n79527), .Q(n119211), .QN(
        n99290) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n6545), .CK(n79527), .Q(n119210), .QN(
        n99291) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n6544), .CK(n79527), .Q(n119209), .QN(
        n99292) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n6543), .CK(n79527), .Q(n119208), .QN(
        n99293) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n6542), .CK(n79527), .Q(n119207), .QN(
        n99294) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n6541), .CK(n79527), .Q(n119206), .QN(
        n99295) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n6540), .CK(n79527), .Q(n119205), .QN(
        n99296) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n6539), .CK(n79527), .Q(n119204), .QN(
        n99297) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n6538), .CK(n79527), .Q(n119203), .QN(
        n99298) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n6537), .CK(n79527), .Q(n119202), .QN(
        n99299) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n6536), .CK(n79527), .Q(n119201), .QN(
        n99300) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n6535), .CK(n79527), .Q(n119200), .QN(
        n99301) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n6534), .CK(n79527), .Q(n119199), .QN(
        n99302) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n6533), .CK(n79527), .Q(n119198), .QN(
        n99303) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n6532), .CK(n79527), .Q(n119197), .QN(
        n99304) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n6531), .CK(n79527), .Q(n119196), .QN(
        n99305) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n6530), .CK(n79527), .Q(n119195), .QN(
        n99306) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n6529), .CK(n79527), .Q(n119194), .QN(
        n99307) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n6528), .CK(n79527), .Q(n119193), .QN(
        n99308) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n6527), .CK(n79527), .Q(n119192), .QN(
        n99309) );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n6714), .CK(n79527), .Q(n119350), .QN(
        n99118) );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n6713), .CK(n79527), .Q(n119349), .QN(
        n99119) );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n6712), .CK(n79527), .Q(n119348), .QN(
        n99120) );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n6711), .CK(n79527), .Q(n119347), .QN(
        n99121) );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n6710), .CK(n79527), .Q(n119346), .QN(
        n99122) );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n6709), .CK(n79527), .Q(n119345), .QN(
        n99123) );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n6708), .CK(n79527), .Q(n119344), .QN(
        n99124) );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n6707), .CK(n79527), .Q(n119343), .QN(
        n99125) );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n6706), .CK(n79527), .Q(n119342), .QN(
        n99126) );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n6705), .CK(n79527), .Q(n119341), .QN(
        n99127) );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n6704), .CK(n79527), .Q(n119340), .QN(
        n99128) );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n6703), .CK(n79527), .Q(n119339), .QN(
        n99129) );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n6702), .CK(n79527), .Q(n119338), .QN(
        n99130) );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n6701), .CK(n79527), .Q(n119337), .QN(
        n99131) );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n6700), .CK(n79527), .Q(n119336), .QN(
        n99132) );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n6699), .CK(n79527), .Q(n119335), .QN(
        n99133) );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n6698), .CK(n79527), .Q(n119334), .QN(
        n99134) );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n6697), .CK(n79527), .Q(n119333), .QN(
        n99135) );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n6696), .CK(n79527), .Q(n119332), .QN(
        n99136) );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n6695), .CK(n79527), .Q(n119331), .QN(
        n99137) );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n6694), .CK(n79527), .Q(n119330), .QN(
        n99138) );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n6693), .CK(n79527), .Q(n119329), .QN(
        n99139) );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n6692), .CK(n79527), .Q(n119328), .QN(
        n99140) );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n6691), .CK(n79527), .Q(n119327), .QN(
        n99141) );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n6690), .CK(n79527), .Q(n119326), .QN(
        n99142) );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n6689), .CK(n79527), .Q(n119325), .QN(
        n99143) );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n6688), .CK(n79527), .Q(n119324), .QN(
        n99144) );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n6687), .CK(n79527), .Q(n119323), .QN(
        n99145) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n6686), .CK(n79527), .Q(n119322), .QN(
        n99146) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n6685), .CK(n79527), .Q(n119321), .QN(
        n99147) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n6684), .CK(n79527), .Q(n119320), .QN(
        n99148) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n6683), .CK(n79527), .Q(n119319), .QN(
        n99149) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n6682), .CK(n79527), .Q(n119318), .QN(
        n99150) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n6681), .CK(n79527), .Q(n119317), .QN(
        n99151) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n6680), .CK(n79527), .Q(n119316), .QN(
        n99152) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n6679), .CK(n79527), .Q(n119315), .QN(
        n99153) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n6678), .CK(n79527), .Q(n119314), .QN(
        n99154) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n6677), .CK(n79527), .Q(n119313), .QN(
        n99155) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n6676), .CK(n79527), .Q(n119312), .QN(
        n99156) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n6675), .CK(n79527), .Q(n119311), .QN(
        n99157) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n6674), .CK(n79527), .Q(n119310), .QN(
        n99158) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n6673), .CK(n79527), .Q(n119309), .QN(
        n99159) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n6672), .CK(n79527), .Q(n119308), .QN(
        n99160) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n6671), .CK(n79527), .Q(n119307), .QN(
        n99161) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n6670), .CK(n79527), .Q(n119306), .QN(
        n99162) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n6669), .CK(n79527), .Q(n119305), .QN(
        n99163) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n6668), .CK(n79527), .Q(n119304), .QN(
        n99164) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n6667), .CK(n79527), .Q(n119303), .QN(
        n99165) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n6666), .CK(n79527), .Q(n119302), .QN(
        n99166) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n6665), .CK(n79527), .Q(n119358), .QN(
        n99167) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n6664), .CK(n79527), .Q(n119357), .QN(
        n99168) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n6663), .CK(n79527), .Q(n119356), .QN(
        n99169) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n6662), .CK(n79527), .Q(n119355), .QN(
        n99170) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n6661), .CK(n79527), .Q(n119365), .QN(
        n99171) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n6660), .CK(n79527), .Q(n119364), .QN(
        n99172) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n6659), .CK(n79527), .Q(n119363), .QN(
        n99173) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n6658), .CK(n79527), .Q(n119362), .QN(
        n99174) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n6657), .CK(n79527), .Q(n119361), .QN(
        n99175) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n6656), .CK(n79527), .Q(n119360), .QN(
        n99176) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n6655), .CK(n79527), .Q(n119359), .QN(
        n99177) );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n6778), .CK(n79527), .Q(n110572), .QN(
        n99052) );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n6777), .CK(n79527), .Q(n110571), .QN(
        n99053) );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n6776), .CK(n79527), .Q(n110570), .QN(
        n99054) );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n6775), .CK(n79527), .Q(n110569), .QN(
        n99055) );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n6774), .CK(n79527), .Q(n110568), .QN(
        n99056) );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n6773), .CK(n79527), .Q(n110567), .QN(
        n99057) );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n6772), .CK(n79527), .Q(n110566), .QN(
        n99058) );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n6771), .CK(n79527), .Q(n110565), .QN(
        n99059) );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n6770), .CK(n79527), .Q(n110564), .QN(
        n99060) );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n6769), .CK(n79527), .Q(n110563), .QN(
        n99061) );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n6768), .CK(n79527), .Q(n110562), .QN(
        n99062) );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n6767), .CK(n79527), .Q(n110561), .QN(
        n99063) );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n6766), .CK(n79527), .Q(n110560), .QN(
        n99064) );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n6765), .CK(n79527), .Q(n110559), .QN(
        n99065) );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n6764), .CK(n79527), .Q(n110622), .QN(
        n99066) );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n6763), .CK(n79527), .Q(n110621), .QN(
        n99067) );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n6762), .CK(n79527), .Q(n110620), .QN(
        n99068) );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n6761), .CK(n79527), .Q(n110619), .QN(
        n99069) );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n6760), .CK(n79527), .Q(n110618), .QN(
        n99070) );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n6759), .CK(n79527), .Q(n110617), .QN(
        n99071) );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n6758), .CK(n79527), .Q(n110616), .QN(
        n99072) );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n6757), .CK(n79527), .Q(n110615), .QN(
        n99073) );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n6756), .CK(n79527), .Q(n110614), .QN(
        n99074) );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n6755), .CK(n79527), .Q(n110613), .QN(
        n99075) );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n6754), .CK(n79527), .Q(n110612), .QN(
        n99076) );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n6753), .CK(n79527), .Q(n110611), .QN(
        n99077) );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n6752), .CK(n79527), .Q(n110610), .QN(
        n99078) );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n6751), .CK(n79527), .Q(n110609), .QN(
        n99079) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n6750), .CK(n79527), .Q(n110608), .QN(
        n99080) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n6749), .CK(n79527), .Q(n110607), .QN(
        n99081) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n6748), .CK(n79527), .Q(n110606), .QN(
        n99082) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n6747), .CK(n79527), .Q(n110605), .QN(
        n99083) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n6746), .CK(n79527), .Q(n110604), .QN(
        n99084) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n6745), .CK(n79527), .Q(n110603), .QN(
        n99085) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n6744), .CK(n79527), .Q(n110602), .QN(
        n99086) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n6743), .CK(n79527), .Q(n110601), .QN(
        n99087) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n6742), .CK(n79527), .Q(n110600), .QN(
        n99088) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n6741), .CK(n79527), .Q(n110599), .QN(
        n99089) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n6740), .CK(n79527), .Q(n110598), .QN(
        n99090) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n6739), .CK(n79527), .Q(n110597), .QN(
        n99091) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n6738), .CK(n79527), .Q(n110596), .QN(
        n99092) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n6737), .CK(n79527), .Q(n110595), .QN(
        n99093) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n6736), .CK(n79527), .Q(n110594), .QN(
        n99094) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n6735), .CK(n79527), .Q(n110593), .QN(
        n99095) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n6734), .CK(n79527), .Q(n110592), .QN(
        n99096) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n6733), .CK(n79527), .Q(n110591), .QN(
        n99097) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n6732), .CK(n79527), .Q(n110590), .QN(
        n99098) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n6731), .CK(n79527), .Q(n110589), .QN(
        n99099) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n6730), .CK(n79527), .Q(n110588), .QN(
        n99100) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n6729), .CK(n79527), .Q(n110587), .QN(
        n99101) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n6728), .CK(n79527), .Q(n110586), .QN(
        n99102) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n6727), .CK(n79527), .Q(n110585), .QN(
        n99103) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n6726), .CK(n79527), .Q(n110584), .QN(
        n99104) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n6725), .CK(n79527), .Q(n110583), .QN(
        n99105) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n6724), .CK(n79527), .Q(n110582), .QN(
        n99106) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n6723), .CK(n79527), .Q(n110581), .QN(
        n99107) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n6722), .CK(n79527), .Q(n110576), .QN(
        n99108) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n6721), .CK(n79527), .Q(n110575), .QN(
        n99109) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n6720), .CK(n79527), .Q(n110574), .QN(
        n99110) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n6719), .CK(n79527), .Q(n110573), .QN(
        n99111) );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n6522), .CK(n79527), .Q(n119251), .QN(
        n99316) );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n6521), .CK(n79527), .Q(n119250), .QN(
        n99317) );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n6520), .CK(n79527), .Q(n119249), .QN(
        n99318) );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n6519), .CK(n79527), .Q(n119248), .QN(
        n99319) );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n6518), .CK(n79527), .Q(n119247), .QN(
        n99320) );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n6517), .CK(n79527), .Q(n119246), .QN(
        n99321) );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n6516), .CK(n79527), .Q(n119245), .QN(
        n99322) );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n6515), .CK(n79527), .Q(n119244), .QN(
        n99323) );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n6514), .CK(n79527), .Q(n119243), .QN(
        n99324) );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n6513), .CK(n79527), .Q(n119242), .QN(
        n99325) );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n6512), .CK(n79527), .Q(n119241), .QN(
        n99326) );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n6511), .CK(n79527), .Q(n119240), .QN(
        n99327) );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n6510), .CK(n79527), .Q(n119239), .QN(
        n99328) );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n6509), .CK(n79527), .Q(n119238), .QN(
        n99329) );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n6508), .CK(n79527), .Q(n119285), .QN(
        n99330) );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n6507), .CK(n79527), .Q(n119284), .QN(
        n99331) );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n6506), .CK(n79527), .Q(n119283), .QN(
        n99332) );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n6505), .CK(n79527), .Q(n119282), .QN(
        n99333) );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n6504), .CK(n79527), .Q(n119281), .QN(
        n99334) );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n6503), .CK(n79527), .Q(n119280), .QN(
        n99335) );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n6502), .CK(n79527), .Q(n119279), .QN(
        n99336) );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n6501), .CK(n79527), .Q(n119278), .QN(
        n99337) );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n6500), .CK(n79527), .Q(n119277), .QN(
        n99338) );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n6499), .CK(n79527), .Q(n119276), .QN(
        n99339) );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n6498), .CK(n79527), .Q(n119275), .QN(
        n99340) );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n6497), .CK(n79527), .Q(n119274), .QN(
        n99341) );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n6496), .CK(n79527), .Q(n119273), .QN(
        n99342) );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n6495), .CK(n79527), .Q(n119272), .QN(
        n99343) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n6494), .CK(n79527), .Q(n119271), .QN(
        n99344) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n6493), .CK(n79527), .Q(n119270), .QN(
        n99345) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n6492), .CK(n79527), .Q(n119269), .QN(
        n99346) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n6491), .CK(n79527), .Q(n119268), .QN(
        n99347) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n6490), .CK(n79527), .Q(n119267), .QN(
        n99348) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n6489), .CK(n79527), .Q(n119266), .QN(
        n99349) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n6488), .CK(n79527), .Q(n119265), .QN(
        n99350) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n6487), .CK(n79527), .Q(n119264), .QN(
        n99351) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n6486), .CK(n79527), .Q(n119263), .QN(
        n99352) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n6485), .CK(n79527), .Q(n119262), .QN(
        n99353) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n6484), .CK(n79527), .Q(n119261), .QN(
        n99354) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n6483), .CK(n79527), .Q(n119260), .QN(
        n99355) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n6482), .CK(n79527), .Q(n119259), .QN(
        n99356) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n6481), .CK(n79527), .Q(n119258), .QN(
        n99357) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n6480), .CK(n79527), .Q(n119257), .QN(
        n99358) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n6479), .CK(n79527), .Q(n119256), .QN(
        n99359) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n6478), .CK(n79527), .Q(n119255), .QN(
        n99360) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n6477), .CK(n79527), .Q(n119254), .QN(
        n99361) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n6476), .CK(n79527), .Q(n119253), .QN(
        n99362) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n6475), .CK(n79527), .Q(n119252), .QN(
        n99363) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n6474), .CK(n79527), .Q(n119297), .QN(
        n99364) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n6473), .CK(n79527), .Q(n119296), .QN(
        n99365) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n6472), .CK(n79527), .Q(n119295), .QN(
        n99366) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n6471), .CK(n79527), .Q(n119294), .QN(
        n99367) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n6470), .CK(n79527), .Q(n119293), .QN(
        n99368) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n6469), .CK(n79527), .Q(n119292), .QN(
        n99369) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n6468), .CK(n79527), .Q(n119291), .QN(
        n99370) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n6467), .CK(n79527), .Q(n119290), .QN(
        n99371) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n6466), .CK(n79527), .Q(n119289), .QN(
        n99372) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n6465), .CK(n79527), .Q(n119288), .QN(
        n99373) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n6464), .CK(n79527), .Q(n119287), .QN(
        n99374) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n6463), .CK(n79527), .Q(n119286), .QN(
        n99375) );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n6650), .CK(n79527), .Q(n119127), .QN(
        n99184) );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n6649), .CK(n79527), .Q(n119126), .QN(
        n99185) );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n6648), .CK(n79527), .Q(n119125), .QN(
        n99186) );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n6647), .CK(n79527), .Q(n119124), .QN(
        n99187) );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n6646), .CK(n79527), .Q(n119123), .QN(
        n99188) );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n6645), .CK(n79527), .Q(n119122), .QN(
        n99189) );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n6644), .CK(n79527), .Q(n119121), .QN(
        n99190) );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n6643), .CK(n79527), .Q(n119120), .QN(
        n99191) );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n6642), .CK(n79527), .Q(n119119), .QN(
        n99192) );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n6641), .CK(n79527), .Q(n119118), .QN(
        n99193) );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n6640), .CK(n79527), .Q(n119117), .QN(
        n99194) );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n6639), .CK(n79527), .Q(n119116), .QN(
        n99195) );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n6638), .CK(n79527), .Q(n119115), .QN(
        n99196) );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n6637), .CK(n79527), .Q(n119114), .QN(
        n99197) );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n6636), .CK(n79527), .Q(n119173), .QN(
        n99198) );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n6635), .CK(n79527), .Q(n119172), .QN(
        n99199) );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n6634), .CK(n79527), .Q(n119171), .QN(
        n99200) );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n6633), .CK(n79527), .Q(n119170), .QN(
        n99201) );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n6632), .CK(n79527), .Q(n119169), .QN(
        n99202) );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n6631), .CK(n79527), .Q(n119168), .QN(
        n99203) );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n6630), .CK(n79527), .Q(n119167), .QN(
        n99204) );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n6629), .CK(n79527), .Q(n119166), .QN(
        n99205) );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n6628), .CK(n79527), .Q(n119165), .QN(
        n99206) );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n6627), .CK(n79527), .Q(n119164), .QN(
        n99207) );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n6626), .CK(n79527), .Q(n119163), .QN(
        n99208) );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n6625), .CK(n79527), .Q(n119162), .QN(
        n99209) );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n6624), .CK(n79527), .Q(n119161), .QN(
        n99210) );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n6623), .CK(n79527), .Q(n119160), .QN(
        n99211) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n6622), .CK(n79527), .Q(n119159), .QN(
        n99212) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n6621), .CK(n79527), .Q(n119158), .QN(
        n99213) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n6620), .CK(n79527), .Q(n119157), .QN(
        n99214) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n6619), .CK(n79527), .Q(n119156), .QN(
        n99215) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n6618), .CK(n79527), .Q(n119155), .QN(
        n99216) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n6617), .CK(n79527), .Q(n119154), .QN(
        n99217) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n6616), .CK(n79527), .Q(n119153), .QN(
        n99218) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n6615), .CK(n79527), .Q(n119152), .QN(
        n99219) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n6614), .CK(n79527), .Q(n119151), .QN(
        n99220) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n6613), .CK(n79527), .Q(n119150), .QN(
        n99221) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n6612), .CK(n79527), .Q(n119149), .QN(
        n99222) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n6611), .CK(n79527), .Q(n119148), .QN(
        n99223) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n6610), .CK(n79527), .Q(n119147), .QN(
        n99224) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n6609), .CK(n79527), .Q(n119146), .QN(
        n99225) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n6608), .CK(n79527), .Q(n119145), .QN(
        n99226) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n6607), .CK(n79527), .Q(n119144), .QN(
        n99227) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n6606), .CK(n79527), .Q(n119143), .QN(
        n99228) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n6605), .CK(n79527), .Q(n119142), .QN(
        n99229) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n6604), .CK(n79527), .Q(n119141), .QN(
        n99230) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n6603), .CK(n79527), .Q(n119140), .QN(
        n99231) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n6602), .CK(n79527), .Q(n119139), .QN(
        n99232) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n6601), .CK(n79527), .Q(n119138), .QN(
        n99233) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n6600), .CK(n79527), .Q(n119137), .QN(
        n99234) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n6599), .CK(n79527), .Q(n119136), .QN(
        n99235) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n6598), .CK(n79527), .Q(n119135), .QN(
        n99236) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n6597), .CK(n79527), .Q(n119134), .QN(
        n99237) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n6596), .CK(n79527), .Q(n119133), .QN(
        n99238) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n6595), .CK(n79527), .Q(n119132), .QN(
        n99239) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n6594), .CK(n79527), .Q(n119131), .QN(
        n99240) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n6593), .CK(n79527), .Q(n119130), .QN(
        n99241) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n6592), .CK(n79527), .Q(n119129), .QN(
        n99242) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n6591), .CK(n79527), .Q(n119128), .QN(
        n99243) );
  DFF_X1 \OUT1_reg[3]  ( .D(n5381), .CK(n79527), .Q(OUT1[3]) );
  DFF_X1 \OUT1_reg[2]  ( .D(n5379), .CK(n79527), .Q(OUT1[2]) );
  DFF_X1 \OUT1_reg[1]  ( .D(n5377), .CK(n79527), .Q(OUT1[1]) );
  DFF_X1 \OUT1_reg[0]  ( .D(n5375), .CK(n79527), .Q(OUT1[0]) );
  DFF_X1 \OUT1_reg[59]  ( .D(n5493), .CK(n79527), .Q(OUT1[59]) );
  DFF_X1 \OUT1_reg[58]  ( .D(n5491), .CK(n79527), .Q(OUT1[58]) );
  DFF_X1 \OUT1_reg[57]  ( .D(n5489), .CK(n79527), .Q(OUT1[57]) );
  DFF_X1 \OUT1_reg[56]  ( .D(n5487), .CK(n79527), .Q(OUT1[56]) );
  DFF_X1 \OUT1_reg[55]  ( .D(n5485), .CK(n79527), .Q(OUT1[55]) );
  DFF_X1 \OUT1_reg[54]  ( .D(n5483), .CK(n79527), .Q(OUT1[54]) );
  DFF_X1 \OUT1_reg[53]  ( .D(n5481), .CK(n79527), .Q(OUT1[53]) );
  DFF_X1 \OUT1_reg[52]  ( .D(n5479), .CK(n79527), .Q(OUT1[52]) );
  DFF_X1 \OUT1_reg[51]  ( .D(n5477), .CK(n79527), .Q(OUT1[51]) );
  DFF_X1 \OUT1_reg[50]  ( .D(n5475), .CK(n79527), .Q(OUT1[50]) );
  DFF_X1 \OUT1_reg[49]  ( .D(n5473), .CK(n79527), .Q(OUT1[49]) );
  DFF_X1 \OUT1_reg[48]  ( .D(n5471), .CK(n79527), .Q(OUT1[48]) );
  DFF_X1 \OUT1_reg[47]  ( .D(n5469), .CK(n79527), .Q(OUT1[47]) );
  DFF_X1 \OUT1_reg[46]  ( .D(n5467), .CK(n79527), .Q(OUT1[46]) );
  DFF_X1 \OUT2_reg[29]  ( .D(n5340), .CK(n79527), .Q(OUT2[29]) );
  DFF_X1 \OUT2_reg[28]  ( .D(n5339), .CK(n79527), .Q(OUT2[28]) );
  DFF_X1 \OUT2_reg[27]  ( .D(n5338), .CK(n79527), .Q(OUT2[27]) );
  DFF_X1 \OUT2_reg[26]  ( .D(n5337), .CK(n79527), .Q(OUT2[26]) );
  DFF_X1 \OUT2_reg[25]  ( .D(n5336), .CK(n79527), .Q(OUT2[25]) );
  DFF_X1 \OUT2_reg[24]  ( .D(n5335), .CK(n79527), .Q(OUT2[24]) );
  DFF_X1 \OUT2_reg[23]  ( .D(n5334), .CK(n79527), .Q(OUT2[23]) );
  DFF_X1 \OUT2_reg[22]  ( .D(n5333), .CK(n79527), .Q(OUT2[22]) );
  DFF_X1 \OUT2_reg[21]  ( .D(n5332), .CK(n79527), .Q(OUT2[21]) );
  DFF_X1 \OUT2_reg[20]  ( .D(n5331), .CK(n79527), .Q(OUT2[20]) );
  DFF_X1 \OUT2_reg[19]  ( .D(n5330), .CK(n79527), .Q(OUT2[19]) );
  DFF_X1 \OUT2_reg[18]  ( .D(n5329), .CK(n79527), .Q(OUT2[18]) );
  DFF_X1 \OUT2_reg[17]  ( .D(n5328), .CK(n79527), .Q(OUT2[17]) );
  DFF_X1 \OUT2_reg[16]  ( .D(n5327), .CK(n79527), .Q(OUT2[16]) );
  DFF_X1 \OUT2_reg[15]  ( .D(n5326), .CK(n79527), .Q(OUT2[15]) );
  DFF_X1 \OUT2_reg[14]  ( .D(n5325), .CK(n79527), .Q(OUT2[14]) );
  DFF_X1 \OUT2_reg[13]  ( .D(n5324), .CK(n79527), .Q(OUT2[13]) );
  DFF_X1 \OUT2_reg[12]  ( .D(n5323), .CK(n79527), .Q(OUT2[12]) );
  DFF_X1 \OUT2_reg[11]  ( .D(n5322), .CK(n79527), .Q(OUT2[11]) );
  NOR3_X2 U81228 ( .A1(n120216), .A2(ADD_RD1[1]), .A3(n116475), .ZN(n116457)
         );
  NOR3_X2 U81241 ( .A1(n120216), .A2(ADD_RD1[2]), .A3(n116478), .ZN(n116453)
         );
  NAND3_X1 U83316 ( .A1(n113987), .A2(n113988), .A3(n113989), .ZN(n113893) );
  NAND3_X1 U83317 ( .A1(n113989), .A2(n113988), .A3(ADD_WR[0]), .ZN(n113901)
         );
  NAND3_X1 U83318 ( .A1(n113989), .A2(n113987), .A3(ADD_WR[3]), .ZN(n114054)
         );
  NAND3_X1 U83319 ( .A1(ADD_WR[0]), .A2(n113989), .A3(ADD_WR[3]), .ZN(n114121)
         );
  NAND3_X1 U83320 ( .A1(n113987), .A2(n113988), .A3(n114302), .ZN(n114141) );
  NAND3_X1 U83321 ( .A1(ADD_WR[0]), .A2(n113988), .A3(n114302), .ZN(n114144)
         );
  NAND3_X1 U83322 ( .A1(ADD_WR[3]), .A2(n113987), .A3(n114302), .ZN(n114371)
         );
  NAND3_X1 U83323 ( .A1(ADD_WR[3]), .A2(ADD_WR[0]), .A3(n114302), .ZN(n114374)
         );
  NAND3_X1 U83324 ( .A1(ENABLE), .A2(n120628), .A3(RD1), .ZN(n114658) );
  NAND3_X1 U83325 ( .A1(ENABLE), .A2(n120628), .A3(RD2), .ZN(n116491) );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n5502), .CK(n79527), .Q(n95528), .QN(
        n114644) );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n5500), .CK(n79527), .Q(n95527), .QN(
        n114704) );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n5498), .CK(n79527), .Q(n95526), .QN(
        n114730) );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n5496), .CK(n79527), .Q(n95525), .QN(
        n114756) );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n5566), .CK(n79527), .Q(n117996), .QN(
        n114578) );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n5565), .CK(n79527), .Q(n117995), .QN(
        n114580) );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n5564), .CK(n79527), .Q(n117994), .QN(
        n114581) );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n5563), .CK(n79527), .Q(n117993), .QN(
        n114582) );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n5694), .CK(n79527), .QN(n114510) );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n5693), .CK(n79527), .QN(n114512) );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n5692), .CK(n79527), .QN(n114513) );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n5691), .CK(n79527), .QN(n114514) );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n5758), .CK(n79527), .QN(n114444) );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n5757), .CK(n79527), .QN(n114446) );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n5756), .CK(n79527), .QN(n114447) );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n5755), .CK(n79527), .QN(n114448) );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n5822), .CK(n79527), .QN(n114378) );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n5821), .CK(n79527), .QN(n114380) );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n5820), .CK(n79527), .QN(n114381) );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n5819), .CK(n79527), .QN(n114382) );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n5950), .CK(n79527), .Q(n117988), .QN(
        n114306) );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n5949), .CK(n79527), .Q(n117987), .QN(
        n114308) );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n5948), .CK(n79527), .Q(n117986), .QN(
        n114309) );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n5947), .CK(n79527), .Q(n117985), .QN(
        n114310) );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n6142), .CK(n79527), .Q(n117984), .QN(
        n114235) );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n6141), .CK(n79527), .Q(n117983), .QN(
        n114237) );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n6140), .CK(n79527), .Q(n117982), .QN(
        n114238) );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n6139), .CK(n79527), .Q(n117981), .QN(
        n114239) );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n6334), .CK(n79527), .QN(n114146) );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n6333), .CK(n79527), .QN(n114148) );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n6332), .CK(n79527), .QN(n114149) );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n6331), .CK(n79527), .QN(n114150) );
  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n7358), .CK(n79527), .Q(n109906), .QN(
        n113903) );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n7357), .CK(n79527), .Q(n109905), .QN(
        n113905) );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n7356), .CK(n79527), .Q(n109904), .QN(
        n113906) );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n7355), .CK(n79527), .Q(n109903), .QN(
        n113907) );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n7102), .CK(n79527), .Q(n111048), .QN(
        n113981) );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n7101), .CK(n79527), .Q(n111047), .QN(
        n113983) );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n7100), .CK(n79527), .Q(n111046), .QN(
        n113984) );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n7099), .CK(n79527), .Q(n111045), .QN(
        n113985) );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n7422), .CK(n79527), .Q(n109898), .QN(
        n113896) );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n7421), .CK(n79527), .Q(n109897), .QN(
        n113898) );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n7420), .CK(n79527), .Q(n109896), .QN(
        n113899) );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n7419), .CK(n79527), .Q(n109895), .QN(
        n113900) );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n6846), .CK(n79527), .Q(n111044), .QN(
        n114123) );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n6845), .CK(n79527), .Q(n111043), .QN(
        n114125) );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n6844), .CK(n79527), .Q(n111042), .QN(
        n114126) );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n6843), .CK(n79527), .Q(n111041), .QN(
        n114127) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n6161), .CK(n79527), .Q(n109997), .QN(
        n114215) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n6160), .CK(n79527), .Q(n109996), .QN(
        n114216) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n6159), .CK(n79527), .Q(n109995), .QN(
        n114217) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n6158), .CK(n79527), .Q(n109994), .QN(
        n114218) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n6157), .CK(n79527), .Q(n109993), .QN(
        n114219) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n6156), .CK(n79527), .Q(n109992), .QN(
        n114220) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n6155), .CK(n79527), .Q(n109991), .QN(
        n114221) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n6154), .CK(n79527), .Q(n109990), .QN(
        n114222) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n6153), .CK(n79527), .Q(n109989), .QN(
        n114223) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n6152), .CK(n79527), .Q(n109988), .QN(
        n114224) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n6151), .CK(n79527), .Q(n109987), .QN(
        n114225) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n6150), .CK(n79527), .Q(n109986), .QN(
        n114226) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n6149), .CK(n79527), .Q(n109985), .QN(
        n114227) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n6148), .CK(n79527), .Q(n109984), .QN(
        n114228) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n6147), .CK(n79527), .Q(n109983), .QN(
        n114229) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n6146), .CK(n79527), .Q(n109982), .QN(
        n114230) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n6145), .CK(n79527), .Q(n109981), .QN(
        n114231) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n6144), .CK(n79527), .Q(n109980), .QN(
        n114232) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n6143), .CK(n79527), .Q(n109979), .QN(
        n114233) );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n7166), .CK(n79527), .QN(n113915) );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n7165), .CK(n79527), .QN(n113917) );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n7164), .CK(n79527), .QN(n113918) );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n7163), .CK(n79527), .QN(n113919) );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n5494), .CK(n79527), .Q(n95488), .QN(
        n114782) );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n5492), .CK(n79527), .Q(n95487), .QN(
        n114810) );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n5490), .CK(n79527), .Q(n95486), .QN(
        n114838) );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n5488), .CK(n79527), .Q(n95485), .QN(
        n114866) );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n5486), .CK(n79527), .Q(n95484), .QN(
        n114894) );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n5484), .CK(n79527), .Q(n95483), .QN(
        n114922) );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n5482), .CK(n79527), .Q(n95482), .QN(
        n114950) );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n5480), .CK(n79527), .Q(n95481), .QN(
        n114978) );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n5478), .CK(n79527), .Q(n95480), .QN(
        n115006) );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n5476), .CK(n79527), .Q(n95479), .QN(
        n115034) );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n5474), .CK(n79527), .Q(n95478), .QN(
        n115062) );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n5472), .CK(n79527), .Q(n95477), .QN(
        n115090) );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n5470), .CK(n79527), .Q(n95476), .QN(
        n115118) );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n5468), .CK(n79527), .Q(n95475), .QN(
        n115146) );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n5466), .CK(n79527), .Q(n95474), .QN(
        n115174) );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n5464), .CK(n79527), .Q(n95473), .QN(
        n115202) );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n5462), .CK(n79527), .Q(n95472), .QN(
        n115230) );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n5460), .CK(n79527), .Q(n95471), .QN(
        n115258) );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n5458), .CK(n79527), .Q(n95470), .QN(
        n115286) );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n5456), .CK(n79527), .Q(n95469), .QN(
        n115314) );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n5454), .CK(n79527), .Q(n95468), .QN(
        n115342) );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n5452), .CK(n79527), .Q(n95467), .QN(
        n115370) );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n5450), .CK(n79527), .Q(n95466), .QN(
        n115398) );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n5448), .CK(n79527), .Q(n95465), .QN(
        n115426) );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n5446), .CK(n79527), .Q(n95464), .QN(
        n115454) );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n5444), .CK(n79527), .Q(n95463), .QN(
        n115482) );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n5442), .CK(n79527), .Q(n95462), .QN(
        n115510) );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n5440), .CK(n79527), .Q(n95461), .QN(
        n115538) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n5438), .CK(n79527), .Q(n95460), .QN(
        n115566) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5436), .CK(n79527), .Q(n95459), .QN(
        n115594) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5434), .CK(n79527), .Q(n95458), .QN(
        n115622) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5432), .CK(n79527), .Q(n95457), .QN(
        n115650) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n5430), .CK(n79527), .Q(n95456), .QN(
        n115678) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n5428), .CK(n79527), .Q(n95455), .QN(
        n115706) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n5426), .CK(n79527), .Q(n95454), .QN(
        n115734) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n5424), .CK(n79527), .Q(n95453), .QN(
        n115762) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n5422), .CK(n79527), .Q(n95452), .QN(
        n115790) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n5420), .CK(n79527), .Q(n95451), .QN(
        n115818) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n5418), .CK(n79527), .Q(n95450), .QN(
        n115846) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n5416), .CK(n79527), .Q(n95449), .QN(
        n115874) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n5414), .CK(n79527), .Q(n95448), .QN(
        n115902) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n5412), .CK(n79527), .Q(n95447), .QN(
        n115930) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n5410), .CK(n79527), .Q(n95446), .QN(
        n115958) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n5408), .CK(n79527), .Q(n95445), .QN(
        n115986) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n5406), .CK(n79527), .Q(n95444), .QN(
        n116014) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n5404), .CK(n79527), .Q(n95443), .QN(
        n116042) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n5402), .CK(n79527), .Q(n95442), .QN(
        n116070) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n5400), .CK(n79527), .Q(n95441), .QN(
        n116098) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n5398), .CK(n79527), .Q(n95440), .QN(
        n116126) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n5396), .CK(n79527), .Q(n95439), .QN(
        n116154) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n5394), .CK(n79527), .Q(n95438), .QN(
        n116182) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n5392), .CK(n79527), .Q(n95437), .QN(
        n116210) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n5390), .CK(n79527), .Q(n95436), .QN(
        n116238) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n5388), .CK(n79527), .Q(n95435), .QN(
        n116266) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n5386), .CK(n79527), .Q(n95434), .QN(
        n116294) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n5384), .CK(n79527), .Q(n95433), .QN(
        n116322) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n5382), .CK(n79527), .Q(n95432), .QN(
        n116350) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n5380), .CK(n79527), .Q(n95431), .QN(
        n116378) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n5378), .CK(n79527), .Q(n95430), .QN(
        n116406) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n5376), .CK(n79527), .Q(n95429), .QN(
        n116434) );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n5562), .CK(n79527), .Q(n118084), .QN(
        n114583) );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n5561), .CK(n79527), .Q(n118083), .QN(
        n114584) );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n5560), .CK(n79527), .Q(n118082), .QN(
        n114585) );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n5559), .CK(n79527), .Q(n118081), .QN(
        n114586) );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n5558), .CK(n79527), .Q(n118080), .QN(
        n114587) );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n5557), .CK(n79527), .Q(n118079), .QN(
        n114588) );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n5556), .CK(n79527), .Q(n118078), .QN(
        n114589) );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n5555), .CK(n79527), .Q(n118077), .QN(
        n114590) );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n5554), .CK(n79527), .Q(n118076), .QN(
        n114591) );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n5553), .CK(n79527), .Q(n118075), .QN(
        n114592) );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n5552), .CK(n79527), .Q(n118074), .QN(
        n114593) );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n5551), .CK(n79527), .Q(n118073), .QN(
        n114594) );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n5550), .CK(n79527), .Q(n118072), .QN(
        n114595) );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n5549), .CK(n79527), .Q(n118071), .QN(
        n114596) );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n5548), .CK(n79527), .Q(n118070), .QN(
        n114597) );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n5547), .CK(n79527), .Q(n111040), .QN(
        n114598) );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n5546), .CK(n79527), .Q(n111039), .QN(
        n114599) );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n5545), .CK(n79527), .Q(n111038), .QN(
        n114600) );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n5544), .CK(n79527), .Q(n111037), .QN(
        n114601) );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n5543), .CK(n79527), .Q(n111036), .QN(
        n114602) );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n5542), .CK(n79527), .Q(n111035), .QN(
        n114603) );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n5541), .CK(n79527), .Q(n111034), .QN(
        n114604) );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n5540), .CK(n79527), .Q(n111033), .QN(
        n114605) );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n5539), .CK(n79527), .Q(n111032), .QN(
        n114606) );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n5538), .CK(n79527), .Q(n111031), .QN(
        n114607) );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n5537), .CK(n79527), .Q(n111030), .QN(
        n114608) );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n5536), .CK(n79527), .Q(n111029), .QN(
        n114609) );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n5535), .CK(n79527), .Q(n111028), .QN(
        n114610) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n5534), .CK(n79527), .Q(n111027), .QN(
        n114611) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5533), .CK(n79527), .Q(n111026), .QN(
        n114612) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5532), .CK(n79527), .Q(n111025), .QN(
        n114613) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5531), .CK(n79527), .Q(n111024), .QN(
        n114614) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n5530), .CK(n79527), .Q(n111023), .QN(
        n114615) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n5529), .CK(n79527), .Q(n111022), .QN(
        n114616) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n5528), .CK(n79527), .Q(n111021), .QN(
        n114617) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n5527), .CK(n79527), .Q(n111020), .QN(
        n114618) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n5526), .CK(n79527), .Q(n111019), .QN(
        n114619) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n5525), .CK(n79527), .Q(n111018), .QN(
        n114620) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n5524), .CK(n79527), .Q(n111017), .QN(
        n114621) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n5523), .CK(n79527), .Q(n111016), .QN(
        n114622) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n5522), .CK(n79527), .Q(n111015), .QN(
        n114623) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n5521), .CK(n79527), .Q(n111014), .QN(
        n114624) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n5520), .CK(n79527), .Q(n111013), .QN(
        n114625) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n5519), .CK(n79527), .Q(n111012), .QN(
        n114626) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n5518), .CK(n79527), .Q(n111011), .QN(
        n114627) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n5517), .CK(n79527), .Q(n111010), .QN(
        n114628) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n5516), .CK(n79527), .Q(n111009), .QN(
        n114629) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n5515), .CK(n79527), .Q(n111008), .QN(
        n114630) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n5514), .CK(n79527), .Q(n111007), .QN(
        n114631) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n5513), .CK(n79527), .Q(n111006), .QN(
        n114632) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n5512), .CK(n79527), .Q(n111005), .QN(
        n114633) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n5511), .CK(n79527), .Q(n111004), .QN(
        n114634) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n5510), .CK(n79527), .Q(n111003), .QN(
        n114635) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n5509), .CK(n79527), .Q(n111002), .QN(
        n114636) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n5508), .CK(n79527), .Q(n111001), .QN(
        n114637) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n5507), .CK(n79527), .Q(n111000), .QN(
        n114638) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n5506), .CK(n79527), .Q(n110999), .QN(
        n114639) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n5505), .CK(n79527), .Q(n110998), .QN(
        n114640) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n5504), .CK(n79527), .Q(n110997), .QN(
        n114641) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n5503), .CK(n79527), .Q(n110996), .QN(
        n114642) );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n5690), .CK(n79527), .QN(n114515) );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n5689), .CK(n79527), .QN(n114516) );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n5688), .CK(n79527), .QN(n114517) );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n5687), .CK(n79527), .QN(n114518) );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n5686), .CK(n79527), .QN(n114519) );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n5685), .CK(n79527), .QN(n114520) );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n5684), .CK(n79527), .QN(n114521) );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n5683), .CK(n79527), .QN(n114522) );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n5682), .CK(n79527), .QN(n114523) );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n5681), .CK(n79527), .QN(n114524) );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n5680), .CK(n79527), .QN(n114525) );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n5679), .CK(n79527), .QN(n114526) );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n5678), .CK(n79527), .QN(n114527) );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n5677), .CK(n79527), .QN(n114528) );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n5676), .CK(n79527), .QN(n114529) );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n5675), .CK(n79527), .QN(n114530) );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n5674), .CK(n79527), .QN(n114531) );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n5673), .CK(n79527), .QN(n114532) );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n5672), .CK(n79527), .QN(n114533) );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n5671), .CK(n79527), .QN(n114534) );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n5670), .CK(n79527), .QN(n114535) );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n5669), .CK(n79527), .QN(n114536) );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n5668), .CK(n79527), .QN(n114537) );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n5667), .CK(n79527), .QN(n114538) );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n5666), .CK(n79527), .QN(n114539) );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n5665), .CK(n79527), .QN(n114540) );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n5664), .CK(n79527), .QN(n114541) );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n5663), .CK(n79527), .QN(n114542) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n5662), .CK(n79527), .QN(n114543) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5661), .CK(n79527), .QN(n114544) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5660), .CK(n79527), .QN(n114545) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5659), .CK(n79527), .QN(n114546) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n5658), .CK(n79527), .QN(n114547) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n5657), .CK(n79527), .QN(n114548) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n5656), .CK(n79527), .QN(n114549) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n5655), .CK(n79527), .QN(n114550) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n5654), .CK(n79527), .QN(n114551) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n5653), .CK(n79527), .QN(n114552) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n5652), .CK(n79527), .QN(n114553) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n5651), .CK(n79527), .QN(n114554) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n5650), .CK(n79527), .QN(n114555) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n5649), .CK(n79527), .QN(n114556) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n5648), .CK(n79527), .QN(n114557) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n5647), .CK(n79527), .QN(n114558) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n5646), .CK(n79527), .QN(n114559) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n5645), .CK(n79527), .QN(n114560) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n5644), .CK(n79527), .QN(n114561) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n5643), .CK(n79527), .QN(n114562) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n5642), .CK(n79527), .QN(n114563) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n5641), .CK(n79527), .QN(n114564) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n5640), .CK(n79527), .QN(n114565) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n5639), .CK(n79527), .QN(n114566) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n5638), .CK(n79527), .QN(n114567) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n5637), .CK(n79527), .QN(n114568) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n5636), .CK(n79527), .QN(n114569) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n5635), .CK(n79527), .QN(n114570) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n5634), .CK(n79527), .QN(n114571) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n5633), .CK(n79527), .QN(n114572) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n5632), .CK(n79527), .QN(n114573) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n5631), .CK(n79527), .QN(n114574) );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n5754), .CK(n79527), .QN(n114449) );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n5753), .CK(n79527), .QN(n114450) );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n5752), .CK(n79527), .QN(n114451) );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n5751), .CK(n79527), .QN(n114452) );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n5750), .CK(n79527), .QN(n114453) );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n5749), .CK(n79527), .QN(n114454) );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n5748), .CK(n79527), .QN(n114455) );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n5747), .CK(n79527), .QN(n114456) );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n5746), .CK(n79527), .QN(n114457) );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n5745), .CK(n79527), .QN(n114458) );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n5744), .CK(n79527), .QN(n114459) );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n5743), .CK(n79527), .QN(n114460) );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n5742), .CK(n79527), .QN(n114461) );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n5741), .CK(n79527), .QN(n114462) );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n5740), .CK(n79527), .QN(n114463) );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n5739), .CK(n79527), .QN(n114464) );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n5738), .CK(n79527), .QN(n114465) );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n5737), .CK(n79527), .QN(n114466) );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n5736), .CK(n79527), .QN(n114467) );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n5735), .CK(n79527), .QN(n114468) );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n5734), .CK(n79527), .QN(n114469) );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n5733), .CK(n79527), .QN(n114470) );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n5732), .CK(n79527), .QN(n114471) );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n5731), .CK(n79527), .QN(n114472) );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n5730), .CK(n79527), .QN(n114473) );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n5729), .CK(n79527), .QN(n114474) );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n5728), .CK(n79527), .QN(n114475) );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n5727), .CK(n79527), .QN(n114476) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n5726), .CK(n79527), .QN(n114477) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5725), .CK(n79527), .QN(n114478) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5724), .CK(n79527), .QN(n114479) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5723), .CK(n79527), .QN(n114480) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n5722), .CK(n79527), .QN(n114481) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n5721), .CK(n79527), .QN(n114482) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n5720), .CK(n79527), .QN(n114483) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n5719), .CK(n79527), .QN(n114484) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n5718), .CK(n79527), .QN(n114485) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n5717), .CK(n79527), .QN(n114486) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n5716), .CK(n79527), .QN(n114487) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n5715), .CK(n79527), .QN(n114488) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n5714), .CK(n79527), .QN(n114489) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n5713), .CK(n79527), .QN(n114490) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n5712), .CK(n79527), .QN(n114491) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n5711), .CK(n79527), .QN(n114492) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n5710), .CK(n79527), .QN(n114493) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n5709), .CK(n79527), .QN(n114494) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n5708), .CK(n79527), .QN(n114495) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n5707), .CK(n79527), .QN(n114496) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n5706), .CK(n79527), .QN(n114497) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n5705), .CK(n79527), .QN(n114498) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n5704), .CK(n79527), .QN(n114499) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n5703), .CK(n79527), .QN(n114500) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n5702), .CK(n79527), .QN(n114501) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n5701), .CK(n79527), .QN(n114502) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n5700), .CK(n79527), .QN(n114503) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n5699), .CK(n79527), .QN(n114504) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n5698), .CK(n79527), .QN(n114505) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n5697), .CK(n79527), .QN(n114506) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n5696), .CK(n79527), .QN(n114507) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n5695), .CK(n79527), .QN(n114508) );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n5818), .CK(n79527), .QN(n114383) );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n5817), .CK(n79527), .QN(n114384) );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n5816), .CK(n79527), .QN(n114385) );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n5815), .CK(n79527), .QN(n114386) );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n5814), .CK(n79527), .QN(n114387) );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n5813), .CK(n79527), .QN(n114388) );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n5812), .CK(n79527), .QN(n114389) );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n5811), .CK(n79527), .QN(n114390) );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n5810), .CK(n79527), .QN(n114391) );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n5809), .CK(n79527), .QN(n114392) );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n5808), .CK(n79527), .QN(n114393) );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n5807), .CK(n79527), .QN(n114394) );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n5806), .CK(n79527), .QN(n114395) );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n5805), .CK(n79527), .QN(n114396) );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n5804), .CK(n79527), .QN(n114397) );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n5803), .CK(n79527), .QN(n114398) );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n5802), .CK(n79527), .QN(n114399) );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n5801), .CK(n79527), .QN(n114400) );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n5800), .CK(n79527), .QN(n114401) );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n5799), .CK(n79527), .QN(n114402) );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n5798), .CK(n79527), .QN(n114403) );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n5797), .CK(n79527), .QN(n114404) );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n5796), .CK(n79527), .QN(n114405) );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n5795), .CK(n79527), .QN(n114406) );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n5794), .CK(n79527), .QN(n114407) );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n5793), .CK(n79527), .QN(n114408) );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n5792), .CK(n79527), .QN(n114409) );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n5791), .CK(n79527), .QN(n114410) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n5790), .CK(n79527), .QN(n114411) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5789), .CK(n79527), .QN(n114412) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5788), .CK(n79527), .QN(n114413) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5787), .CK(n79527), .QN(n114414) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n5786), .CK(n79527), .QN(n114415) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n5785), .CK(n79527), .QN(n114416) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n5784), .CK(n79527), .QN(n114417) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n5783), .CK(n79527), .QN(n114418) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n5782), .CK(n79527), .QN(n114419) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n5781), .CK(n79527), .QN(n114420) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n5780), .CK(n79527), .QN(n114421) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n5779), .CK(n79527), .QN(n114422) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n5778), .CK(n79527), .QN(n114423) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n5777), .CK(n79527), .QN(n114424) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n5776), .CK(n79527), .QN(n114425) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n5775), .CK(n79527), .QN(n114426) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n5774), .CK(n79527), .QN(n114427) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n5773), .CK(n79527), .QN(n114428) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n5772), .CK(n79527), .QN(n114429) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n5771), .CK(n79527), .QN(n114430) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n5770), .CK(n79527), .QN(n114431) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n5769), .CK(n79527), .QN(n114432) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n5768), .CK(n79527), .QN(n114433) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n5767), .CK(n79527), .QN(n114434) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n5766), .CK(n79527), .QN(n114435) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n5765), .CK(n79527), .QN(n114436) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n5764), .CK(n79527), .QN(n114437) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n5763), .CK(n79527), .QN(n114438) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n5762), .CK(n79527), .QN(n114439) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n5761), .CK(n79527), .QN(n114440) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n5760), .CK(n79527), .QN(n114441) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n5759), .CK(n79527), .QN(n114442) );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n5946), .CK(n79527), .Q(n118444), .QN(
        n114311) );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n5945), .CK(n79527), .Q(n118443), .QN(
        n114312) );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n5944), .CK(n79527), .Q(n118442), .QN(
        n114313) );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n5943), .CK(n79527), .Q(n118441), .QN(
        n114314) );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n5942), .CK(n79527), .Q(n118440), .QN(
        n114315) );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n5941), .CK(n79527), .Q(n118439), .QN(
        n114316) );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n5940), .CK(n79527), .Q(n118438), .QN(
        n114317) );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n5939), .CK(n79527), .Q(n118437), .QN(
        n114318) );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n5938), .CK(n79527), .Q(n118436), .QN(
        n114319) );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n5937), .CK(n79527), .Q(n118435), .QN(
        n114320) );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n5936), .CK(n79527), .Q(n118434), .QN(
        n114321) );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n5935), .CK(n79527), .Q(n118433), .QN(
        n114322) );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n5934), .CK(n79527), .Q(n118432), .QN(
        n114323) );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n5933), .CK(n79527), .Q(n118431), .QN(
        n114324) );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n5932), .CK(n79527), .Q(n118430), .QN(
        n114325) );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n5931), .CK(n79527), .Q(n118429), .QN(
        n114326) );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n5930), .CK(n79527), .Q(n118428), .QN(
        n114327) );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n5929), .CK(n79527), .Q(n118427), .QN(
        n114328) );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n5928), .CK(n79527), .Q(n118426), .QN(
        n114329) );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n5927), .CK(n79527), .Q(n118425), .QN(
        n114330) );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n5926), .CK(n79527), .Q(n118424), .QN(
        n114331) );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n5925), .CK(n79527), .Q(n118423), .QN(
        n114332) );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n5924), .CK(n79527), .Q(n118422), .QN(
        n114333) );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n5923), .CK(n79527), .Q(n118421), .QN(
        n114334) );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n5922), .CK(n79527), .Q(n118420), .QN(
        n114335) );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n5921), .CK(n79527), .Q(n118419), .QN(
        n114336) );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n5920), .CK(n79527), .Q(n118418), .QN(
        n114337) );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n5919), .CK(n79527), .Q(n118417), .QN(
        n114338) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5918), .CK(n79527), .Q(n118416), .QN(
        n114339) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5917), .CK(n79527), .Q(n118415), .QN(
        n114340) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5916), .CK(n79527), .Q(n118414), .QN(
        n114341) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5915), .CK(n79527), .Q(n118413), .QN(
        n114342) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n5914), .CK(n79527), .Q(n118412), .QN(
        n114343) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n5913), .CK(n79527), .Q(n118411), .QN(
        n114344) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n5912), .CK(n79527), .Q(n118410), .QN(
        n114345) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n5911), .CK(n79527), .Q(n118409), .QN(
        n114346) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n5910), .CK(n79527), .Q(n118408), .QN(
        n114347) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n5909), .CK(n79527), .Q(n118407), .QN(
        n114348) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n5908), .CK(n79527), .Q(n118406), .QN(
        n114349) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n5907), .CK(n79527), .Q(n118405), .QN(
        n114350) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n5906), .CK(n79527), .Q(n118404), .QN(
        n114351) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n5905), .CK(n79527), .Q(n118403), .QN(
        n114352) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n5904), .CK(n79527), .Q(n118402), .QN(
        n114353) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n5903), .CK(n79527), .Q(n118401), .QN(
        n114354) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n5902), .CK(n79527), .Q(n118400), .QN(
        n114355) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n5901), .CK(n79527), .Q(n118399), .QN(
        n114356) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n5900), .CK(n79527), .Q(n118398), .QN(
        n114357) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n5899), .CK(n79527), .Q(n118397), .QN(
        n114358) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n5898), .CK(n79527), .Q(n118396), .QN(
        n114359) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n5897), .CK(n79527), .Q(n118395), .QN(
        n114360) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n5896), .CK(n79527), .Q(n118394), .QN(
        n114361) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n5895), .CK(n79527), .Q(n118393), .QN(
        n114362) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n5894), .CK(n79527), .Q(n118392), .QN(
        n114363) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n5893), .CK(n79527), .Q(n118391), .QN(
        n114364) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n5892), .CK(n79527), .Q(n118390), .QN(
        n114365) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n5891), .CK(n79527), .Q(n118389), .QN(
        n114366) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n5890), .CK(n79527), .Q(n118388), .QN(
        n114367) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n5889), .CK(n79527), .Q(n118387), .QN(
        n114368) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n5888), .CK(n79527), .Q(n118386), .QN(
        n114369) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n5887), .CK(n79527), .Q(n118385), .QN(
        n114370) );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n6138), .CK(n79527), .Q(n118384), .QN(
        n114240) );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n6137), .CK(n79527), .Q(n118383), .QN(
        n114241) );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n6136), .CK(n79527), .Q(n118382), .QN(
        n114242) );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n6135), .CK(n79527), .Q(n118381), .QN(
        n114243) );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n6134), .CK(n79527), .Q(n118380), .QN(
        n114244) );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n6133), .CK(n79527), .Q(n118379), .QN(
        n114245) );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n6132), .CK(n79527), .Q(n118378), .QN(
        n114246) );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n6131), .CK(n79527), .Q(n118377), .QN(
        n114247) );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n6130), .CK(n79527), .Q(n118376), .QN(
        n114248) );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n6129), .CK(n79527), .Q(n118375), .QN(
        n114249) );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n6128), .CK(n79527), .Q(n118374), .QN(
        n114250) );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n6127), .CK(n79527), .Q(n118373), .QN(
        n114251) );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n6126), .CK(n79527), .Q(n118372), .QN(
        n114252) );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n6125), .CK(n79527), .Q(n118371), .QN(
        n114253) );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n6124), .CK(n79527), .Q(n118370), .QN(
        n114254) );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n6123), .CK(n79527), .Q(n118369), .QN(
        n114255) );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n6122), .CK(n79527), .Q(n118368), .QN(
        n114256) );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n6121), .CK(n79527), .Q(n118367), .QN(
        n114257) );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n6120), .CK(n79527), .Q(n118366), .QN(
        n114258) );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n6119), .CK(n79527), .Q(n118365), .QN(
        n114259) );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n6118), .CK(n79527), .Q(n118364), .QN(
        n114260) );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n6117), .CK(n79527), .Q(n118363), .QN(
        n114261) );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n6116), .CK(n79527), .Q(n118362), .QN(
        n114262) );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n6115), .CK(n79527), .Q(n118361), .QN(
        n114263) );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n6114), .CK(n79527), .Q(n118360), .QN(
        n114264) );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n6113), .CK(n79527), .Q(n118359), .QN(
        n114265) );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n6112), .CK(n79527), .Q(n118358), .QN(
        n114266) );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n6111), .CK(n79527), .Q(n118357), .QN(
        n114267) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n6110), .CK(n79527), .Q(n118356), .QN(
        n114268) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n6109), .CK(n79527), .Q(n118355), .QN(
        n114269) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n6108), .CK(n79527), .Q(n118354), .QN(
        n114270) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n6107), .CK(n79527), .Q(n118353), .QN(
        n114271) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n6106), .CK(n79527), .Q(n118352), .QN(
        n114272) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n6105), .CK(n79527), .Q(n118351), .QN(
        n114273) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n6104), .CK(n79527), .Q(n118350), .QN(
        n114274) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n6103), .CK(n79527), .Q(n118349), .QN(
        n114275) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n6102), .CK(n79527), .Q(n118348), .QN(
        n114276) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n6101), .CK(n79527), .Q(n118347), .QN(
        n114277) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n6100), .CK(n79527), .Q(n118346), .QN(
        n114278) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n6099), .CK(n79527), .Q(n118345), .QN(
        n114279) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n6098), .CK(n79527), .Q(n118344), .QN(
        n114280) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n6097), .CK(n79527), .Q(n118343), .QN(
        n114281) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n6096), .CK(n79527), .Q(n118342), .QN(
        n114282) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n6095), .CK(n79527), .Q(n118341), .QN(
        n114283) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n6094), .CK(n79527), .Q(n118340), .QN(
        n114284) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n6093), .CK(n79527), .Q(n118339), .QN(
        n114285) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n6092), .CK(n79527), .Q(n118338), .QN(
        n114286) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n6091), .CK(n79527), .Q(n118337), .QN(
        n114287) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n6090), .CK(n79527), .Q(n118336), .QN(
        n114288) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n6089), .CK(n79527), .Q(n118335), .QN(
        n114289) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n6088), .CK(n79527), .Q(n118334), .QN(
        n114290) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n6087), .CK(n79527), .Q(n118333), .QN(
        n114291) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n6086), .CK(n79527), .Q(n118332), .QN(
        n114292) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n6085), .CK(n79527), .Q(n118331), .QN(
        n114293) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n6084), .CK(n79527), .Q(n118330), .QN(
        n114294) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n6083), .CK(n79527), .Q(n118329), .QN(
        n114295) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n6082), .CK(n79527), .Q(n118328), .QN(
        n114296) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n6081), .CK(n79527), .Q(n118327), .QN(
        n114297) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n6080), .CK(n79527), .Q(n118326), .QN(
        n114298) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n6079), .CK(n79527), .Q(n118325), .QN(
        n114299) );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n6330), .CK(n79527), .QN(n114151) );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n6329), .CK(n79527), .QN(n114152) );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n6328), .CK(n79527), .QN(n114153) );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n6327), .CK(n79527), .QN(n114154) );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n6326), .CK(n79527), .QN(n114155) );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n6325), .CK(n79527), .QN(n114156) );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n6324), .CK(n79527), .QN(n114157) );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n6323), .CK(n79527), .QN(n114158) );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n6322), .CK(n79527), .QN(n114159) );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n6321), .CK(n79527), .QN(n114160) );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n6320), .CK(n79527), .QN(n114161) );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n6319), .CK(n79527), .QN(n114162) );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n6318), .CK(n79527), .QN(n114163) );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n6317), .CK(n79527), .QN(n114164) );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n6316), .CK(n79527), .QN(n114165) );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n6315), .CK(n79527), .QN(n114166) );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n6314), .CK(n79527), .QN(n114167) );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n6313), .CK(n79527), .QN(n114168) );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n6312), .CK(n79527), .QN(n114169) );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n6311), .CK(n79527), .QN(n114170) );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n6310), .CK(n79527), .QN(n114171) );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n6309), .CK(n79527), .QN(n114172) );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n6308), .CK(n79527), .QN(n114173) );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n6307), .CK(n79527), .QN(n114174) );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n6306), .CK(n79527), .QN(n114175) );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n6305), .CK(n79527), .QN(n114176) );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n6304), .CK(n79527), .QN(n114177) );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n6303), .CK(n79527), .QN(n114178) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n6302), .CK(n79527), .QN(n114179) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n6301), .CK(n79527), .QN(n114180) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n6300), .CK(n79527), .QN(n114181) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n6299), .CK(n79527), .QN(n114182) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n6298), .CK(n79527), .QN(n114183) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n6297), .CK(n79527), .QN(n114184) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n6296), .CK(n79527), .QN(n114185) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n6295), .CK(n79527), .QN(n114186) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n6294), .CK(n79527), .QN(n114187) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n6293), .CK(n79527), .QN(n114188) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n6292), .CK(n79527), .QN(n114189) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n6291), .CK(n79527), .QN(n114190) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n6290), .CK(n79527), .QN(n114191) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n6289), .CK(n79527), .QN(n114192) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n6288), .CK(n79527), .QN(n114193) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n6287), .CK(n79527), .QN(n114194) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n6286), .CK(n79527), .QN(n114195) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n6285), .CK(n79527), .QN(n114196) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n6284), .CK(n79527), .QN(n114197) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n6283), .CK(n79527), .QN(n114198) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n6282), .CK(n79527), .QN(n114199) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n6281), .CK(n79527), .QN(n114200) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n6280), .CK(n79527), .QN(n114201) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n6279), .CK(n79527), .QN(n114202) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n6278), .CK(n79527), .QN(n114203) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n6277), .CK(n79527), .QN(n114204) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n6276), .CK(n79527), .QN(n114205) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n6275), .CK(n79527), .QN(n114206) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n6274), .CK(n79527), .QN(n114207) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n6273), .CK(n79527), .QN(n114208) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n6272), .CK(n79527), .QN(n114209) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n6271), .CK(n79527), .QN(n114210) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n6910), .CK(n79527), .Q(n117977), .QN(
        n114056) );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n6909), .CK(n79527), .Q(n117976), .QN(
        n114058) );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n6908), .CK(n79527), .Q(n117975), .QN(
        n114059) );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n6907), .CK(n79527), .Q(n117974), .QN(
        n114060) );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n7482), .CK(n79527), .QN(n113772) );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n7481), .CK(n79527), .QN(n113774) );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n7480), .CK(n79527), .QN(n113776) );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n7479), .CK(n79527), .QN(n113778) );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n7478), .CK(n79527), .QN(n113780) );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n7477), .CK(n79527), .QN(n113782) );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n7476), .CK(n79527), .QN(n113784) );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n7475), .CK(n79527), .QN(n113786) );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n7474), .CK(n79527), .QN(n113788) );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n7473), .CK(n79527), .QN(n113790) );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n7472), .CK(n79527), .QN(n113792) );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n7471), .CK(n79527), .QN(n113794) );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n7470), .CK(n79527), .QN(n113796) );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n7469), .CK(n79527), .QN(n113798) );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n7468), .CK(n79527), .QN(n113800) );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n7467), .CK(n79527), .QN(n113802) );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n7466), .CK(n79527), .QN(n113804) );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n7465), .CK(n79527), .QN(n113806) );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n7464), .CK(n79527), .QN(n113808) );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n7463), .CK(n79527), .QN(n113810) );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n7462), .CK(n79527), .QN(n113812) );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n7461), .CK(n79527), .QN(n113814) );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n7460), .CK(n79527), .QN(n113816) );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n7459), .CK(n79527), .QN(n113818) );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n7458), .CK(n79527), .QN(n113820) );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n7457), .CK(n79527), .QN(n113822) );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n7456), .CK(n79527), .QN(n113824) );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n7455), .CK(n79527), .QN(n113826) );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n7454), .CK(n79527), .QN(n113828) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n7453), .CK(n79527), .QN(n113830) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n7452), .CK(n79527), .QN(n113832) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n7451), .CK(n79527), .QN(n113834) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n7450), .CK(n79527), .QN(n113836) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n7449), .CK(n79527), .QN(n113838) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n7448), .CK(n79527), .QN(n113840) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n7447), .CK(n79527), .QN(n113842) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n7446), .CK(n79527), .QN(n113844) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n7445), .CK(n79527), .QN(n113846) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n7444), .CK(n79527), .QN(n113848) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n7443), .CK(n79527), .QN(n113850) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n7442), .CK(n79527), .QN(n113852) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n7441), .CK(n79527), .QN(n113854) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n7440), .CK(n79527), .QN(n113856) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n7439), .CK(n79527), .QN(n113858) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n7438), .CK(n79527), .QN(n113860) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n7437), .CK(n79527), .QN(n113862) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n7436), .CK(n79527), .QN(n113864) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n7435), .CK(n79527), .QN(n113866) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n7434), .CK(n79527), .QN(n113868) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n7433), .CK(n79527), .QN(n113870) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n7432), .CK(n79527), .QN(n113872) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n7431), .CK(n79527), .QN(n113874) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n7430), .CK(n79527), .QN(n113876) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n7429), .CK(n79527), .QN(n113878) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n7428), .CK(n79527), .QN(n113880) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n7427), .CK(n79527), .QN(n113882) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n7426), .CK(n79527), .QN(n113884) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n7425), .CK(n79527), .QN(n113886) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n7424), .CK(n79527), .QN(n113888) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n7423), .CK(n79527), .QN(n113890) );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n7034), .CK(n79527), .QN(n113992) );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n7033), .CK(n79527), .QN(n113993) );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n7032), .CK(n79527), .QN(n113994) );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n7031), .CK(n79527), .QN(n113995) );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n7030), .CK(n79527), .QN(n113996) );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n7029), .CK(n79527), .QN(n113997) );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n7028), .CK(n79527), .QN(n113998) );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n7027), .CK(n79527), .QN(n113999) );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n7026), .CK(n79527), .QN(n114000) );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n7025), .CK(n79527), .QN(n114001) );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n7024), .CK(n79527), .QN(n114002) );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n7023), .CK(n79527), .QN(n114003) );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n7022), .CK(n79527), .QN(n114004) );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n7021), .CK(n79527), .QN(n114005) );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n7020), .CK(n79527), .QN(n114006) );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n7019), .CK(n79527), .QN(n114007) );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n7018), .CK(n79527), .QN(n114008) );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n7017), .CK(n79527), .QN(n114009) );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n7016), .CK(n79527), .QN(n114010) );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n7015), .CK(n79527), .QN(n114011) );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n7014), .CK(n79527), .QN(n114012) );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n7013), .CK(n79527), .QN(n114013) );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n7012), .CK(n79527), .QN(n114014) );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n7011), .CK(n79527), .QN(n114015) );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n7010), .CK(n79527), .QN(n114016) );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n7009), .CK(n79527), .QN(n114017) );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n7008), .CK(n79527), .QN(n114018) );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n7007), .CK(n79527), .QN(n114019) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n7006), .CK(n79527), .QN(n114020) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n7005), .CK(n79527), .QN(n114021) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n7004), .CK(n79527), .QN(n114022) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n7003), .CK(n79527), .QN(n114023) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n7002), .CK(n79527), .QN(n114024) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n7001), .CK(n79527), .QN(n114025) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n7000), .CK(n79527), .QN(n114026) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n6999), .CK(n79527), .QN(n114027) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n6998), .CK(n79527), .QN(n114028) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n6997), .CK(n79527), .QN(n114029) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n6996), .CK(n79527), .QN(n114030) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n6995), .CK(n79527), .QN(n114031) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n6994), .CK(n79527), .QN(n114032) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n6993), .CK(n79527), .QN(n114033) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n6992), .CK(n79527), .QN(n114034) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n6991), .CK(n79527), .QN(n114035) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n6990), .CK(n79527), .QN(n114036) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n6989), .CK(n79527), .QN(n114037) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n6988), .CK(n79527), .QN(n114038) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n6987), .CK(n79527), .QN(n114039) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n6986), .CK(n79527), .QN(n114040) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n6985), .CK(n79527), .QN(n114041) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n6984), .CK(n79527), .QN(n114042) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n6983), .CK(n79527), .QN(n114043) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n6982), .CK(n79527), .QN(n114044) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n6981), .CK(n79527), .QN(n114045) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n6980), .CK(n79527), .QN(n114046) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n6979), .CK(n79527), .QN(n114047) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n6978), .CK(n79527), .QN(n114048) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n6977), .CK(n79527), .QN(n114049) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n6976), .CK(n79527), .QN(n114050) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n6975), .CK(n79527), .QN(n114051) );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n7162), .CK(n79527), .QN(n113920) );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n7161), .CK(n79527), .QN(n113921) );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n7160), .CK(n79527), .QN(n113922) );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n7159), .CK(n79527), .QN(n113923) );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n7158), .CK(n79527), .QN(n113924) );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n7157), .CK(n79527), .QN(n113925) );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n7156), .CK(n79527), .QN(n113926) );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n7155), .CK(n79527), .QN(n113927) );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n7154), .CK(n79527), .QN(n113928) );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n7153), .CK(n79527), .QN(n113929) );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n7152), .CK(n79527), .QN(n113930) );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n7151), .CK(n79527), .QN(n113931) );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n7150), .CK(n79527), .QN(n113932) );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n7149), .CK(n79527), .QN(n113933) );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n7148), .CK(n79527), .QN(n113934) );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n7147), .CK(n79527), .QN(n113935) );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n7146), .CK(n79527), .QN(n113936) );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n7145), .CK(n79527), .QN(n113937) );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n7144), .CK(n79527), .QN(n113938) );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n7143), .CK(n79527), .QN(n113939) );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n7142), .CK(n79527), .QN(n113940) );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n7141), .CK(n79527), .QN(n113941) );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n7140), .CK(n79527), .QN(n113942) );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n7139), .CK(n79527), .QN(n113943) );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n7138), .CK(n79527), .QN(n113944) );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n7137), .CK(n79527), .QN(n113945) );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n7136), .CK(n79527), .QN(n113946) );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n7135), .CK(n79527), .QN(n113947) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n7134), .CK(n79527), .QN(n113948) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n7133), .CK(n79527), .QN(n113949) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n7132), .CK(n79527), .QN(n113950) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n7131), .CK(n79527), .QN(n113951) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n7130), .CK(n79527), .QN(n113952) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n7129), .CK(n79527), .QN(n113953) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n7128), .CK(n79527), .QN(n113954) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n7127), .CK(n79527), .QN(n113955) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n7126), .CK(n79527), .QN(n113956) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n7125), .CK(n79527), .QN(n113957) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n7124), .CK(n79527), .QN(n113958) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n7123), .CK(n79527), .QN(n113959) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n7122), .CK(n79527), .QN(n113960) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n7121), .CK(n79527), .QN(n113961) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n7120), .CK(n79527), .QN(n113962) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n7119), .CK(n79527), .QN(n113963) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n7118), .CK(n79527), .QN(n113964) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n7117), .CK(n79527), .QN(n113965) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n7116), .CK(n79527), .QN(n113966) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n7115), .CK(n79527), .QN(n113967) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n7114), .CK(n79527), .QN(n113968) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n7113), .CK(n79527), .QN(n113969) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n7112), .CK(n79527), .QN(n113970) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n7111), .CK(n79527), .QN(n113971) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n7110), .CK(n79527), .QN(n113972) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n7109), .CK(n79527), .QN(n113973) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n7108), .CK(n79527), .QN(n113974) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n7107), .CK(n79527), .QN(n113975) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n7106), .CK(n79527), .QN(n113976) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n7105), .CK(n79527), .QN(n113977) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n7104), .CK(n79527), .QN(n113978) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n7103), .CK(n79527), .QN(n113979) );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n6906), .CK(n79527), .Q(n118264), .QN(
        n114061) );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n6905), .CK(n79527), .Q(n118263), .QN(
        n114062) );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n6904), .CK(n79527), .Q(n118262), .QN(
        n114063) );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n6903), .CK(n79527), .Q(n118261), .QN(
        n114064) );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n6902), .CK(n79527), .Q(n118260), .QN(
        n114065) );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n6901), .CK(n79527), .Q(n118259), .QN(
        n114066) );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n6900), .CK(n79527), .Q(n118258), .QN(
        n114067) );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n6899), .CK(n79527), .Q(n118257), .QN(
        n114068) );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n6898), .CK(n79527), .Q(n118256), .QN(
        n114069) );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n6897), .CK(n79527), .Q(n118255), .QN(
        n114070) );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n6896), .CK(n79527), .Q(n118254), .QN(
        n114071) );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n6895), .CK(n79527), .Q(n118253), .QN(
        n114072) );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n6894), .CK(n79527), .Q(n118252), .QN(
        n114073) );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n6893), .CK(n79527), .Q(n118251), .QN(
        n114074) );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n6892), .CK(n79527), .Q(n118250), .QN(
        n114075) );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n6891), .CK(n79527), .Q(n118249), .QN(
        n114076) );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n6890), .CK(n79527), .Q(n118248), .QN(
        n114077) );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n6889), .CK(n79527), .Q(n118247), .QN(
        n114078) );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n6888), .CK(n79527), .Q(n118246), .QN(
        n114079) );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n6887), .CK(n79527), .Q(n118245), .QN(
        n114080) );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n6886), .CK(n79527), .Q(n118244), .QN(
        n114081) );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n6885), .CK(n79527), .Q(n118243), .QN(
        n114082) );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n6884), .CK(n79527), .Q(n118242), .QN(
        n114083) );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n6883), .CK(n79527), .Q(n118241), .QN(
        n114084) );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n6882), .CK(n79527), .Q(n118240), .QN(
        n114085) );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n6881), .CK(n79527), .Q(n118239), .QN(
        n114086) );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n6880), .CK(n79527), .Q(n118238), .QN(
        n114087) );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n6879), .CK(n79527), .Q(n118237), .QN(
        n114088) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n6878), .CK(n79527), .Q(n118236), .QN(
        n114089) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n6877), .CK(n79527), .Q(n118235), .QN(
        n114090) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n6876), .CK(n79527), .Q(n118234), .QN(
        n114091) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n6875), .CK(n79527), .Q(n118233), .QN(
        n114092) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n6874), .CK(n79527), .Q(n118232), .QN(
        n114093) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n6873), .CK(n79527), .Q(n118231), .QN(
        n114094) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n6872), .CK(n79527), .Q(n118230), .QN(
        n114095) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n6871), .CK(n79527), .Q(n118229), .QN(
        n114096) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n6870), .CK(n79527), .Q(n118228), .QN(
        n114097) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n6869), .CK(n79527), .Q(n118227), .QN(
        n114098) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n6868), .CK(n79527), .Q(n118226), .QN(
        n114099) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n6867), .CK(n79527), .Q(n118225), .QN(
        n114100) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n6866), .CK(n79527), .Q(n118224), .QN(
        n114101) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n6865), .CK(n79527), .Q(n118223), .QN(
        n114102) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n6864), .CK(n79527), .Q(n118222), .QN(
        n114103) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n6863), .CK(n79527), .Q(n118221), .QN(
        n114104) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n6862), .CK(n79527), .Q(n118220), .QN(
        n114105) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n6861), .CK(n79527), .Q(n118219), .QN(
        n114106) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n6860), .CK(n79527), .Q(n118218), .QN(
        n114107) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n6859), .CK(n79527), .Q(n118217), .QN(
        n114108) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n6858), .CK(n79527), .Q(n118216), .QN(
        n114109) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n6857), .CK(n79527), .Q(n118215), .QN(
        n114110) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n6856), .CK(n79527), .Q(n118214), .QN(
        n114111) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n6855), .CK(n79527), .Q(n118213), .QN(
        n114112) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n6854), .CK(n79527), .Q(n118212), .QN(
        n114113) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n6853), .CK(n79527), .Q(n118211), .QN(
        n114114) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n6852), .CK(n79527), .Q(n118210), .QN(
        n114115) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n6851), .CK(n79527), .Q(n118209), .QN(
        n114116) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n6850), .CK(n79527), .Q(n118208), .QN(
        n114117) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n6849), .CK(n79527), .Q(n118207), .QN(
        n114118) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n6848), .CK(n79527), .Q(n118206), .QN(
        n114119) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n6847), .CK(n79527), .Q(n118205), .QN(
        n114120) );
  DFF_X1 \OUT1_reg[63]  ( .D(n5501), .CK(n79527), .Q(OUT1[63]) );
  DFF_X1 \OUT1_reg[62]  ( .D(n5499), .CK(n79527), .Q(OUT1[62]) );
  DFF_X1 \OUT1_reg[61]  ( .D(n5497), .CK(n79527), .Q(OUT1[61]) );
  DFF_X1 \OUT1_reg[60]  ( .D(n5495), .CK(n79527), .Q(OUT1[60]) );
  DFF_X1 \OUT2_reg[63]  ( .D(n5374), .CK(n79527), .Q(OUT2[63]) );
  DFF_X1 \OUT2_reg[62]  ( .D(n5373), .CK(n79527), .Q(OUT2[62]) );
  DFF_X1 \OUT2_reg[61]  ( .D(n5372), .CK(n79527), .Q(OUT2[61]) );
  DFF_X1 \OUT2_reg[60]  ( .D(n5371), .CK(n79527), .Q(OUT2[60]) );
  DFF_X1 \OUT2_reg[59]  ( .D(n5370), .CK(n79527), .Q(OUT2[59]) );
  DFF_X1 \OUT2_reg[58]  ( .D(n5369), .CK(n79527), .Q(OUT2[58]) );
  DFF_X1 \OUT2_reg[57]  ( .D(n5368), .CK(n79527), .Q(OUT2[57]) );
  DFF_X1 \OUT2_reg[56]  ( .D(n5367), .CK(n79527), .Q(OUT2[56]) );
  DFF_X1 \OUT2_reg[55]  ( .D(n5366), .CK(n79527), .Q(OUT2[55]) );
  DFF_X1 \OUT2_reg[54]  ( .D(n5365), .CK(n79527), .Q(OUT2[54]) );
  DFF_X1 \OUT2_reg[53]  ( .D(n5364), .CK(n79527), .Q(OUT2[53]) );
  DFF_X1 \OUT2_reg[52]  ( .D(n5363), .CK(n79527), .Q(OUT2[52]) );
  DFF_X1 \OUT2_reg[51]  ( .D(n5362), .CK(n79527), .Q(OUT2[51]) );
  DFF_X1 \OUT2_reg[50]  ( .D(n5361), .CK(n79527), .Q(OUT2[50]) );
  DFF_X1 \OUT2_reg[49]  ( .D(n5360), .CK(n79527), .Q(OUT2[49]) );
  DFF_X1 \OUT2_reg[48]  ( .D(n5359), .CK(n79527), .Q(OUT2[48]) );
  DFF_X1 \OUT2_reg[47]  ( .D(n5358), .CK(n79527), .Q(OUT2[47]) );
  DFF_X1 \OUT2_reg[46]  ( .D(n5357), .CK(n79527), .Q(OUT2[46]) );
  DFF_X1 \OUT2_reg[45]  ( .D(n5356), .CK(n79527), .Q(OUT2[45]) );
  DFF_X1 \OUT2_reg[44]  ( .D(n5355), .CK(n79527), .Q(OUT2[44]) );
  DFF_X1 \OUT2_reg[43]  ( .D(n5354), .CK(n79527), .Q(OUT2[43]) );
  DFF_X1 \OUT2_reg[42]  ( .D(n5353), .CK(n79527), .Q(OUT2[42]) );
  DFF_X1 \OUT2_reg[41]  ( .D(n5352), .CK(n79527), .Q(OUT2[41]) );
  DFF_X1 \OUT2_reg[40]  ( .D(n5351), .CK(n79527), .Q(OUT2[40]) );
  DFF_X1 \OUT2_reg[39]  ( .D(n5350), .CK(n79527), .Q(OUT2[39]) );
  DFF_X1 \OUT2_reg[38]  ( .D(n5349), .CK(n79527), .Q(OUT2[38]) );
  DFF_X1 \OUT2_reg[37]  ( .D(n5348), .CK(n79527), .Q(OUT2[37]) );
  DFF_X1 \OUT2_reg[36]  ( .D(n5347), .CK(n79527), .Q(OUT2[36]) );
  DFF_X1 \OUT2_reg[35]  ( .D(n5346), .CK(n79527), .Q(OUT2[35]) );
  DFF_X1 \OUT2_reg[34]  ( .D(n5345), .CK(n79527), .Q(OUT2[34]) );
  DFF_X1 \OUT2_reg[33]  ( .D(n5344), .CK(n79527), .Q(OUT2[33]) );
  DFF_X1 \OUT2_reg[32]  ( .D(n5343), .CK(n79527), .Q(OUT2[32]) );
  DFF_X1 \OUT2_reg[31]  ( .D(n5342), .CK(n79527), .Q(OUT2[31]) );
  DFF_X1 \OUT2_reg[30]  ( .D(n5341), .CK(n79527), .Q(OUT2[30]) );
  NOR3_X1 U83326 ( .A1(n120018), .A2(ADD_RD2[2]), .A3(n117973), .ZN(n117945)
         );
  NOR3_X1 U83327 ( .A1(n120018), .A2(ADD_RD2[1]), .A3(n117971), .ZN(n117953)
         );
  NOR3_X1 U83328 ( .A1(n117971), .A2(n120018), .A3(n117973), .ZN(n117948) );
  NOR3_X1 U83329 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n120018), .ZN(n117954) );
  NOR3_X1 U83330 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n120216), .ZN(n116445) );
  BUF_X1 U83331 ( .A(n120827), .Z(n120829) );
  BUF_X1 U83332 ( .A(n120828), .Z(n120833) );
  BUF_X1 U83333 ( .A(n120828), .Z(n120832) );
  BUF_X1 U83334 ( .A(n120827), .Z(n120831) );
  BUF_X1 U83335 ( .A(n120827), .Z(n120830) );
  BUF_X1 U83336 ( .A(n116528), .Z(n119863) );
  BUF_X1 U83337 ( .A(n116528), .Z(n119864) );
  BUF_X1 U83338 ( .A(n116528), .Z(n119865) );
  BUF_X1 U83339 ( .A(n116528), .Z(n119866) );
  BUF_X1 U83340 ( .A(n116528), .Z(n119862) );
  BUF_X1 U83341 ( .A(n113767), .Z(n120822) );
  BUF_X1 U83342 ( .A(n113767), .Z(n120823) );
  BUF_X1 U83343 ( .A(n113767), .Z(n120824) );
  BUF_X1 U83344 ( .A(n113767), .Z(n120825) );
  BUF_X1 U83345 ( .A(n120543), .Z(n120545) );
  BUF_X1 U83346 ( .A(n120246), .Z(n120248) );
  BUF_X1 U83347 ( .A(n120259), .Z(n120261) );
  BUF_X1 U83348 ( .A(n120518), .Z(n120520) );
  BUF_X1 U83349 ( .A(n120568), .Z(n120570) );
  BUF_X1 U83350 ( .A(n120372), .Z(n120374) );
  BUF_X1 U83351 ( .A(n120335), .Z(n120337) );
  BUF_X1 U83352 ( .A(n120284), .Z(n120286) );
  BUF_X1 U83353 ( .A(n120409), .Z(n120411) );
  BUF_X1 U83354 ( .A(n120310), .Z(n120312) );
  BUF_X1 U83355 ( .A(n120297), .Z(n120299) );
  BUF_X1 U83356 ( .A(n120544), .Z(n120549) );
  BUF_X1 U83357 ( .A(n120544), .Z(n120548) );
  BUF_X1 U83358 ( .A(n120543), .Z(n120547) );
  BUF_X1 U83359 ( .A(n120543), .Z(n120546) );
  BUF_X1 U83360 ( .A(n120246), .Z(n120249) );
  BUF_X1 U83361 ( .A(n120246), .Z(n120250) );
  BUF_X1 U83362 ( .A(n120247), .Z(n120251) );
  BUF_X1 U83363 ( .A(n120259), .Z(n120262) );
  BUF_X1 U83364 ( .A(n120259), .Z(n120263) );
  BUF_X1 U83365 ( .A(n120247), .Z(n120252) );
  BUF_X1 U83366 ( .A(n120518), .Z(n120521) );
  BUF_X1 U83367 ( .A(n120518), .Z(n120522) );
  BUF_X1 U83368 ( .A(n120519), .Z(n120523) );
  BUF_X1 U83369 ( .A(n120568), .Z(n120571) );
  BUF_X1 U83370 ( .A(n120568), .Z(n120572) );
  BUF_X1 U83371 ( .A(n120569), .Z(n120573) );
  BUF_X1 U83372 ( .A(n120519), .Z(n120524) );
  BUF_X1 U83373 ( .A(n120372), .Z(n120375) );
  BUF_X1 U83374 ( .A(n120372), .Z(n120376) );
  BUF_X1 U83375 ( .A(n120373), .Z(n120377) );
  BUF_X1 U83376 ( .A(n120335), .Z(n120338) );
  BUF_X1 U83377 ( .A(n120335), .Z(n120339) );
  BUF_X1 U83378 ( .A(n120336), .Z(n120340) );
  BUF_X1 U83379 ( .A(n120284), .Z(n120287) );
  BUF_X1 U83380 ( .A(n120284), .Z(n120288) );
  BUF_X1 U83381 ( .A(n120285), .Z(n120289) );
  BUF_X1 U83382 ( .A(n120260), .Z(n120264) );
  BUF_X1 U83383 ( .A(n120409), .Z(n120412) );
  BUF_X1 U83384 ( .A(n120409), .Z(n120413) );
  BUF_X1 U83385 ( .A(n120410), .Z(n120414) );
  BUF_X1 U83386 ( .A(n120310), .Z(n120313) );
  BUF_X1 U83387 ( .A(n120310), .Z(n120314) );
  BUF_X1 U83388 ( .A(n120311), .Z(n120315) );
  BUF_X1 U83389 ( .A(n120569), .Z(n120574) );
  BUF_X1 U83390 ( .A(n120373), .Z(n120378) );
  BUF_X1 U83391 ( .A(n120336), .Z(n120341) );
  BUF_X1 U83392 ( .A(n120285), .Z(n120290) );
  BUF_X1 U83393 ( .A(n120260), .Z(n120265) );
  BUF_X1 U83394 ( .A(n120297), .Z(n120300) );
  BUF_X1 U83395 ( .A(n120297), .Z(n120301) );
  BUF_X1 U83396 ( .A(n120298), .Z(n120302) );
  BUF_X1 U83397 ( .A(n120410), .Z(n120415) );
  BUF_X1 U83398 ( .A(n120298), .Z(n120303) );
  BUF_X1 U83399 ( .A(n120311), .Z(n120316) );
  BUF_X1 U83400 ( .A(n114139), .Z(n120434) );
  BUF_X1 U83401 ( .A(n114139), .Z(n120435) );
  BUF_X1 U83402 ( .A(n114139), .Z(n120436) );
  BUF_X1 U83403 ( .A(n114139), .Z(n120437) );
  BUF_X1 U83404 ( .A(n114139), .Z(n120438) );
  BUF_X1 U83405 ( .A(n114645), .Z(n120240) );
  BUF_X1 U83406 ( .A(n114645), .Z(n120241) );
  BUF_X1 U83407 ( .A(n114645), .Z(n120242) );
  BUF_X1 U83408 ( .A(n114645), .Z(n120243) );
  BUF_X1 U83409 ( .A(n114645), .Z(n120244) );
  BUF_X1 U83410 ( .A(n113897), .Z(n120611) );
  BUF_X1 U83411 ( .A(n113897), .Z(n120612) );
  BUF_X1 U83412 ( .A(n113897), .Z(n120613) );
  BUF_X1 U83413 ( .A(n113897), .Z(n120614) );
  BUF_X1 U83414 ( .A(n113897), .Z(n120615) );
  BUF_X1 U83415 ( .A(n113904), .Z(n120599) );
  BUF_X1 U83416 ( .A(n113904), .Z(n120600) );
  BUF_X1 U83417 ( .A(n113904), .Z(n120601) );
  BUF_X1 U83418 ( .A(n113904), .Z(n120602) );
  BUF_X1 U83419 ( .A(n113904), .Z(n120603) );
  BUF_X1 U83420 ( .A(n113991), .Z(n120537) );
  BUF_X1 U83421 ( .A(n113991), .Z(n120538) );
  BUF_X1 U83422 ( .A(n113991), .Z(n120539) );
  BUF_X1 U83423 ( .A(n113991), .Z(n120540) );
  BUF_X1 U83424 ( .A(n113991), .Z(n120541) );
  BUF_X1 U83425 ( .A(n114214), .Z(n120379) );
  BUF_X1 U83426 ( .A(n114579), .Z(n120253) );
  BUF_X1 U83427 ( .A(n114579), .Z(n120254) );
  BUF_X1 U83428 ( .A(n114579), .Z(n120255) );
  BUF_X1 U83429 ( .A(n114133), .Z(n120464) );
  BUF_X1 U83430 ( .A(n114133), .Z(n120465) );
  BUF_X1 U83431 ( .A(n114133), .Z(n120466) );
  BUF_X1 U83432 ( .A(n114133), .Z(n120467) );
  BUF_X1 U83433 ( .A(n114133), .Z(n120468) );
  BUF_X1 U83434 ( .A(n114137), .Z(n120440) );
  BUF_X1 U83435 ( .A(n114137), .Z(n120441) );
  BUF_X1 U83436 ( .A(n114137), .Z(n120442) );
  BUF_X1 U83437 ( .A(n114137), .Z(n120443) );
  BUF_X1 U83438 ( .A(n114137), .Z(n120444) );
  BUF_X1 U83439 ( .A(n114057), .Z(n120512) );
  BUF_X1 U83440 ( .A(n114057), .Z(n120513) );
  BUF_X1 U83441 ( .A(n114057), .Z(n120514) );
  BUF_X1 U83442 ( .A(n114057), .Z(n120515) );
  BUF_X1 U83443 ( .A(n114057), .Z(n120516) );
  BUF_X1 U83444 ( .A(n114129), .Z(n120488) );
  BUF_X1 U83445 ( .A(n114129), .Z(n120489) );
  BUF_X1 U83446 ( .A(n114129), .Z(n120490) );
  BUF_X1 U83447 ( .A(n114129), .Z(n120491) );
  BUF_X1 U83448 ( .A(n114129), .Z(n120492) );
  BUF_X1 U83449 ( .A(n114131), .Z(n120476) );
  BUF_X1 U83450 ( .A(n114131), .Z(n120477) );
  BUF_X1 U83451 ( .A(n114131), .Z(n120478) );
  BUF_X1 U83452 ( .A(n114131), .Z(n120479) );
  BUF_X1 U83453 ( .A(n114131), .Z(n120480) );
  BUF_X1 U83454 ( .A(n114135), .Z(n120452) );
  BUF_X1 U83455 ( .A(n114135), .Z(n120453) );
  BUF_X1 U83456 ( .A(n114135), .Z(n120454) );
  BUF_X1 U83457 ( .A(n114135), .Z(n120455) );
  BUF_X1 U83458 ( .A(n114135), .Z(n120456) );
  BUF_X1 U83459 ( .A(n113912), .Z(n120575) );
  BUF_X1 U83460 ( .A(n113912), .Z(n120576) );
  BUF_X1 U83461 ( .A(n113912), .Z(n120577) );
  BUF_X1 U83462 ( .A(n113912), .Z(n120578) );
  BUF_X1 U83463 ( .A(n113912), .Z(n120579) );
  BUF_X1 U83464 ( .A(n114124), .Z(n120500) );
  BUF_X1 U83465 ( .A(n114124), .Z(n120501) );
  BUF_X1 U83466 ( .A(n114124), .Z(n120502) );
  BUF_X1 U83467 ( .A(n114124), .Z(n120503) );
  BUF_X1 U83468 ( .A(n114124), .Z(n120504) );
  BUF_X1 U83469 ( .A(n113982), .Z(n120550) );
  BUF_X1 U83470 ( .A(n113982), .Z(n120551) );
  BUF_X1 U83471 ( .A(n113982), .Z(n120552) );
  BUF_X1 U83472 ( .A(n113982), .Z(n120553) );
  BUF_X1 U83473 ( .A(n113982), .Z(n120554) );
  BUF_X1 U83474 ( .A(n113910), .Z(n120587) );
  BUF_X1 U83475 ( .A(n113910), .Z(n120588) );
  BUF_X1 U83476 ( .A(n113910), .Z(n120589) );
  BUF_X1 U83477 ( .A(n113910), .Z(n120590) );
  BUF_X1 U83478 ( .A(n113910), .Z(n120591) );
  BUF_X1 U83479 ( .A(n113916), .Z(n120562) );
  BUF_X1 U83480 ( .A(n113916), .Z(n120563) );
  BUF_X1 U83481 ( .A(n113916), .Z(n120564) );
  BUF_X1 U83482 ( .A(n113916), .Z(n120565) );
  BUF_X1 U83483 ( .A(n113916), .Z(n120566) );
  BUF_X1 U83484 ( .A(n114301), .Z(n120354) );
  BUF_X1 U83485 ( .A(n114301), .Z(n120355) );
  BUF_X1 U83486 ( .A(n114301), .Z(n120356) );
  BUF_X1 U83487 ( .A(n114301), .Z(n120357) );
  BUF_X1 U83488 ( .A(n114301), .Z(n120358) );
  BUF_X1 U83489 ( .A(n114236), .Z(n120366) );
  BUF_X1 U83490 ( .A(n114236), .Z(n120367) );
  BUF_X1 U83491 ( .A(n114236), .Z(n120368) );
  BUF_X1 U83492 ( .A(n114236), .Z(n120369) );
  BUF_X1 U83493 ( .A(n114236), .Z(n120370) );
  BUF_X1 U83494 ( .A(n114307), .Z(n120329) );
  BUF_X1 U83495 ( .A(n114307), .Z(n120330) );
  BUF_X1 U83496 ( .A(n114307), .Z(n120331) );
  BUF_X1 U83497 ( .A(n114307), .Z(n120332) );
  BUF_X1 U83498 ( .A(n114307), .Z(n120333) );
  BUF_X1 U83499 ( .A(n114212), .Z(n120391) );
  BUF_X1 U83500 ( .A(n114212), .Z(n120392) );
  BUF_X1 U83501 ( .A(n114212), .Z(n120393) );
  BUF_X1 U83502 ( .A(n114212), .Z(n120394) );
  BUF_X1 U83503 ( .A(n114212), .Z(n120395) );
  BUF_X1 U83504 ( .A(n114373), .Z(n120317) );
  BUF_X1 U83505 ( .A(n114373), .Z(n120318) );
  BUF_X1 U83506 ( .A(n114373), .Z(n120319) );
  BUF_X1 U83507 ( .A(n114373), .Z(n120320) );
  BUF_X1 U83508 ( .A(n114373), .Z(n120321) );
  BUF_X1 U83509 ( .A(n114511), .Z(n120278) );
  BUF_X1 U83510 ( .A(n114511), .Z(n120279) );
  BUF_X1 U83511 ( .A(n114511), .Z(n120280) );
  BUF_X1 U83512 ( .A(n114511), .Z(n120281) );
  BUF_X1 U83513 ( .A(n114511), .Z(n120282) );
  BUF_X1 U83514 ( .A(n114576), .Z(n120266) );
  BUF_X1 U83515 ( .A(n114576), .Z(n120267) );
  BUF_X1 U83516 ( .A(n114576), .Z(n120268) );
  BUF_X1 U83517 ( .A(n114576), .Z(n120269) );
  BUF_X1 U83518 ( .A(n114576), .Z(n120270) );
  BUF_X1 U83519 ( .A(n114579), .Z(n120256) );
  BUF_X1 U83520 ( .A(n114579), .Z(n120257) );
  BUF_X1 U83521 ( .A(n114147), .Z(n120403) );
  BUF_X1 U83522 ( .A(n114147), .Z(n120404) );
  BUF_X1 U83523 ( .A(n114147), .Z(n120405) );
  BUF_X1 U83524 ( .A(n114147), .Z(n120406) );
  BUF_X1 U83525 ( .A(n114147), .Z(n120407) );
  BUF_X1 U83526 ( .A(n114379), .Z(n120304) );
  BUF_X1 U83527 ( .A(n114379), .Z(n120305) );
  BUF_X1 U83528 ( .A(n114379), .Z(n120306) );
  BUF_X1 U83529 ( .A(n114379), .Z(n120307) );
  BUF_X1 U83530 ( .A(n114214), .Z(n120380) );
  BUF_X1 U83531 ( .A(n114214), .Z(n120381) );
  BUF_X1 U83532 ( .A(n114214), .Z(n120382) );
  BUF_X1 U83533 ( .A(n114214), .Z(n120383) );
  BUF_X1 U83534 ( .A(n114140), .Z(n120428) );
  BUF_X1 U83535 ( .A(n114140), .Z(n120429) );
  BUF_X1 U83536 ( .A(n114140), .Z(n120430) );
  BUF_X1 U83537 ( .A(n114140), .Z(n120431) );
  BUF_X1 U83538 ( .A(n114140), .Z(n120432) );
  BUF_X1 U83539 ( .A(n114143), .Z(n120416) );
  BUF_X1 U83540 ( .A(n114143), .Z(n120417) );
  BUF_X1 U83541 ( .A(n114143), .Z(n120418) );
  BUF_X1 U83542 ( .A(n114143), .Z(n120419) );
  BUF_X1 U83543 ( .A(n114143), .Z(n120420) );
  BUF_X1 U83544 ( .A(n114304), .Z(n120342) );
  BUF_X1 U83545 ( .A(n114304), .Z(n120343) );
  BUF_X1 U83546 ( .A(n114304), .Z(n120344) );
  BUF_X1 U83547 ( .A(n114304), .Z(n120345) );
  BUF_X1 U83548 ( .A(n114304), .Z(n120346) );
  BUF_X1 U83549 ( .A(n114445), .Z(n120291) );
  BUF_X1 U83550 ( .A(n114445), .Z(n120292) );
  BUF_X1 U83551 ( .A(n114445), .Z(n120293) );
  BUF_X1 U83552 ( .A(n114445), .Z(n120294) );
  BUF_X1 U83553 ( .A(n114445), .Z(n120295) );
  BUF_X1 U83554 ( .A(n114053), .Z(n120525) );
  BUF_X1 U83555 ( .A(n114053), .Z(n120526) );
  BUF_X1 U83556 ( .A(n114053), .Z(n120527) );
  BUF_X1 U83557 ( .A(n114053), .Z(n120528) );
  BUF_X1 U83558 ( .A(n114053), .Z(n120529) );
  BUF_X1 U83559 ( .A(n114379), .Z(n120308) );
  BUF_X1 U83560 ( .A(n114689), .Z(n120100) );
  BUF_X1 U83561 ( .A(n114689), .Z(n120096) );
  BUF_X1 U83562 ( .A(n114689), .Z(n120097) );
  BUF_X1 U83563 ( .A(n114689), .Z(n120098) );
  BUF_X1 U83564 ( .A(n114689), .Z(n120099) );
  BUF_X1 U83565 ( .A(n113767), .Z(n120821) );
  BUF_X1 U83566 ( .A(n113766), .Z(n120827) );
  BUF_X1 U83567 ( .A(n113766), .Z(n120828) );
  OAI21_X1 U83568 ( .B1(n113894), .B2(n114141), .A(n120624), .ZN(n114139) );
  NAND2_X1 U83569 ( .A1(n116447), .A2(n116463), .ZN(n114689) );
  BUF_X1 U83570 ( .A(n116522), .Z(n119887) );
  BUF_X1 U83571 ( .A(n116522), .Z(n119888) );
  BUF_X1 U83572 ( .A(n116522), .Z(n119889) );
  BUF_X1 U83573 ( .A(n116522), .Z(n119890) );
  BUF_X1 U83574 ( .A(n114691), .Z(n120088) );
  BUF_X1 U83575 ( .A(n114698), .Z(n120064) );
  BUF_X1 U83576 ( .A(n116522), .Z(n119886) );
  BUF_X1 U83577 ( .A(n114691), .Z(n120084) );
  BUF_X1 U83578 ( .A(n114698), .Z(n120060) );
  BUF_X1 U83579 ( .A(n114691), .Z(n120085) );
  BUF_X1 U83580 ( .A(n114698), .Z(n120061) );
  BUF_X1 U83581 ( .A(n114691), .Z(n120086) );
  BUF_X1 U83582 ( .A(n114698), .Z(n120062) );
  BUF_X1 U83583 ( .A(n114691), .Z(n120087) );
  BUF_X1 U83584 ( .A(n114698), .Z(n120063) );
  BUF_X1 U83585 ( .A(n116490), .Z(n120025) );
  BUF_X1 U83586 ( .A(n116490), .Z(n120026) );
  BUF_X1 U83587 ( .A(n116490), .Z(n120027) );
  BUF_X1 U83588 ( .A(n116490), .Z(n120028) );
  BUF_X1 U83589 ( .A(n114662), .Z(n120202) );
  BUF_X1 U83590 ( .A(n116490), .Z(n120024) );
  BUF_X1 U83591 ( .A(n114662), .Z(n120198) );
  BUF_X1 U83592 ( .A(n114662), .Z(n120199) );
  BUF_X1 U83593 ( .A(n114662), .Z(n120200) );
  BUF_X1 U83594 ( .A(n114662), .Z(n120201) );
  BUF_X1 U83595 ( .A(n114657), .Z(n120226) );
  BUF_X1 U83596 ( .A(n114657), .Z(n120222) );
  BUF_X1 U83597 ( .A(n114657), .Z(n120223) );
  BUF_X1 U83598 ( .A(n114657), .Z(n120224) );
  BUF_X1 U83599 ( .A(n114657), .Z(n120225) );
  BUF_X1 U83600 ( .A(n116495), .Z(n120001) );
  BUF_X1 U83601 ( .A(n116502), .Z(n119977) );
  BUF_X1 U83602 ( .A(n116507), .Z(n119953) );
  BUF_X1 U83603 ( .A(n116495), .Z(n120002) );
  BUF_X1 U83604 ( .A(n116502), .Z(n119978) );
  BUF_X1 U83605 ( .A(n116507), .Z(n119954) );
  BUF_X1 U83606 ( .A(n116495), .Z(n120003) );
  BUF_X1 U83607 ( .A(n116502), .Z(n119979) );
  BUF_X1 U83608 ( .A(n116507), .Z(n119955) );
  BUF_X1 U83609 ( .A(n116495), .Z(n120004) );
  BUF_X1 U83610 ( .A(n116502), .Z(n119980) );
  BUF_X1 U83611 ( .A(n116507), .Z(n119956) );
  BUF_X1 U83612 ( .A(n114669), .Z(n120178) );
  BUF_X1 U83613 ( .A(n114675), .Z(n120154) );
  BUF_X1 U83614 ( .A(n116495), .Z(n120000) );
  BUF_X1 U83615 ( .A(n116502), .Z(n119976) );
  BUF_X1 U83616 ( .A(n116507), .Z(n119952) );
  BUF_X1 U83617 ( .A(n114669), .Z(n120174) );
  BUF_X1 U83618 ( .A(n114675), .Z(n120150) );
  BUF_X1 U83619 ( .A(n114669), .Z(n120175) );
  BUF_X1 U83620 ( .A(n114675), .Z(n120151) );
  BUF_X1 U83621 ( .A(n114669), .Z(n120176) );
  BUF_X1 U83622 ( .A(n114675), .Z(n120152) );
  BUF_X1 U83623 ( .A(n114669), .Z(n120177) );
  BUF_X1 U83624 ( .A(n114675), .Z(n120153) );
  BUF_X1 U83625 ( .A(n116523), .Z(n119881) );
  BUF_X1 U83626 ( .A(n116523), .Z(n119882) );
  BUF_X1 U83627 ( .A(n116523), .Z(n119883) );
  BUF_X1 U83628 ( .A(n116523), .Z(n119884) );
  BUF_X1 U83629 ( .A(n116523), .Z(n119880) );
  BUF_X1 U83630 ( .A(n116529), .Z(n119857) );
  BUF_X1 U83631 ( .A(n116529), .Z(n119858) );
  BUF_X1 U83632 ( .A(n116529), .Z(n119859) );
  BUF_X1 U83633 ( .A(n116529), .Z(n119860) );
  BUF_X1 U83634 ( .A(n114693), .Z(n120082) );
  BUF_X1 U83635 ( .A(n114700), .Z(n120058) );
  BUF_X1 U83636 ( .A(n116529), .Z(n119856) );
  BUF_X1 U83637 ( .A(n114693), .Z(n120078) );
  BUF_X1 U83638 ( .A(n114700), .Z(n120054) );
  BUF_X1 U83639 ( .A(n114693), .Z(n120079) );
  BUF_X1 U83640 ( .A(n114700), .Z(n120055) );
  BUF_X1 U83641 ( .A(n114693), .Z(n120080) );
  BUF_X1 U83642 ( .A(n114700), .Z(n120056) );
  BUF_X1 U83643 ( .A(n114693), .Z(n120081) );
  BUF_X1 U83644 ( .A(n114700), .Z(n120057) );
  BUF_X1 U83645 ( .A(n116492), .Z(n120013) );
  BUF_X1 U83646 ( .A(n116499), .Z(n119989) );
  BUF_X1 U83647 ( .A(n116487), .Z(n120037) );
  BUF_X1 U83648 ( .A(n116504), .Z(n119965) );
  BUF_X1 U83649 ( .A(n116492), .Z(n120014) );
  BUF_X1 U83650 ( .A(n116499), .Z(n119990) );
  BUF_X1 U83651 ( .A(n116487), .Z(n120038) );
  BUF_X1 U83652 ( .A(n116504), .Z(n119966) );
  BUF_X1 U83653 ( .A(n116492), .Z(n120015) );
  BUF_X1 U83654 ( .A(n116499), .Z(n119991) );
  BUF_X1 U83655 ( .A(n116487), .Z(n120039) );
  BUF_X1 U83656 ( .A(n116504), .Z(n119967) );
  BUF_X1 U83657 ( .A(n116492), .Z(n120016) );
  BUF_X1 U83658 ( .A(n116499), .Z(n119992) );
  BUF_X1 U83659 ( .A(n116487), .Z(n120040) );
  BUF_X1 U83660 ( .A(n116504), .Z(n119968) );
  BUF_X1 U83661 ( .A(n114672), .Z(n120166) );
  BUF_X1 U83662 ( .A(n114672), .Z(n120163) );
  BUF_X1 U83663 ( .A(n114672), .Z(n120164) );
  BUF_X1 U83664 ( .A(n114672), .Z(n120165) );
  BUF_X1 U83665 ( .A(n114654), .Z(n120238) );
  BUF_X1 U83666 ( .A(n114654), .Z(n120235) );
  BUF_X1 U83667 ( .A(n114654), .Z(n120236) );
  BUF_X1 U83668 ( .A(n114654), .Z(n120237) );
  BUF_X1 U83669 ( .A(n114659), .Z(n120214) );
  BUF_X1 U83670 ( .A(n114666), .Z(n120190) );
  BUF_X1 U83671 ( .A(n114659), .Z(n120211) );
  BUF_X1 U83672 ( .A(n114666), .Z(n120187) );
  BUF_X1 U83673 ( .A(n114659), .Z(n120212) );
  BUF_X1 U83674 ( .A(n114666), .Z(n120188) );
  BUF_X1 U83675 ( .A(n114659), .Z(n120213) );
  BUF_X1 U83676 ( .A(n114666), .Z(n120189) );
  BUF_X1 U83677 ( .A(n114690), .Z(n120094) );
  BUF_X1 U83678 ( .A(n114690), .Z(n120090) );
  BUF_X1 U83679 ( .A(n114690), .Z(n120091) );
  BUF_X1 U83680 ( .A(n114690), .Z(n120092) );
  BUF_X1 U83681 ( .A(n114690), .Z(n120093) );
  BUF_X1 U83682 ( .A(n116521), .Z(n119893) );
  BUF_X1 U83683 ( .A(n116521), .Z(n119894) );
  BUF_X1 U83684 ( .A(n116521), .Z(n119895) );
  BUF_X1 U83685 ( .A(n116521), .Z(n119896) );
  BUF_X1 U83686 ( .A(n116521), .Z(n119892) );
  BUF_X1 U83687 ( .A(n114688), .Z(n120106) );
  BUF_X1 U83688 ( .A(n114688), .Z(n120102) );
  BUF_X1 U83689 ( .A(n114688), .Z(n120103) );
  BUF_X1 U83690 ( .A(n114688), .Z(n120104) );
  BUF_X1 U83691 ( .A(n114688), .Z(n120105) );
  BUF_X1 U83692 ( .A(n116519), .Z(n119905) );
  BUF_X1 U83693 ( .A(n116519), .Z(n119906) );
  BUF_X1 U83694 ( .A(n116519), .Z(n119907) );
  BUF_X1 U83695 ( .A(n116519), .Z(n119908) );
  BUF_X1 U83696 ( .A(n116519), .Z(n119904) );
  BUF_X1 U83697 ( .A(n116520), .Z(n119899) );
  BUF_X1 U83698 ( .A(n116520), .Z(n119900) );
  BUF_X1 U83699 ( .A(n116520), .Z(n119901) );
  BUF_X1 U83700 ( .A(n116520), .Z(n119902) );
  BUF_X1 U83701 ( .A(n116520), .Z(n119898) );
  BUF_X1 U83702 ( .A(n114670), .Z(n120172) );
  BUF_X1 U83703 ( .A(n114676), .Z(n120148) );
  BUF_X1 U83704 ( .A(n114670), .Z(n120168) );
  BUF_X1 U83705 ( .A(n114676), .Z(n120144) );
  BUF_X1 U83706 ( .A(n114670), .Z(n120169) );
  BUF_X1 U83707 ( .A(n114676), .Z(n120145) );
  BUF_X1 U83708 ( .A(n114670), .Z(n120170) );
  BUF_X1 U83709 ( .A(n114676), .Z(n120146) );
  BUF_X1 U83710 ( .A(n114670), .Z(n120171) );
  BUF_X1 U83711 ( .A(n114676), .Z(n120147) );
  BUF_X1 U83712 ( .A(n116497), .Z(n119995) );
  BUF_X1 U83713 ( .A(n116503), .Z(n119971) );
  BUF_X1 U83714 ( .A(n116508), .Z(n119947) );
  BUF_X1 U83715 ( .A(n116497), .Z(n119996) );
  BUF_X1 U83716 ( .A(n116503), .Z(n119972) );
  BUF_X1 U83717 ( .A(n116508), .Z(n119948) );
  BUF_X1 U83718 ( .A(n116497), .Z(n119997) );
  BUF_X1 U83719 ( .A(n116503), .Z(n119973) );
  BUF_X1 U83720 ( .A(n116508), .Z(n119949) );
  BUF_X1 U83721 ( .A(n116497), .Z(n119998) );
  BUF_X1 U83722 ( .A(n116503), .Z(n119974) );
  BUF_X1 U83723 ( .A(n116508), .Z(n119950) );
  BUF_X1 U83724 ( .A(n114664), .Z(n120196) );
  BUF_X1 U83725 ( .A(n116497), .Z(n119994) );
  BUF_X1 U83726 ( .A(n116503), .Z(n119970) );
  BUF_X1 U83727 ( .A(n116508), .Z(n119946) );
  BUF_X1 U83728 ( .A(n114664), .Z(n120192) );
  BUF_X1 U83729 ( .A(n114664), .Z(n120193) );
  BUF_X1 U83730 ( .A(n114664), .Z(n120194) );
  BUF_X1 U83731 ( .A(n114664), .Z(n120195) );
  NAND2_X1 U83732 ( .A1(n120628), .A2(n120248), .ZN(n114645) );
  NAND2_X1 U83733 ( .A1(n120628), .A2(n120617), .ZN(n113897) );
  NAND2_X1 U83734 ( .A1(n120628), .A2(n120605), .ZN(n113904) );
  BUF_X1 U83735 ( .A(n114213), .Z(n120389) );
  BUF_X1 U83736 ( .A(n114132), .Z(n120470) );
  BUF_X1 U83737 ( .A(n114136), .Z(n120446) );
  BUF_X1 U83738 ( .A(n114128), .Z(n120494) );
  BUF_X1 U83739 ( .A(n114130), .Z(n120482) );
  BUF_X1 U83740 ( .A(n114134), .Z(n120458) );
  BUF_X1 U83741 ( .A(n113911), .Z(n120581) );
  BUF_X1 U83742 ( .A(n114122), .Z(n120506) );
  BUF_X1 U83743 ( .A(n113980), .Z(n120556) );
  BUF_X1 U83744 ( .A(n113909), .Z(n120593) );
  BUF_X1 U83745 ( .A(n114300), .Z(n120360) );
  BUF_X1 U83746 ( .A(n114211), .Z(n120397) );
  BUF_X1 U83747 ( .A(n114372), .Z(n120323) );
  BUF_X1 U83748 ( .A(n114575), .Z(n120272) );
  BUF_X1 U83749 ( .A(n114142), .Z(n120422) );
  BUF_X1 U83750 ( .A(n114303), .Z(n120348) );
  BUF_X1 U83751 ( .A(n114213), .Z(n120385) );
  BUF_X1 U83752 ( .A(n114052), .Z(n120531) );
  BUF_X1 U83753 ( .A(n113895), .Z(n120617) );
  BUF_X1 U83754 ( .A(n113902), .Z(n120605) );
  BUF_X1 U83755 ( .A(n114132), .Z(n120471) );
  BUF_X1 U83756 ( .A(n114132), .Z(n120472) );
  BUF_X1 U83757 ( .A(n114132), .Z(n120473) );
  BUF_X1 U83758 ( .A(n114132), .Z(n120474) );
  BUF_X1 U83759 ( .A(n114136), .Z(n120447) );
  BUF_X1 U83760 ( .A(n114136), .Z(n120448) );
  BUF_X1 U83761 ( .A(n114136), .Z(n120449) );
  BUF_X1 U83762 ( .A(n114136), .Z(n120450) );
  BUF_X1 U83763 ( .A(n114128), .Z(n120495) );
  BUF_X1 U83764 ( .A(n114128), .Z(n120496) );
  BUF_X1 U83765 ( .A(n114128), .Z(n120497) );
  BUF_X1 U83766 ( .A(n114128), .Z(n120498) );
  BUF_X1 U83767 ( .A(n114130), .Z(n120483) );
  BUF_X1 U83768 ( .A(n114130), .Z(n120484) );
  BUF_X1 U83769 ( .A(n114130), .Z(n120485) );
  BUF_X1 U83770 ( .A(n114130), .Z(n120486) );
  BUF_X1 U83771 ( .A(n114134), .Z(n120459) );
  BUF_X1 U83772 ( .A(n114134), .Z(n120460) );
  BUF_X1 U83773 ( .A(n114134), .Z(n120461) );
  BUF_X1 U83774 ( .A(n114134), .Z(n120462) );
  BUF_X1 U83775 ( .A(n113911), .Z(n120582) );
  BUF_X1 U83776 ( .A(n113911), .Z(n120583) );
  BUF_X1 U83777 ( .A(n113911), .Z(n120584) );
  BUF_X1 U83778 ( .A(n113911), .Z(n120585) );
  BUF_X1 U83779 ( .A(n114122), .Z(n120507) );
  BUF_X1 U83780 ( .A(n114122), .Z(n120508) );
  BUF_X1 U83781 ( .A(n114122), .Z(n120509) );
  BUF_X1 U83782 ( .A(n114122), .Z(n120510) );
  BUF_X1 U83783 ( .A(n113980), .Z(n120557) );
  BUF_X1 U83784 ( .A(n113980), .Z(n120558) );
  BUF_X1 U83785 ( .A(n113980), .Z(n120559) );
  BUF_X1 U83786 ( .A(n113980), .Z(n120560) );
  BUF_X1 U83787 ( .A(n113909), .Z(n120594) );
  BUF_X1 U83788 ( .A(n113909), .Z(n120595) );
  BUF_X1 U83789 ( .A(n113909), .Z(n120596) );
  BUF_X1 U83790 ( .A(n113909), .Z(n120597) );
  BUF_X1 U83791 ( .A(n114300), .Z(n120361) );
  BUF_X1 U83792 ( .A(n114300), .Z(n120362) );
  BUF_X1 U83793 ( .A(n114300), .Z(n120363) );
  BUF_X1 U83794 ( .A(n114300), .Z(n120364) );
  BUF_X1 U83795 ( .A(n114211), .Z(n120398) );
  BUF_X1 U83796 ( .A(n114211), .Z(n120399) );
  BUF_X1 U83797 ( .A(n114211), .Z(n120400) );
  BUF_X1 U83798 ( .A(n114211), .Z(n120401) );
  BUF_X1 U83799 ( .A(n114372), .Z(n120324) );
  BUF_X1 U83800 ( .A(n114372), .Z(n120325) );
  BUF_X1 U83801 ( .A(n114372), .Z(n120326) );
  BUF_X1 U83802 ( .A(n114372), .Z(n120327) );
  BUF_X1 U83803 ( .A(n114575), .Z(n120273) );
  BUF_X1 U83804 ( .A(n114575), .Z(n120274) );
  BUF_X1 U83805 ( .A(n114575), .Z(n120275) );
  BUF_X1 U83806 ( .A(n114575), .Z(n120276) );
  BUF_X1 U83807 ( .A(n114213), .Z(n120386) );
  BUF_X1 U83808 ( .A(n114142), .Z(n120423) );
  BUF_X1 U83809 ( .A(n114142), .Z(n120424) );
  BUF_X1 U83810 ( .A(n114142), .Z(n120425) );
  BUF_X1 U83811 ( .A(n114142), .Z(n120426) );
  BUF_X1 U83812 ( .A(n114303), .Z(n120349) );
  BUF_X1 U83813 ( .A(n114303), .Z(n120350) );
  BUF_X1 U83814 ( .A(n114303), .Z(n120351) );
  BUF_X1 U83815 ( .A(n114303), .Z(n120352) );
  BUF_X1 U83816 ( .A(n114213), .Z(n120387) );
  BUF_X1 U83817 ( .A(n114052), .Z(n120532) );
  BUF_X1 U83818 ( .A(n114052), .Z(n120533) );
  BUF_X1 U83819 ( .A(n114052), .Z(n120534) );
  BUF_X1 U83820 ( .A(n114052), .Z(n120535) );
  BUF_X1 U83821 ( .A(n113895), .Z(n120618) );
  BUF_X1 U83822 ( .A(n113895), .Z(n120619) );
  BUF_X1 U83823 ( .A(n113895), .Z(n120620) );
  BUF_X1 U83824 ( .A(n113895), .Z(n120621) );
  BUF_X1 U83825 ( .A(n113902), .Z(n120606) );
  BUF_X1 U83826 ( .A(n113902), .Z(n120607) );
  BUF_X1 U83827 ( .A(n113902), .Z(n120608) );
  BUF_X1 U83828 ( .A(n113902), .Z(n120609) );
  BUF_X1 U83829 ( .A(n116513), .Z(n119941) );
  BUF_X1 U83830 ( .A(n116515), .Z(n119929) );
  BUF_X1 U83831 ( .A(n116517), .Z(n119917) );
  BUF_X1 U83832 ( .A(n116513), .Z(n119942) );
  BUF_X1 U83833 ( .A(n116515), .Z(n119930) );
  BUF_X1 U83834 ( .A(n116517), .Z(n119918) );
  BUF_X1 U83835 ( .A(n116513), .Z(n119943) );
  BUF_X1 U83836 ( .A(n116515), .Z(n119931) );
  BUF_X1 U83837 ( .A(n116517), .Z(n119919) );
  BUF_X1 U83838 ( .A(n116513), .Z(n119944) );
  BUF_X1 U83839 ( .A(n116515), .Z(n119932) );
  BUF_X1 U83840 ( .A(n116517), .Z(n119920) );
  BUF_X1 U83841 ( .A(n114686), .Z(n120118) );
  BUF_X1 U83842 ( .A(n114686), .Z(n120114) );
  BUF_X1 U83843 ( .A(n114696), .Z(n120072) );
  BUF_X1 U83844 ( .A(n114686), .Z(n120115) );
  BUF_X1 U83845 ( .A(n114684), .Z(n120130) );
  BUF_X1 U83846 ( .A(n114682), .Z(n120142) );
  BUF_X1 U83847 ( .A(n114696), .Z(n120076) );
  BUF_X1 U83848 ( .A(n116513), .Z(n119940) );
  BUF_X1 U83849 ( .A(n116515), .Z(n119928) );
  BUF_X1 U83850 ( .A(n116517), .Z(n119916) );
  BUF_X1 U83851 ( .A(n114684), .Z(n120126) );
  BUF_X1 U83852 ( .A(n114682), .Z(n120138) );
  BUF_X1 U83853 ( .A(n114684), .Z(n120127) );
  BUF_X1 U83854 ( .A(n114682), .Z(n120139) );
  BUF_X1 U83855 ( .A(n114696), .Z(n120073) );
  BUF_X1 U83856 ( .A(n114686), .Z(n120116) );
  BUF_X1 U83857 ( .A(n114686), .Z(n120117) );
  BUF_X1 U83858 ( .A(n114684), .Z(n120128) );
  BUF_X1 U83859 ( .A(n114682), .Z(n120140) );
  BUF_X1 U83860 ( .A(n114696), .Z(n120074) );
  BUF_X1 U83861 ( .A(n114684), .Z(n120129) );
  BUF_X1 U83862 ( .A(n114682), .Z(n120141) );
  BUF_X1 U83863 ( .A(n114696), .Z(n120075) );
  BUF_X1 U83864 ( .A(n116531), .Z(n119851) );
  BUF_X1 U83865 ( .A(n116526), .Z(n119875) );
  BUF_X1 U83866 ( .A(n116531), .Z(n119852) );
  BUF_X1 U83867 ( .A(n116526), .Z(n119876) );
  BUF_X1 U83868 ( .A(n116531), .Z(n119853) );
  BUF_X1 U83869 ( .A(n116526), .Z(n119877) );
  BUF_X1 U83870 ( .A(n116531), .Z(n119854) );
  BUF_X1 U83871 ( .A(n116526), .Z(n119878) );
  BUF_X1 U83872 ( .A(n114702), .Z(n120052) );
  BUF_X1 U83873 ( .A(n116531), .Z(n119850) );
  BUF_X1 U83874 ( .A(n116526), .Z(n119874) );
  BUF_X1 U83875 ( .A(n114702), .Z(n120048) );
  BUF_X1 U83876 ( .A(n114702), .Z(n120049) );
  BUF_X1 U83877 ( .A(n114702), .Z(n120050) );
  BUF_X1 U83878 ( .A(n114702), .Z(n120051) );
  BUF_X1 U83879 ( .A(n114213), .Z(n120388) );
  NAND2_X1 U83880 ( .A1(n120625), .A2(n120360), .ZN(n114301) );
  NAND2_X1 U83881 ( .A1(n120625), .A2(n120374), .ZN(n114236) );
  NAND2_X1 U83882 ( .A1(n120625), .A2(n120411), .ZN(n114147) );
  NAND2_X1 U83883 ( .A1(n120625), .A2(n120385), .ZN(n114214) );
  NAND2_X1 U83884 ( .A1(n120626), .A2(n120506), .ZN(n114124) );
  NAND2_X1 U83885 ( .A1(n120627), .A2(n120556), .ZN(n113982) );
  NAND2_X1 U83886 ( .A1(n120626), .A2(n120470), .ZN(n114133) );
  NAND2_X1 U83887 ( .A1(n120626), .A2(n120446), .ZN(n114137) );
  NAND2_X1 U83888 ( .A1(n120627), .A2(n120520), .ZN(n114057) );
  NAND2_X1 U83889 ( .A1(n120626), .A2(n120494), .ZN(n114129) );
  NAND2_X1 U83890 ( .A1(n120626), .A2(n120482), .ZN(n114131) );
  NAND2_X1 U83891 ( .A1(n120626), .A2(n120458), .ZN(n114135) );
  NAND2_X1 U83892 ( .A1(n120627), .A2(n120581), .ZN(n113912) );
  NAND2_X1 U83893 ( .A1(n120627), .A2(n120593), .ZN(n113910) );
  NAND2_X1 U83894 ( .A1(n120627), .A2(n120570), .ZN(n113916) );
  NAND2_X1 U83895 ( .A1(n120626), .A2(n120337), .ZN(n114307) );
  NAND2_X1 U83896 ( .A1(n120626), .A2(n120397), .ZN(n114212) );
  NAND2_X1 U83897 ( .A1(n120627), .A2(n120323), .ZN(n114373) );
  NAND2_X1 U83898 ( .A1(n120627), .A2(n120286), .ZN(n114511) );
  NAND2_X1 U83899 ( .A1(n120627), .A2(n120272), .ZN(n114576) );
  NAND2_X1 U83900 ( .A1(n120627), .A2(n120261), .ZN(n114579) );
  NAND2_X1 U83901 ( .A1(n120627), .A2(n120545), .ZN(n113991) );
  NAND2_X1 U83902 ( .A1(n120626), .A2(n120434), .ZN(n114140) );
  NAND2_X1 U83903 ( .A1(n120626), .A2(n120422), .ZN(n114143) );
  NAND2_X1 U83904 ( .A1(n120626), .A2(n120348), .ZN(n114304) );
  NAND2_X1 U83905 ( .A1(n120627), .A2(n120299), .ZN(n114445) );
  NAND2_X1 U83906 ( .A1(n120627), .A2(n120531), .ZN(n114053) );
  NAND2_X1 U83907 ( .A1(n120626), .A2(n120312), .ZN(n114379) );
  BUF_X1 U83908 ( .A(n116514), .Z(n119935) );
  BUF_X1 U83909 ( .A(n116518), .Z(n119911) );
  BUF_X1 U83910 ( .A(n116514), .Z(n119936) );
  BUF_X1 U83911 ( .A(n116518), .Z(n119912) );
  BUF_X1 U83912 ( .A(n116514), .Z(n119937) );
  BUF_X1 U83913 ( .A(n116518), .Z(n119913) );
  BUF_X1 U83914 ( .A(n116514), .Z(n119938) );
  BUF_X1 U83915 ( .A(n116518), .Z(n119914) );
  BUF_X1 U83916 ( .A(n114685), .Z(n120124) );
  BUF_X1 U83917 ( .A(n114685), .Z(n120120) );
  BUF_X1 U83918 ( .A(n114685), .Z(n120121) );
  BUF_X1 U83919 ( .A(n114685), .Z(n120122) );
  BUF_X1 U83920 ( .A(n114685), .Z(n120123) );
  BUF_X1 U83921 ( .A(n114683), .Z(n120136) );
  BUF_X1 U83922 ( .A(n114703), .Z(n120046) );
  BUF_X1 U83923 ( .A(n116514), .Z(n119934) );
  BUF_X1 U83924 ( .A(n116518), .Z(n119910) );
  BUF_X1 U83925 ( .A(n114683), .Z(n120132) );
  BUF_X1 U83926 ( .A(n114703), .Z(n120042) );
  BUF_X1 U83927 ( .A(n114683), .Z(n120133) );
  BUF_X1 U83928 ( .A(n114703), .Z(n120043) );
  BUF_X1 U83929 ( .A(n114683), .Z(n120134) );
  BUF_X1 U83930 ( .A(n114703), .Z(n120044) );
  BUF_X1 U83931 ( .A(n114683), .Z(n120135) );
  BUF_X1 U83932 ( .A(n114703), .Z(n120045) );
  BUF_X1 U83933 ( .A(n116516), .Z(n119923) );
  BUF_X1 U83934 ( .A(n116532), .Z(n119845) );
  BUF_X1 U83935 ( .A(n116527), .Z(n119869) );
  BUF_X1 U83936 ( .A(n116516), .Z(n119924) );
  BUF_X1 U83937 ( .A(n116532), .Z(n119846) );
  BUF_X1 U83938 ( .A(n116527), .Z(n119870) );
  BUF_X1 U83939 ( .A(n116516), .Z(n119925) );
  BUF_X1 U83940 ( .A(n116532), .Z(n119847) );
  BUF_X1 U83941 ( .A(n116527), .Z(n119871) );
  BUF_X1 U83942 ( .A(n116516), .Z(n119926) );
  BUF_X1 U83943 ( .A(n116532), .Z(n119848) );
  BUF_X1 U83944 ( .A(n116527), .Z(n119872) );
  BUF_X1 U83945 ( .A(n114687), .Z(n120112) );
  BUF_X1 U83946 ( .A(n114697), .Z(n120070) );
  BUF_X1 U83947 ( .A(n116516), .Z(n119922) );
  BUF_X1 U83948 ( .A(n116532), .Z(n119844) );
  BUF_X1 U83949 ( .A(n116527), .Z(n119868) );
  BUF_X1 U83950 ( .A(n114687), .Z(n120108) );
  BUF_X1 U83951 ( .A(n114697), .Z(n120066) );
  BUF_X1 U83952 ( .A(n114687), .Z(n120109) );
  BUF_X1 U83953 ( .A(n114697), .Z(n120067) );
  BUF_X1 U83954 ( .A(n114687), .Z(n120110) );
  BUF_X1 U83955 ( .A(n114697), .Z(n120068) );
  BUF_X1 U83956 ( .A(n114687), .Z(n120111) );
  BUF_X1 U83957 ( .A(n114697), .Z(n120069) );
  BUF_X1 U83958 ( .A(n116493), .Z(n120007) );
  BUF_X1 U83959 ( .A(n116488), .Z(n120031) );
  BUF_X1 U83960 ( .A(n116505), .Z(n119959) );
  BUF_X1 U83961 ( .A(n116493), .Z(n120008) );
  BUF_X1 U83962 ( .A(n116488), .Z(n120032) );
  BUF_X1 U83963 ( .A(n116505), .Z(n119960) );
  BUF_X1 U83964 ( .A(n116493), .Z(n120009) );
  BUF_X1 U83965 ( .A(n116488), .Z(n120033) );
  BUF_X1 U83966 ( .A(n116505), .Z(n119961) );
  BUF_X1 U83967 ( .A(n116493), .Z(n120010) );
  BUF_X1 U83968 ( .A(n116488), .Z(n120034) );
  BUF_X1 U83969 ( .A(n116505), .Z(n119962) );
  BUF_X1 U83970 ( .A(n114655), .Z(n120232) );
  BUF_X1 U83971 ( .A(n114667), .Z(n120184) );
  BUF_X1 U83972 ( .A(n116493), .Z(n120006) );
  BUF_X1 U83973 ( .A(n116488), .Z(n120030) );
  BUF_X1 U83974 ( .A(n116505), .Z(n119958) );
  BUF_X1 U83975 ( .A(n114655), .Z(n120228) );
  BUF_X1 U83976 ( .A(n114667), .Z(n120180) );
  BUF_X1 U83977 ( .A(n114655), .Z(n120229) );
  BUF_X1 U83978 ( .A(n114667), .Z(n120181) );
  BUF_X1 U83979 ( .A(n114655), .Z(n120230) );
  BUF_X1 U83980 ( .A(n114667), .Z(n120182) );
  BUF_X1 U83981 ( .A(n114655), .Z(n120231) );
  BUF_X1 U83982 ( .A(n114667), .Z(n120183) );
  BUF_X1 U83983 ( .A(n116500), .Z(n119983) );
  BUF_X1 U83984 ( .A(n116500), .Z(n119984) );
  BUF_X1 U83985 ( .A(n116500), .Z(n119985) );
  BUF_X1 U83986 ( .A(n116500), .Z(n119986) );
  BUF_X1 U83987 ( .A(n114660), .Z(n120208) );
  BUF_X1 U83988 ( .A(n114673), .Z(n120160) );
  BUF_X1 U83989 ( .A(n116500), .Z(n119982) );
  BUF_X1 U83990 ( .A(n114660), .Z(n120204) );
  BUF_X1 U83991 ( .A(n114673), .Z(n120156) );
  BUF_X1 U83992 ( .A(n114660), .Z(n120205) );
  BUF_X1 U83993 ( .A(n114673), .Z(n120157) );
  BUF_X1 U83994 ( .A(n114660), .Z(n120206) );
  BUF_X1 U83995 ( .A(n114673), .Z(n120158) );
  BUF_X1 U83996 ( .A(n114660), .Z(n120207) );
  BUF_X1 U83997 ( .A(n114673), .Z(n120159) );
  BUF_X1 U83998 ( .A(n114672), .Z(n120162) );
  BUF_X1 U83999 ( .A(n116492), .Z(n120012) );
  BUF_X1 U84000 ( .A(n116499), .Z(n119988) );
  BUF_X1 U84001 ( .A(n116487), .Z(n120036) );
  BUF_X1 U84002 ( .A(n116504), .Z(n119964) );
  BUF_X1 U84003 ( .A(n114654), .Z(n120234) );
  BUF_X1 U84004 ( .A(n114659), .Z(n120210) );
  BUF_X1 U84005 ( .A(n114666), .Z(n120186) );
  NAND2_X1 U84006 ( .A1(n120628), .A2(n120829), .ZN(n113767) );
  OAI21_X1 U84007 ( .B1(n113893), .B2(n113894), .A(n120623), .ZN(n113766) );
  AND2_X1 U84008 ( .A1(n117949), .A2(n117948), .ZN(n116528) );
  BUF_X1 U84009 ( .A(n113914), .Z(n120568) );
  BUF_X1 U84010 ( .A(n113990), .Z(n120543) );
  BUF_X1 U84011 ( .A(n114643), .Z(n120246) );
  BUF_X1 U84012 ( .A(n114577), .Z(n120259) );
  BUF_X1 U84013 ( .A(n114055), .Z(n120518) );
  BUF_X1 U84014 ( .A(n114234), .Z(n120372) );
  BUF_X1 U84015 ( .A(n114305), .Z(n120335) );
  BUF_X1 U84016 ( .A(n114509), .Z(n120284) );
  BUF_X1 U84017 ( .A(n114145), .Z(n120409) );
  BUF_X1 U84018 ( .A(n114377), .Z(n120310) );
  BUF_X1 U84019 ( .A(n114443), .Z(n120297) );
  BUF_X1 U84020 ( .A(n113990), .Z(n120544) );
  BUF_X1 U84021 ( .A(n113914), .Z(n120569) );
  BUF_X1 U84022 ( .A(n114643), .Z(n120247) );
  BUF_X1 U84023 ( .A(n114055), .Z(n120519) );
  BUF_X1 U84024 ( .A(n114234), .Z(n120373) );
  BUF_X1 U84025 ( .A(n114305), .Z(n120336) );
  BUF_X1 U84026 ( .A(n114509), .Z(n120285) );
  BUF_X1 U84027 ( .A(n114577), .Z(n120260) );
  BUF_X1 U84028 ( .A(n114145), .Z(n120410) );
  BUF_X1 U84029 ( .A(n114443), .Z(n120298) );
  BUF_X1 U84030 ( .A(n114377), .Z(n120311) );
  NOR3_X1 U84031 ( .A1(n116478), .A2(n120216), .A3(n116475), .ZN(n116447) );
  NOR3_X1 U84032 ( .A1(n116470), .A2(n116469), .A3(n116471), .ZN(n116463) );
  NOR3_X1 U84033 ( .A1(n117967), .A2(n117970), .A3(n117958), .ZN(n117949) );
  OAI21_X1 U84034 ( .B1(n113901), .B2(n113908), .A(n120623), .ZN(n113909) );
  OAI21_X1 U84035 ( .B1(n113908), .B2(n114054), .A(n120623), .ZN(n114122) );
  OAI21_X1 U84036 ( .B1(n113913), .B2(n114121), .A(n120624), .ZN(n114132) );
  OAI21_X1 U84037 ( .B1(n113986), .B2(n114121), .A(n120624), .ZN(n114136) );
  OAI21_X1 U84038 ( .B1(n113908), .B2(n114121), .A(n120623), .ZN(n114128) );
  OAI21_X1 U84039 ( .B1(n113913), .B2(n114054), .A(n120624), .ZN(n114130) );
  OAI21_X1 U84040 ( .B1(n113986), .B2(n114054), .A(n120624), .ZN(n114134) );
  OAI21_X1 U84041 ( .B1(n113986), .B2(n114141), .A(n120625), .ZN(n114300) );
  OAI21_X1 U84042 ( .B1(n113908), .B2(n114144), .A(n120624), .ZN(n114211) );
  OAI21_X1 U84043 ( .B1(n113894), .B2(n114374), .A(n120625), .ZN(n114372) );
  OAI21_X1 U84044 ( .B1(n113913), .B2(n114374), .A(n120624), .ZN(n114575) );
  OAI21_X1 U84045 ( .B1(n113913), .B2(n114141), .A(n120624), .ZN(n114213) );
  OAI21_X1 U84046 ( .B1(n113894), .B2(n114144), .A(n120624), .ZN(n114142) );
  OAI21_X1 U84047 ( .B1(n113986), .B2(n114144), .A(n120625), .ZN(n114303) );
  OAI21_X1 U84048 ( .B1(n113894), .B2(n114054), .A(n120623), .ZN(n114052) );
  OAI21_X1 U84049 ( .B1(n113893), .B2(n113986), .A(n120623), .ZN(n113980) );
  OAI21_X1 U84050 ( .B1(n113893), .B2(n113908), .A(n120623), .ZN(n113902) );
  OAI21_X1 U84051 ( .B1(n113893), .B2(n113913), .A(n120623), .ZN(n113911) );
  OAI21_X1 U84052 ( .B1(n113894), .B2(n113901), .A(n120623), .ZN(n113895) );
  BUF_X1 U84053 ( .A(n114658), .Z(n120216) );
  BUF_X1 U84054 ( .A(n116491), .Z(n120018) );
  BUF_X1 U84055 ( .A(n116491), .Z(n120021) );
  BUF_X1 U84056 ( .A(n116491), .Z(n120019) );
  BUF_X1 U84057 ( .A(n116491), .Z(n120020) );
  BUF_X1 U84058 ( .A(n114658), .Z(n120219) );
  BUF_X1 U84059 ( .A(n114658), .Z(n120218) );
  BUF_X1 U84060 ( .A(n114658), .Z(n120217) );
  NAND2_X1 U84061 ( .A1(n116457), .A2(n116463), .ZN(n114697) );
  NAND2_X1 U84062 ( .A1(n116453), .A2(n116446), .ZN(n114660) );
  NAND2_X1 U84063 ( .A1(n116453), .A2(n116463), .ZN(n114673) );
  NAND2_X1 U84064 ( .A1(n116453), .A2(n116464), .ZN(n114702) );
  NAND2_X1 U84065 ( .A1(n117948), .A2(n117959), .ZN(n116532) );
  NAND2_X1 U84066 ( .A1(n117948), .A2(n117968), .ZN(n116526) );
  NAND2_X1 U84067 ( .A1(n117945), .A2(n117959), .ZN(n116500) );
  NAND2_X1 U84068 ( .A1(n117945), .A2(n117961), .ZN(n116516) );
  NAND2_X1 U84069 ( .A1(n117945), .A2(n117968), .ZN(n116531) );
  NAND2_X1 U84070 ( .A1(n117945), .A2(n117962), .ZN(n116527) );
  NAND2_X1 U84071 ( .A1(n114375), .A2(n114376), .ZN(n113894) );
  NAND2_X1 U84072 ( .A1(n116445), .A2(n116459), .ZN(n114687) );
  BUF_X1 U84073 ( .A(n113892), .Z(n120624) );
  BUF_X1 U84074 ( .A(n113892), .Z(n120623) );
  BUF_X1 U84075 ( .A(n113892), .Z(n120625) );
  BUF_X1 U84076 ( .A(n113892), .Z(n120627) );
  BUF_X1 U84077 ( .A(n113892), .Z(n120626) );
  NAND2_X1 U84078 ( .A1(n116453), .A2(n116448), .ZN(n114659) );
  NAND2_X1 U84079 ( .A1(n116453), .A2(n116459), .ZN(n114666) );
  NAND2_X1 U84080 ( .A1(n116454), .A2(n116457), .ZN(n114685) );
  NAND2_X1 U84081 ( .A1(n116448), .A2(n116457), .ZN(n114686) );
  NAND2_X1 U84082 ( .A1(n116464), .A2(n116457), .ZN(n114696) );
  NAND2_X1 U84083 ( .A1(n116457), .A2(n116459), .ZN(n114688) );
  NAND2_X1 U84084 ( .A1(n116458), .A2(n116453), .ZN(n114667) );
  NAND2_X1 U84085 ( .A1(n116452), .A2(n116453), .ZN(n114682) );
  NAND2_X1 U84086 ( .A1(n117947), .A2(n117948), .ZN(n116488) );
  NAND2_X1 U84087 ( .A1(n117946), .A2(n117948), .ZN(n116505) );
  NAND2_X1 U84088 ( .A1(n117962), .A2(n117948), .ZN(n116515) );
  NAND2_X1 U84089 ( .A1(n117955), .A2(n117945), .ZN(n116493) );
  NAND2_X1 U84090 ( .A1(n117948), .A2(n117961), .ZN(n116521) );
  NAND2_X1 U84091 ( .A1(n117946), .A2(n117953), .ZN(n116517) );
  NAND2_X1 U84092 ( .A1(n117953), .A2(n117968), .ZN(n116519) );
  OAI22_X1 U84093 ( .A1(n113907), .A2(n120053), .B1(n114582), .B2(n120047), 
        .ZN(n114781) );
  OAI22_X1 U84094 ( .A1(n113906), .A2(n120053), .B1(n114581), .B2(n120047), 
        .ZN(n114755) );
  OAI22_X1 U84095 ( .A1(n113905), .A2(n120053), .B1(n114580), .B2(n120047), 
        .ZN(n114729) );
  OAI22_X1 U84096 ( .A1(n113903), .A2(n120053), .B1(n114578), .B2(n120047), 
        .ZN(n114701) );
  NAND2_X1 U84097 ( .A1(n116446), .A2(n116447), .ZN(n114655) );
  NAND2_X1 U84098 ( .A1(n116458), .A2(n116447), .ZN(n114703) );
  NAND2_X1 U84099 ( .A1(n117946), .A2(n117954), .ZN(n116514) );
  NAND2_X1 U84100 ( .A1(n117949), .A2(n117954), .ZN(n116513) );
  NAND2_X1 U84101 ( .A1(n117962), .A2(n117954), .ZN(n116518) );
  NAND2_X1 U84102 ( .A1(n116448), .A2(n116445), .ZN(n114684) );
  NAND2_X1 U84103 ( .A1(n117954), .A2(n117959), .ZN(n116520) );
  NAND2_X1 U84104 ( .A1(n116464), .A2(n116445), .ZN(n114683) );
  BUF_X1 U84105 ( .A(n113891), .Z(n120630) );
  BUF_X1 U84106 ( .A(n113889), .Z(n120633) );
  BUF_X1 U84107 ( .A(n113887), .Z(n120636) );
  BUF_X1 U84108 ( .A(n113885), .Z(n120639) );
  BUF_X1 U84109 ( .A(n113883), .Z(n120642) );
  BUF_X1 U84110 ( .A(n113881), .Z(n120645) );
  BUF_X1 U84111 ( .A(n113879), .Z(n120648) );
  BUF_X1 U84112 ( .A(n113877), .Z(n120651) );
  BUF_X1 U84113 ( .A(n113875), .Z(n120654) );
  BUF_X1 U84114 ( .A(n113873), .Z(n120657) );
  BUF_X1 U84115 ( .A(n113871), .Z(n120660) );
  BUF_X1 U84116 ( .A(n113869), .Z(n120663) );
  BUF_X1 U84117 ( .A(n113867), .Z(n120666) );
  BUF_X1 U84118 ( .A(n113865), .Z(n120669) );
  BUF_X1 U84119 ( .A(n113863), .Z(n120672) );
  BUF_X1 U84120 ( .A(n113861), .Z(n120675) );
  BUF_X1 U84121 ( .A(n113859), .Z(n120678) );
  BUF_X1 U84122 ( .A(n113857), .Z(n120681) );
  BUF_X1 U84123 ( .A(n113855), .Z(n120684) );
  BUF_X1 U84124 ( .A(n113853), .Z(n120687) );
  BUF_X1 U84125 ( .A(n113851), .Z(n120690) );
  BUF_X1 U84126 ( .A(n113849), .Z(n120693) );
  BUF_X1 U84127 ( .A(n113847), .Z(n120696) );
  BUF_X1 U84128 ( .A(n113845), .Z(n120699) );
  BUF_X1 U84129 ( .A(n113843), .Z(n120702) );
  BUF_X1 U84130 ( .A(n113841), .Z(n120705) );
  BUF_X1 U84131 ( .A(n113839), .Z(n120708) );
  BUF_X1 U84132 ( .A(n113837), .Z(n120711) );
  BUF_X1 U84133 ( .A(n113835), .Z(n120714) );
  BUF_X1 U84134 ( .A(n113833), .Z(n120717) );
  BUF_X1 U84135 ( .A(n113831), .Z(n120720) );
  BUF_X1 U84136 ( .A(n113829), .Z(n120723) );
  BUF_X1 U84137 ( .A(n113827), .Z(n120726) );
  BUF_X1 U84138 ( .A(n113825), .Z(n120729) );
  BUF_X1 U84139 ( .A(n113823), .Z(n120732) );
  BUF_X1 U84140 ( .A(n113821), .Z(n120735) );
  BUF_X1 U84141 ( .A(n113819), .Z(n120738) );
  BUF_X1 U84142 ( .A(n113817), .Z(n120741) );
  BUF_X1 U84143 ( .A(n113815), .Z(n120744) );
  BUF_X1 U84144 ( .A(n113813), .Z(n120747) );
  BUF_X1 U84145 ( .A(n113811), .Z(n120750) );
  BUF_X1 U84146 ( .A(n113809), .Z(n120753) );
  BUF_X1 U84147 ( .A(n113807), .Z(n120756) );
  BUF_X1 U84148 ( .A(n113805), .Z(n120759) );
  BUF_X1 U84149 ( .A(n113803), .Z(n120762) );
  BUF_X1 U84150 ( .A(n113801), .Z(n120765) );
  BUF_X1 U84151 ( .A(n113799), .Z(n120768) );
  BUF_X1 U84152 ( .A(n113797), .Z(n120771) );
  BUF_X1 U84153 ( .A(n113795), .Z(n120774) );
  BUF_X1 U84154 ( .A(n113793), .Z(n120777) );
  BUF_X1 U84155 ( .A(n113791), .Z(n120780) );
  BUF_X1 U84156 ( .A(n113789), .Z(n120783) );
  BUF_X1 U84157 ( .A(n113787), .Z(n120786) );
  BUF_X1 U84158 ( .A(n113785), .Z(n120789) );
  BUF_X1 U84159 ( .A(n113783), .Z(n120792) );
  BUF_X1 U84160 ( .A(n113781), .Z(n120795) );
  BUF_X1 U84161 ( .A(n113779), .Z(n120798) );
  BUF_X1 U84162 ( .A(n113777), .Z(n120801) );
  BUF_X1 U84163 ( .A(n113775), .Z(n120804) );
  BUF_X1 U84164 ( .A(n113773), .Z(n120807) );
  BUF_X1 U84165 ( .A(n113771), .Z(n120810) );
  BUF_X1 U84166 ( .A(n113770), .Z(n120813) );
  BUF_X1 U84167 ( .A(n113769), .Z(n120816) );
  BUF_X1 U84168 ( .A(n113768), .Z(n120819) );
  BUF_X1 U84169 ( .A(n116491), .Z(n120022) );
  BUF_X1 U84170 ( .A(n114658), .Z(n120220) );
  BUF_X1 U84171 ( .A(n113771), .Z(n120809) );
  BUF_X1 U84172 ( .A(n113770), .Z(n120812) );
  BUF_X1 U84173 ( .A(n113769), .Z(n120815) );
  BUF_X1 U84174 ( .A(n113768), .Z(n120818) );
  BUF_X1 U84175 ( .A(n113891), .Z(n120629) );
  BUF_X1 U84176 ( .A(n113889), .Z(n120632) );
  BUF_X1 U84177 ( .A(n113887), .Z(n120635) );
  BUF_X1 U84178 ( .A(n113885), .Z(n120638) );
  BUF_X1 U84179 ( .A(n113883), .Z(n120641) );
  BUF_X1 U84180 ( .A(n113881), .Z(n120644) );
  BUF_X1 U84181 ( .A(n113879), .Z(n120647) );
  BUF_X1 U84182 ( .A(n113877), .Z(n120650) );
  BUF_X1 U84183 ( .A(n113875), .Z(n120653) );
  BUF_X1 U84184 ( .A(n113873), .Z(n120656) );
  BUF_X1 U84185 ( .A(n113871), .Z(n120659) );
  BUF_X1 U84186 ( .A(n113869), .Z(n120662) );
  BUF_X1 U84187 ( .A(n113867), .Z(n120665) );
  BUF_X1 U84188 ( .A(n113865), .Z(n120668) );
  BUF_X1 U84189 ( .A(n113863), .Z(n120671) );
  BUF_X1 U84190 ( .A(n113861), .Z(n120674) );
  BUF_X1 U84191 ( .A(n113859), .Z(n120677) );
  BUF_X1 U84192 ( .A(n113857), .Z(n120680) );
  BUF_X1 U84193 ( .A(n113855), .Z(n120683) );
  BUF_X1 U84194 ( .A(n113853), .Z(n120686) );
  BUF_X1 U84195 ( .A(n113851), .Z(n120689) );
  BUF_X1 U84196 ( .A(n113849), .Z(n120692) );
  BUF_X1 U84197 ( .A(n113847), .Z(n120695) );
  BUF_X1 U84198 ( .A(n113845), .Z(n120698) );
  BUF_X1 U84199 ( .A(n113843), .Z(n120701) );
  BUF_X1 U84200 ( .A(n113841), .Z(n120704) );
  BUF_X1 U84201 ( .A(n113839), .Z(n120707) );
  BUF_X1 U84202 ( .A(n113837), .Z(n120710) );
  BUF_X1 U84203 ( .A(n113835), .Z(n120713) );
  BUF_X1 U84204 ( .A(n113833), .Z(n120716) );
  BUF_X1 U84205 ( .A(n113831), .Z(n120719) );
  BUF_X1 U84206 ( .A(n113829), .Z(n120722) );
  BUF_X1 U84207 ( .A(n113827), .Z(n120725) );
  BUF_X1 U84208 ( .A(n113825), .Z(n120728) );
  BUF_X1 U84209 ( .A(n113823), .Z(n120731) );
  BUF_X1 U84210 ( .A(n113821), .Z(n120734) );
  BUF_X1 U84211 ( .A(n113819), .Z(n120737) );
  BUF_X1 U84212 ( .A(n113817), .Z(n120740) );
  BUF_X1 U84213 ( .A(n113815), .Z(n120743) );
  BUF_X1 U84214 ( .A(n113813), .Z(n120746) );
  BUF_X1 U84215 ( .A(n113811), .Z(n120749) );
  BUF_X1 U84216 ( .A(n113809), .Z(n120752) );
  BUF_X1 U84217 ( .A(n113807), .Z(n120755) );
  BUF_X1 U84218 ( .A(n113805), .Z(n120758) );
  BUF_X1 U84219 ( .A(n113803), .Z(n120761) );
  BUF_X1 U84220 ( .A(n113801), .Z(n120764) );
  BUF_X1 U84221 ( .A(n113799), .Z(n120767) );
  BUF_X1 U84222 ( .A(n113797), .Z(n120770) );
  BUF_X1 U84223 ( .A(n113795), .Z(n120773) );
  BUF_X1 U84224 ( .A(n113793), .Z(n120776) );
  BUF_X1 U84225 ( .A(n113791), .Z(n120779) );
  BUF_X1 U84226 ( .A(n113789), .Z(n120782) );
  BUF_X1 U84227 ( .A(n113787), .Z(n120785) );
  BUF_X1 U84228 ( .A(n113785), .Z(n120788) );
  BUF_X1 U84229 ( .A(n113783), .Z(n120791) );
  BUF_X1 U84230 ( .A(n113781), .Z(n120794) );
  BUF_X1 U84231 ( .A(n113779), .Z(n120797) );
  BUF_X1 U84232 ( .A(n113777), .Z(n120800) );
  BUF_X1 U84233 ( .A(n113775), .Z(n120803) );
  BUF_X1 U84234 ( .A(n113773), .Z(n120806) );
  NAND2_X1 U84235 ( .A1(n116458), .A2(n116457), .ZN(n114672) );
  OAI22_X1 U84236 ( .A1(n120833), .A2(n113866), .B1(n120822), .B2(n120665), 
        .ZN(n7435) );
  OAI22_X1 U84237 ( .A1(n120833), .A2(n113864), .B1(n120822), .B2(n120668), 
        .ZN(n7436) );
  OAI22_X1 U84238 ( .A1(n120832), .A2(n113862), .B1(n120822), .B2(n120671), 
        .ZN(n7437) );
  OAI22_X1 U84239 ( .A1(n120832), .A2(n113860), .B1(n120822), .B2(n120674), 
        .ZN(n7438) );
  OAI22_X1 U84240 ( .A1(n120832), .A2(n113858), .B1(n120822), .B2(n120677), 
        .ZN(n7439) );
  OAI22_X1 U84241 ( .A1(n120832), .A2(n113856), .B1(n120822), .B2(n120680), 
        .ZN(n7440) );
  OAI22_X1 U84242 ( .A1(n120832), .A2(n113854), .B1(n120822), .B2(n120683), 
        .ZN(n7441) );
  OAI22_X1 U84243 ( .A1(n120832), .A2(n113852), .B1(n120822), .B2(n120686), 
        .ZN(n7442) );
  OAI22_X1 U84244 ( .A1(n120832), .A2(n113850), .B1(n120822), .B2(n120689), 
        .ZN(n7443) );
  OAI22_X1 U84245 ( .A1(n120832), .A2(n113848), .B1(n120822), .B2(n120692), 
        .ZN(n7444) );
  OAI22_X1 U84246 ( .A1(n120832), .A2(n113846), .B1(n120822), .B2(n120695), 
        .ZN(n7445) );
  OAI22_X1 U84247 ( .A1(n120832), .A2(n113844), .B1(n120822), .B2(n120698), 
        .ZN(n7446) );
  OAI22_X1 U84248 ( .A1(n120832), .A2(n113842), .B1(n120823), .B2(n120701), 
        .ZN(n7447) );
  OAI22_X1 U84249 ( .A1(n120832), .A2(n113840), .B1(n120823), .B2(n120704), 
        .ZN(n7448) );
  OAI22_X1 U84250 ( .A1(n120832), .A2(n113838), .B1(n120823), .B2(n120707), 
        .ZN(n7449) );
  OAI22_X1 U84251 ( .A1(n120831), .A2(n113836), .B1(n120823), .B2(n120710), 
        .ZN(n7450) );
  OAI22_X1 U84252 ( .A1(n120831), .A2(n113834), .B1(n120823), .B2(n120713), 
        .ZN(n7451) );
  OAI22_X1 U84253 ( .A1(n120831), .A2(n113832), .B1(n120823), .B2(n120716), 
        .ZN(n7452) );
  OAI22_X1 U84254 ( .A1(n120831), .A2(n113830), .B1(n120823), .B2(n120719), 
        .ZN(n7453) );
  OAI22_X1 U84255 ( .A1(n120831), .A2(n113828), .B1(n120823), .B2(n120722), 
        .ZN(n7454) );
  OAI22_X1 U84256 ( .A1(n120831), .A2(n113826), .B1(n120823), .B2(n120725), 
        .ZN(n7455) );
  OAI22_X1 U84257 ( .A1(n120831), .A2(n113824), .B1(n120823), .B2(n120728), 
        .ZN(n7456) );
  OAI22_X1 U84258 ( .A1(n120831), .A2(n113822), .B1(n120823), .B2(n120731), 
        .ZN(n7457) );
  OAI22_X1 U84259 ( .A1(n120831), .A2(n113820), .B1(n120823), .B2(n120734), 
        .ZN(n7458) );
  OAI22_X1 U84260 ( .A1(n120831), .A2(n113818), .B1(n120824), .B2(n120737), 
        .ZN(n7459) );
  OAI22_X1 U84261 ( .A1(n120831), .A2(n113816), .B1(n120824), .B2(n120740), 
        .ZN(n7460) );
  OAI22_X1 U84262 ( .A1(n120831), .A2(n113814), .B1(n120824), .B2(n120743), 
        .ZN(n7461) );
  OAI22_X1 U84263 ( .A1(n120830), .A2(n113812), .B1(n120824), .B2(n120746), 
        .ZN(n7462) );
  OAI22_X1 U84264 ( .A1(n120830), .A2(n113810), .B1(n120824), .B2(n120749), 
        .ZN(n7463) );
  OAI22_X1 U84265 ( .A1(n120830), .A2(n113808), .B1(n120824), .B2(n120752), 
        .ZN(n7464) );
  OAI22_X1 U84266 ( .A1(n120830), .A2(n113806), .B1(n120824), .B2(n120755), 
        .ZN(n7465) );
  OAI22_X1 U84267 ( .A1(n120830), .A2(n113804), .B1(n120824), .B2(n120758), 
        .ZN(n7466) );
  OAI22_X1 U84268 ( .A1(n120830), .A2(n113802), .B1(n120824), .B2(n120761), 
        .ZN(n7467) );
  OAI22_X1 U84269 ( .A1(n120830), .A2(n113800), .B1(n120824), .B2(n120764), 
        .ZN(n7468) );
  OAI22_X1 U84270 ( .A1(n120830), .A2(n113798), .B1(n120824), .B2(n120767), 
        .ZN(n7469) );
  OAI22_X1 U84271 ( .A1(n120831), .A2(n113796), .B1(n120824), .B2(n120770), 
        .ZN(n7470) );
  OAI22_X1 U84272 ( .A1(n120830), .A2(n113794), .B1(n120825), .B2(n120773), 
        .ZN(n7471) );
  OAI22_X1 U84273 ( .A1(n120830), .A2(n113792), .B1(n120825), .B2(n120776), 
        .ZN(n7472) );
  OAI22_X1 U84274 ( .A1(n120830), .A2(n113790), .B1(n120825), .B2(n120779), 
        .ZN(n7473) );
  OAI22_X1 U84275 ( .A1(n120830), .A2(n113788), .B1(n120825), .B2(n120782), 
        .ZN(n7474) );
  OAI22_X1 U84276 ( .A1(n120830), .A2(n113786), .B1(n120825), .B2(n120785), 
        .ZN(n7475) );
  OAI22_X1 U84277 ( .A1(n120829), .A2(n113784), .B1(n120825), .B2(n120788), 
        .ZN(n7476) );
  OAI22_X1 U84278 ( .A1(n120829), .A2(n113782), .B1(n120825), .B2(n120791), 
        .ZN(n7477) );
  OAI22_X1 U84279 ( .A1(n120829), .A2(n113780), .B1(n120825), .B2(n120794), 
        .ZN(n7478) );
  OAI22_X1 U84280 ( .A1(n120829), .A2(n113778), .B1(n120825), .B2(n120797), 
        .ZN(n7479) );
  OAI22_X1 U84281 ( .A1(n120829), .A2(n113776), .B1(n120825), .B2(n120800), 
        .ZN(n7480) );
  OAI22_X1 U84282 ( .A1(n120829), .A2(n113774), .B1(n120825), .B2(n120803), 
        .ZN(n7481) );
  OAI22_X1 U84283 ( .A1(n120829), .A2(n113772), .B1(n120825), .B2(n120806), 
        .ZN(n7482) );
  NAND2_X1 U84284 ( .A1(n117949), .A2(n117945), .ZN(n116487) );
  NAND2_X1 U84285 ( .A1(n117949), .A2(n117953), .ZN(n116492) );
  NAND2_X1 U84286 ( .A1(n117955), .A2(n117953), .ZN(n116499) );
  NAND2_X1 U84287 ( .A1(n117961), .A2(n117953), .ZN(n116504) );
  OAI22_X1 U84288 ( .A1(n120511), .A2(n114127), .B1(n120809), .B2(n120505), 
        .ZN(n6843) );
  OAI22_X1 U84289 ( .A1(n120511), .A2(n114126), .B1(n120812), .B2(n120505), 
        .ZN(n6844) );
  OAI22_X1 U84290 ( .A1(n120511), .A2(n114125), .B1(n120815), .B2(n120505), 
        .ZN(n6845) );
  OAI22_X1 U84291 ( .A1(n120511), .A2(n114123), .B1(n120818), .B2(n120505), 
        .ZN(n6846) );
  OAI22_X1 U84292 ( .A1(n120561), .A2(n113985), .B1(n120809), .B2(n120555), 
        .ZN(n7099) );
  OAI22_X1 U84293 ( .A1(n120561), .A2(n113984), .B1(n120812), .B2(n120555), 
        .ZN(n7100) );
  OAI22_X1 U84294 ( .A1(n120561), .A2(n113983), .B1(n120815), .B2(n120555), 
        .ZN(n7101) );
  OAI22_X1 U84295 ( .A1(n120561), .A2(n113981), .B1(n120818), .B2(n120555), 
        .ZN(n7102) );
  OAI22_X1 U84296 ( .A1(n120610), .A2(n113907), .B1(n120809), .B2(n120604), 
        .ZN(n7355) );
  OAI22_X1 U84297 ( .A1(n120610), .A2(n113906), .B1(n120812), .B2(n120604), 
        .ZN(n7356) );
  OAI22_X1 U84298 ( .A1(n120610), .A2(n113905), .B1(n120815), .B2(n120604), 
        .ZN(n7357) );
  OAI22_X1 U84299 ( .A1(n120610), .A2(n113903), .B1(n120818), .B2(n120604), 
        .ZN(n7358) );
  NAND2_X1 U84300 ( .A1(n116446), .A2(n116457), .ZN(n114690) );
  OAI22_X1 U84301 ( .A1(n120252), .A2(n114756), .B1(n120811), .B2(n120245), 
        .ZN(n5496) );
  OAI22_X1 U84302 ( .A1(n120252), .A2(n114730), .B1(n120814), .B2(n120245), 
        .ZN(n5498) );
  OAI22_X1 U84303 ( .A1(n120252), .A2(n114704), .B1(n120817), .B2(n120245), 
        .ZN(n5500) );
  OAI22_X1 U84304 ( .A1(n120252), .A2(n114644), .B1(n120820), .B2(n120245), 
        .ZN(n5502) );
  OAI22_X1 U84305 ( .A1(n120574), .A2(n113919), .B1(n120809), .B2(n120567), 
        .ZN(n7163) );
  OAI22_X1 U84306 ( .A1(n120574), .A2(n113918), .B1(n120812), .B2(n120567), 
        .ZN(n7164) );
  OAI22_X1 U84307 ( .A1(n120574), .A2(n113917), .B1(n120815), .B2(n120567), 
        .ZN(n7165) );
  OAI22_X1 U84308 ( .A1(n120574), .A2(n113915), .B1(n120818), .B2(n120567), 
        .ZN(n7166) );
  OAI22_X1 U84309 ( .A1(n120378), .A2(n114239), .B1(n120810), .B2(n120371), 
        .ZN(n6139) );
  OAI22_X1 U84310 ( .A1(n120378), .A2(n114238), .B1(n120813), .B2(n120371), 
        .ZN(n6140) );
  OAI22_X1 U84311 ( .A1(n120378), .A2(n114237), .B1(n120816), .B2(n120371), 
        .ZN(n6141) );
  OAI22_X1 U84312 ( .A1(n120378), .A2(n114235), .B1(n120819), .B2(n120371), 
        .ZN(n6142) );
  OAI22_X1 U84313 ( .A1(n120290), .A2(n114514), .B1(n120811), .B2(n120283), 
        .ZN(n5691) );
  OAI22_X1 U84314 ( .A1(n120290), .A2(n114513), .B1(n120814), .B2(n120283), 
        .ZN(n5692) );
  OAI22_X1 U84315 ( .A1(n120290), .A2(n114512), .B1(n120817), .B2(n120283), 
        .ZN(n5693) );
  OAI22_X1 U84316 ( .A1(n120290), .A2(n114510), .B1(n120820), .B2(n120283), 
        .ZN(n5694) );
  OAI22_X1 U84317 ( .A1(n120265), .A2(n114582), .B1(n120811), .B2(n120258), 
        .ZN(n5563) );
  OAI22_X1 U84318 ( .A1(n120265), .A2(n114581), .B1(n120814), .B2(n120258), 
        .ZN(n5564) );
  OAI22_X1 U84319 ( .A1(n120265), .A2(n114580), .B1(n120817), .B2(n120258), 
        .ZN(n5565) );
  OAI22_X1 U84320 ( .A1(n120265), .A2(n114578), .B1(n120820), .B2(n120258), 
        .ZN(n5566) );
  OAI22_X1 U84321 ( .A1(n120415), .A2(n114150), .B1(n120810), .B2(n120408), 
        .ZN(n6331) );
  OAI22_X1 U84322 ( .A1(n120415), .A2(n114149), .B1(n120813), .B2(n120408), 
        .ZN(n6332) );
  OAI22_X1 U84323 ( .A1(n120415), .A2(n114148), .B1(n120816), .B2(n120408), 
        .ZN(n6333) );
  OAI22_X1 U84324 ( .A1(n120415), .A2(n114146), .B1(n120819), .B2(n120408), 
        .ZN(n6334) );
  OAI22_X1 U84325 ( .A1(n120316), .A2(n114382), .B1(n120811), .B2(n120309), 
        .ZN(n5819) );
  OAI22_X1 U84326 ( .A1(n120316), .A2(n114381), .B1(n120814), .B2(n120309), 
        .ZN(n5820) );
  OAI22_X1 U84327 ( .A1(n120316), .A2(n114380), .B1(n120817), .B2(n120309), 
        .ZN(n5821) );
  OAI22_X1 U84328 ( .A1(n120316), .A2(n114378), .B1(n120820), .B2(n120309), 
        .ZN(n5822) );
  OAI22_X1 U84329 ( .A1(n120303), .A2(n114448), .B1(n120811), .B2(n120296), 
        .ZN(n5755) );
  OAI22_X1 U84330 ( .A1(n120303), .A2(n114447), .B1(n120814), .B2(n120296), 
        .ZN(n5756) );
  OAI22_X1 U84331 ( .A1(n120303), .A2(n114446), .B1(n120817), .B2(n120296), 
        .ZN(n5757) );
  OAI22_X1 U84332 ( .A1(n120303), .A2(n114444), .B1(n120820), .B2(n120296), 
        .ZN(n5758) );
  NAND2_X1 U84333 ( .A1(n116448), .A2(n116447), .ZN(n114654) );
  OAI22_X1 U84334 ( .A1(n120248), .A2(n116434), .B1(n120631), .B2(n120240), 
        .ZN(n5376) );
  OAI22_X1 U84335 ( .A1(n120248), .A2(n116406), .B1(n120634), .B2(n120240), 
        .ZN(n5378) );
  OAI22_X1 U84336 ( .A1(n120248), .A2(n116378), .B1(n120637), .B2(n120240), 
        .ZN(n5380) );
  OAI22_X1 U84337 ( .A1(n120248), .A2(n116350), .B1(n120640), .B2(n120240), 
        .ZN(n5382) );
  OAI22_X1 U84338 ( .A1(n120248), .A2(n116322), .B1(n120643), .B2(n120240), 
        .ZN(n5384) );
  OAI22_X1 U84339 ( .A1(n120248), .A2(n116294), .B1(n120646), .B2(n120240), 
        .ZN(n5386) );
  OAI22_X1 U84340 ( .A1(n120248), .A2(n116266), .B1(n120649), .B2(n120240), 
        .ZN(n5388) );
  OAI22_X1 U84341 ( .A1(n120248), .A2(n116238), .B1(n120652), .B2(n120240), 
        .ZN(n5390) );
  OAI22_X1 U84342 ( .A1(n120248), .A2(n116210), .B1(n120655), .B2(n120240), 
        .ZN(n5392) );
  OAI22_X1 U84343 ( .A1(n120248), .A2(n116182), .B1(n120658), .B2(n120240), 
        .ZN(n5394) );
  OAI22_X1 U84344 ( .A1(n120248), .A2(n116154), .B1(n120661), .B2(n120240), 
        .ZN(n5396) );
  OAI22_X1 U84345 ( .A1(n120248), .A2(n116126), .B1(n120664), .B2(n120240), 
        .ZN(n5398) );
  OAI22_X1 U84346 ( .A1(n120249), .A2(n116098), .B1(n120667), .B2(n120241), 
        .ZN(n5400) );
  OAI22_X1 U84347 ( .A1(n120249), .A2(n116070), .B1(n120670), .B2(n120241), 
        .ZN(n5402) );
  OAI22_X1 U84348 ( .A1(n120249), .A2(n116042), .B1(n120673), .B2(n120241), 
        .ZN(n5404) );
  OAI22_X1 U84349 ( .A1(n120249), .A2(n116014), .B1(n120676), .B2(n120241), 
        .ZN(n5406) );
  OAI22_X1 U84350 ( .A1(n120249), .A2(n115986), .B1(n120679), .B2(n120241), 
        .ZN(n5408) );
  OAI22_X1 U84351 ( .A1(n120249), .A2(n115958), .B1(n120682), .B2(n120241), 
        .ZN(n5410) );
  OAI22_X1 U84352 ( .A1(n120249), .A2(n115930), .B1(n120685), .B2(n120241), 
        .ZN(n5412) );
  OAI22_X1 U84353 ( .A1(n120249), .A2(n115902), .B1(n120688), .B2(n120241), 
        .ZN(n5414) );
  OAI22_X1 U84354 ( .A1(n120249), .A2(n115874), .B1(n120691), .B2(n120241), 
        .ZN(n5416) );
  OAI22_X1 U84355 ( .A1(n120249), .A2(n115846), .B1(n120694), .B2(n120241), 
        .ZN(n5418) );
  OAI22_X1 U84356 ( .A1(n120249), .A2(n115818), .B1(n120697), .B2(n120241), 
        .ZN(n5420) );
  OAI22_X1 U84357 ( .A1(n120249), .A2(n115790), .B1(n120700), .B2(n120241), 
        .ZN(n5422) );
  OAI22_X1 U84358 ( .A1(n120249), .A2(n115762), .B1(n120703), .B2(n120242), 
        .ZN(n5424) );
  OAI22_X1 U84359 ( .A1(n120250), .A2(n115734), .B1(n120706), .B2(n120242), 
        .ZN(n5426) );
  OAI22_X1 U84360 ( .A1(n120250), .A2(n115706), .B1(n120709), .B2(n120242), 
        .ZN(n5428) );
  OAI22_X1 U84361 ( .A1(n120250), .A2(n115678), .B1(n120712), .B2(n120242), 
        .ZN(n5430) );
  OAI22_X1 U84362 ( .A1(n120250), .A2(n115650), .B1(n120715), .B2(n120242), 
        .ZN(n5432) );
  OAI22_X1 U84363 ( .A1(n120250), .A2(n115622), .B1(n120718), .B2(n120242), 
        .ZN(n5434) );
  OAI22_X1 U84364 ( .A1(n120250), .A2(n115594), .B1(n120721), .B2(n120242), 
        .ZN(n5436) );
  OAI22_X1 U84365 ( .A1(n120250), .A2(n115566), .B1(n120724), .B2(n120242), 
        .ZN(n5438) );
  OAI22_X1 U84366 ( .A1(n120250), .A2(n115538), .B1(n120727), .B2(n120242), 
        .ZN(n5440) );
  OAI22_X1 U84367 ( .A1(n120250), .A2(n115510), .B1(n120730), .B2(n120242), 
        .ZN(n5442) );
  OAI22_X1 U84368 ( .A1(n120250), .A2(n115482), .B1(n120733), .B2(n120242), 
        .ZN(n5444) );
  OAI22_X1 U84369 ( .A1(n120250), .A2(n115454), .B1(n120736), .B2(n120242), 
        .ZN(n5446) );
  OAI22_X1 U84370 ( .A1(n120250), .A2(n115426), .B1(n120739), .B2(n120243), 
        .ZN(n5448) );
  OAI22_X1 U84371 ( .A1(n120250), .A2(n115398), .B1(n120742), .B2(n120243), 
        .ZN(n5450) );
  OAI22_X1 U84372 ( .A1(n120251), .A2(n115370), .B1(n120745), .B2(n120243), 
        .ZN(n5452) );
  OAI22_X1 U84373 ( .A1(n120251), .A2(n115342), .B1(n120748), .B2(n120243), 
        .ZN(n5454) );
  OAI22_X1 U84374 ( .A1(n120251), .A2(n115314), .B1(n120751), .B2(n120243), 
        .ZN(n5456) );
  OAI22_X1 U84375 ( .A1(n120251), .A2(n115286), .B1(n120754), .B2(n120243), 
        .ZN(n5458) );
  OAI22_X1 U84376 ( .A1(n120251), .A2(n115258), .B1(n120757), .B2(n120243), 
        .ZN(n5460) );
  OAI22_X1 U84377 ( .A1(n120251), .A2(n115230), .B1(n120760), .B2(n120243), 
        .ZN(n5462) );
  OAI22_X1 U84378 ( .A1(n120251), .A2(n115202), .B1(n120763), .B2(n120243), 
        .ZN(n5464) );
  OAI22_X1 U84379 ( .A1(n120251), .A2(n115174), .B1(n120766), .B2(n120243), 
        .ZN(n5466) );
  OAI22_X1 U84380 ( .A1(n120251), .A2(n115146), .B1(n120769), .B2(n120243), 
        .ZN(n5468) );
  OAI22_X1 U84381 ( .A1(n120251), .A2(n115118), .B1(n120772), .B2(n120243), 
        .ZN(n5470) );
  OAI22_X1 U84382 ( .A1(n120251), .A2(n115090), .B1(n120775), .B2(n120244), 
        .ZN(n5472) );
  OAI22_X1 U84383 ( .A1(n120251), .A2(n115062), .B1(n120778), .B2(n120244), 
        .ZN(n5474) );
  OAI22_X1 U84384 ( .A1(n120251), .A2(n115034), .B1(n120781), .B2(n120244), 
        .ZN(n5476) );
  OAI22_X1 U84385 ( .A1(n120252), .A2(n115006), .B1(n120784), .B2(n120244), 
        .ZN(n5478) );
  OAI22_X1 U84386 ( .A1(n120252), .A2(n114978), .B1(n120787), .B2(n120244), 
        .ZN(n5480) );
  OAI22_X1 U84387 ( .A1(n120252), .A2(n114950), .B1(n120790), .B2(n120244), 
        .ZN(n5482) );
  OAI22_X1 U84388 ( .A1(n120252), .A2(n114922), .B1(n120793), .B2(n120244), 
        .ZN(n5484) );
  OAI22_X1 U84389 ( .A1(n120252), .A2(n114894), .B1(n120796), .B2(n120244), 
        .ZN(n5486) );
  OAI22_X1 U84390 ( .A1(n120252), .A2(n114866), .B1(n120799), .B2(n120244), 
        .ZN(n5488) );
  OAI22_X1 U84391 ( .A1(n120252), .A2(n114838), .B1(n120802), .B2(n120244), 
        .ZN(n5490) );
  OAI22_X1 U84392 ( .A1(n120252), .A2(n114810), .B1(n120805), .B2(n120244), 
        .ZN(n5492) );
  OAI22_X1 U84393 ( .A1(n120252), .A2(n114782), .B1(n120808), .B2(n120244), 
        .ZN(n5494) );
  OAI22_X1 U84394 ( .A1(n120261), .A2(n114642), .B1(n120631), .B2(n120253), 
        .ZN(n5503) );
  OAI22_X1 U84395 ( .A1(n120261), .A2(n114641), .B1(n120634), .B2(n120253), 
        .ZN(n5504) );
  OAI22_X1 U84396 ( .A1(n120261), .A2(n114640), .B1(n120637), .B2(n120253), 
        .ZN(n5505) );
  OAI22_X1 U84397 ( .A1(n120261), .A2(n114639), .B1(n120640), .B2(n120253), 
        .ZN(n5506) );
  OAI22_X1 U84398 ( .A1(n120261), .A2(n114638), .B1(n120643), .B2(n120253), 
        .ZN(n5507) );
  OAI22_X1 U84399 ( .A1(n120261), .A2(n114637), .B1(n120646), .B2(n120253), 
        .ZN(n5508) );
  OAI22_X1 U84400 ( .A1(n120261), .A2(n114636), .B1(n120649), .B2(n120253), 
        .ZN(n5509) );
  OAI22_X1 U84401 ( .A1(n120261), .A2(n114635), .B1(n120652), .B2(n120253), 
        .ZN(n5510) );
  OAI22_X1 U84402 ( .A1(n120261), .A2(n114634), .B1(n120655), .B2(n120253), 
        .ZN(n5511) );
  OAI22_X1 U84403 ( .A1(n120261), .A2(n114633), .B1(n120658), .B2(n120253), 
        .ZN(n5512) );
  OAI22_X1 U84404 ( .A1(n120261), .A2(n114632), .B1(n120661), .B2(n120253), 
        .ZN(n5513) );
  OAI22_X1 U84405 ( .A1(n120261), .A2(n114631), .B1(n120664), .B2(n120253), 
        .ZN(n5514) );
  OAI22_X1 U84406 ( .A1(n120262), .A2(n114630), .B1(n120667), .B2(n120254), 
        .ZN(n5515) );
  OAI22_X1 U84407 ( .A1(n120262), .A2(n114629), .B1(n120670), .B2(n120254), 
        .ZN(n5516) );
  OAI22_X1 U84408 ( .A1(n120262), .A2(n114628), .B1(n120673), .B2(n120254), 
        .ZN(n5517) );
  OAI22_X1 U84409 ( .A1(n120262), .A2(n114627), .B1(n120676), .B2(n120254), 
        .ZN(n5518) );
  OAI22_X1 U84410 ( .A1(n120262), .A2(n114626), .B1(n120679), .B2(n120254), 
        .ZN(n5519) );
  OAI22_X1 U84411 ( .A1(n120262), .A2(n114625), .B1(n120682), .B2(n120254), 
        .ZN(n5520) );
  OAI22_X1 U84412 ( .A1(n120262), .A2(n114624), .B1(n120685), .B2(n120254), 
        .ZN(n5521) );
  OAI22_X1 U84413 ( .A1(n120262), .A2(n114623), .B1(n120688), .B2(n120254), 
        .ZN(n5522) );
  OAI22_X1 U84414 ( .A1(n120262), .A2(n114622), .B1(n120691), .B2(n120254), 
        .ZN(n5523) );
  OAI22_X1 U84415 ( .A1(n120262), .A2(n114621), .B1(n120694), .B2(n120254), 
        .ZN(n5524) );
  OAI22_X1 U84416 ( .A1(n120262), .A2(n114620), .B1(n120697), .B2(n120254), 
        .ZN(n5525) );
  OAI22_X1 U84417 ( .A1(n120262), .A2(n114619), .B1(n120700), .B2(n120254), 
        .ZN(n5526) );
  OAI22_X1 U84418 ( .A1(n120262), .A2(n114618), .B1(n120703), .B2(n120255), 
        .ZN(n5527) );
  OAI22_X1 U84419 ( .A1(n120263), .A2(n114617), .B1(n120706), .B2(n120255), 
        .ZN(n5528) );
  OAI22_X1 U84420 ( .A1(n120263), .A2(n114616), .B1(n120709), .B2(n120255), 
        .ZN(n5529) );
  OAI22_X1 U84421 ( .A1(n120263), .A2(n114615), .B1(n120712), .B2(n120255), 
        .ZN(n5530) );
  OAI22_X1 U84422 ( .A1(n120263), .A2(n114614), .B1(n120715), .B2(n120255), 
        .ZN(n5531) );
  OAI22_X1 U84423 ( .A1(n120263), .A2(n114613), .B1(n120718), .B2(n120255), 
        .ZN(n5532) );
  OAI22_X1 U84424 ( .A1(n120263), .A2(n114612), .B1(n120721), .B2(n120255), 
        .ZN(n5533) );
  OAI22_X1 U84425 ( .A1(n120263), .A2(n114611), .B1(n120724), .B2(n120255), 
        .ZN(n5534) );
  OAI22_X1 U84426 ( .A1(n120263), .A2(n114610), .B1(n120727), .B2(n120255), 
        .ZN(n5535) );
  OAI22_X1 U84427 ( .A1(n120263), .A2(n114609), .B1(n120730), .B2(n120255), 
        .ZN(n5536) );
  OAI22_X1 U84428 ( .A1(n120263), .A2(n114608), .B1(n120733), .B2(n120255), 
        .ZN(n5537) );
  OAI22_X1 U84429 ( .A1(n120263), .A2(n114607), .B1(n120736), .B2(n120255), 
        .ZN(n5538) );
  OAI22_X1 U84430 ( .A1(n120263), .A2(n114606), .B1(n120739), .B2(n120256), 
        .ZN(n5539) );
  OAI22_X1 U84431 ( .A1(n120263), .A2(n114605), .B1(n120742), .B2(n120256), 
        .ZN(n5540) );
  OAI22_X1 U84432 ( .A1(n120264), .A2(n114604), .B1(n120745), .B2(n120256), 
        .ZN(n5541) );
  OAI22_X1 U84433 ( .A1(n120264), .A2(n114603), .B1(n120748), .B2(n120256), 
        .ZN(n5542) );
  OAI22_X1 U84434 ( .A1(n120264), .A2(n114602), .B1(n120751), .B2(n120256), 
        .ZN(n5543) );
  OAI22_X1 U84435 ( .A1(n120264), .A2(n114601), .B1(n120754), .B2(n120256), 
        .ZN(n5544) );
  OAI22_X1 U84436 ( .A1(n120264), .A2(n114600), .B1(n120757), .B2(n120256), 
        .ZN(n5545) );
  OAI22_X1 U84437 ( .A1(n120264), .A2(n114599), .B1(n120760), .B2(n120256), 
        .ZN(n5546) );
  OAI22_X1 U84438 ( .A1(n120264), .A2(n114598), .B1(n120763), .B2(n120256), 
        .ZN(n5547) );
  OAI22_X1 U84439 ( .A1(n120286), .A2(n114574), .B1(n120631), .B2(n120278), 
        .ZN(n5631) );
  OAI22_X1 U84440 ( .A1(n120286), .A2(n114573), .B1(n120634), .B2(n120278), 
        .ZN(n5632) );
  OAI22_X1 U84441 ( .A1(n120286), .A2(n114572), .B1(n120637), .B2(n120278), 
        .ZN(n5633) );
  OAI22_X1 U84442 ( .A1(n120286), .A2(n114571), .B1(n120640), .B2(n120278), 
        .ZN(n5634) );
  OAI22_X1 U84443 ( .A1(n120286), .A2(n114570), .B1(n120643), .B2(n120278), 
        .ZN(n5635) );
  OAI22_X1 U84444 ( .A1(n120286), .A2(n114569), .B1(n120646), .B2(n120278), 
        .ZN(n5636) );
  OAI22_X1 U84445 ( .A1(n120286), .A2(n114568), .B1(n120649), .B2(n120278), 
        .ZN(n5637) );
  OAI22_X1 U84446 ( .A1(n120286), .A2(n114567), .B1(n120652), .B2(n120278), 
        .ZN(n5638) );
  OAI22_X1 U84447 ( .A1(n120286), .A2(n114566), .B1(n120655), .B2(n120278), 
        .ZN(n5639) );
  OAI22_X1 U84448 ( .A1(n120286), .A2(n114565), .B1(n120658), .B2(n120278), 
        .ZN(n5640) );
  OAI22_X1 U84449 ( .A1(n120286), .A2(n114564), .B1(n120661), .B2(n120278), 
        .ZN(n5641) );
  OAI22_X1 U84450 ( .A1(n120286), .A2(n114563), .B1(n120664), .B2(n120278), 
        .ZN(n5642) );
  OAI22_X1 U84451 ( .A1(n120287), .A2(n114562), .B1(n120667), .B2(n120279), 
        .ZN(n5643) );
  OAI22_X1 U84452 ( .A1(n120287), .A2(n114561), .B1(n120670), .B2(n120279), 
        .ZN(n5644) );
  OAI22_X1 U84453 ( .A1(n120287), .A2(n114560), .B1(n120673), .B2(n120279), 
        .ZN(n5645) );
  OAI22_X1 U84454 ( .A1(n120287), .A2(n114559), .B1(n120676), .B2(n120279), 
        .ZN(n5646) );
  OAI22_X1 U84455 ( .A1(n120287), .A2(n114558), .B1(n120679), .B2(n120279), 
        .ZN(n5647) );
  OAI22_X1 U84456 ( .A1(n120287), .A2(n114557), .B1(n120682), .B2(n120279), 
        .ZN(n5648) );
  OAI22_X1 U84457 ( .A1(n120287), .A2(n114556), .B1(n120685), .B2(n120279), 
        .ZN(n5649) );
  OAI22_X1 U84458 ( .A1(n120287), .A2(n114555), .B1(n120688), .B2(n120279), 
        .ZN(n5650) );
  OAI22_X1 U84459 ( .A1(n120287), .A2(n114554), .B1(n120691), .B2(n120279), 
        .ZN(n5651) );
  OAI22_X1 U84460 ( .A1(n120287), .A2(n114553), .B1(n120694), .B2(n120279), 
        .ZN(n5652) );
  OAI22_X1 U84461 ( .A1(n120287), .A2(n114552), .B1(n120697), .B2(n120279), 
        .ZN(n5653) );
  OAI22_X1 U84462 ( .A1(n120287), .A2(n114551), .B1(n120700), .B2(n120279), 
        .ZN(n5654) );
  OAI22_X1 U84463 ( .A1(n120287), .A2(n114550), .B1(n120703), .B2(n120280), 
        .ZN(n5655) );
  OAI22_X1 U84464 ( .A1(n120288), .A2(n114549), .B1(n120706), .B2(n120280), 
        .ZN(n5656) );
  OAI22_X1 U84465 ( .A1(n120288), .A2(n114548), .B1(n120709), .B2(n120280), 
        .ZN(n5657) );
  OAI22_X1 U84466 ( .A1(n120288), .A2(n114547), .B1(n120712), .B2(n120280), 
        .ZN(n5658) );
  OAI22_X1 U84467 ( .A1(n120288), .A2(n114546), .B1(n120715), .B2(n120280), 
        .ZN(n5659) );
  OAI22_X1 U84468 ( .A1(n120288), .A2(n114545), .B1(n120718), .B2(n120280), 
        .ZN(n5660) );
  OAI22_X1 U84469 ( .A1(n120288), .A2(n114544), .B1(n120721), .B2(n120280), 
        .ZN(n5661) );
  OAI22_X1 U84470 ( .A1(n120288), .A2(n114543), .B1(n120724), .B2(n120280), 
        .ZN(n5662) );
  OAI22_X1 U84471 ( .A1(n120288), .A2(n114542), .B1(n120727), .B2(n120280), 
        .ZN(n5663) );
  OAI22_X1 U84472 ( .A1(n120288), .A2(n114541), .B1(n120730), .B2(n120280), 
        .ZN(n5664) );
  OAI22_X1 U84473 ( .A1(n120288), .A2(n114540), .B1(n120733), .B2(n120280), 
        .ZN(n5665) );
  OAI22_X1 U84474 ( .A1(n120288), .A2(n114539), .B1(n120736), .B2(n120280), 
        .ZN(n5666) );
  OAI22_X1 U84475 ( .A1(n120288), .A2(n114538), .B1(n120739), .B2(n120281), 
        .ZN(n5667) );
  OAI22_X1 U84476 ( .A1(n120288), .A2(n114537), .B1(n120742), .B2(n120281), 
        .ZN(n5668) );
  OAI22_X1 U84477 ( .A1(n120289), .A2(n114536), .B1(n120745), .B2(n120281), 
        .ZN(n5669) );
  OAI22_X1 U84478 ( .A1(n120289), .A2(n114535), .B1(n120748), .B2(n120281), 
        .ZN(n5670) );
  OAI22_X1 U84479 ( .A1(n120289), .A2(n114534), .B1(n120751), .B2(n120281), 
        .ZN(n5671) );
  OAI22_X1 U84480 ( .A1(n120289), .A2(n114533), .B1(n120754), .B2(n120281), 
        .ZN(n5672) );
  OAI22_X1 U84481 ( .A1(n120289), .A2(n114532), .B1(n120757), .B2(n120281), 
        .ZN(n5673) );
  OAI22_X1 U84482 ( .A1(n120289), .A2(n114531), .B1(n120760), .B2(n120281), 
        .ZN(n5674) );
  OAI22_X1 U84483 ( .A1(n120289), .A2(n114530), .B1(n120763), .B2(n120281), 
        .ZN(n5675) );
  OAI22_X1 U84484 ( .A1(n120289), .A2(n114529), .B1(n120766), .B2(n120281), 
        .ZN(n5676) );
  OAI22_X1 U84485 ( .A1(n120289), .A2(n114528), .B1(n120769), .B2(n120281), 
        .ZN(n5677) );
  OAI22_X1 U84486 ( .A1(n120289), .A2(n114527), .B1(n120772), .B2(n120281), 
        .ZN(n5678) );
  OAI22_X1 U84487 ( .A1(n120289), .A2(n114526), .B1(n120775), .B2(n120282), 
        .ZN(n5679) );
  OAI22_X1 U84488 ( .A1(n120289), .A2(n114525), .B1(n120778), .B2(n120282), 
        .ZN(n5680) );
  OAI22_X1 U84489 ( .A1(n120289), .A2(n114524), .B1(n120781), .B2(n120282), 
        .ZN(n5681) );
  OAI22_X1 U84490 ( .A1(n120290), .A2(n114523), .B1(n120784), .B2(n120282), 
        .ZN(n5682) );
  OAI22_X1 U84491 ( .A1(n120290), .A2(n114522), .B1(n120787), .B2(n120282), 
        .ZN(n5683) );
  OAI22_X1 U84492 ( .A1(n120290), .A2(n114521), .B1(n120790), .B2(n120282), 
        .ZN(n5684) );
  OAI22_X1 U84493 ( .A1(n120290), .A2(n114520), .B1(n120793), .B2(n120282), 
        .ZN(n5685) );
  OAI22_X1 U84494 ( .A1(n120290), .A2(n114519), .B1(n120796), .B2(n120282), 
        .ZN(n5686) );
  OAI22_X1 U84495 ( .A1(n120290), .A2(n114518), .B1(n120799), .B2(n120282), 
        .ZN(n5687) );
  OAI22_X1 U84496 ( .A1(n120290), .A2(n114517), .B1(n120802), .B2(n120282), 
        .ZN(n5688) );
  OAI22_X1 U84497 ( .A1(n120290), .A2(n114516), .B1(n120805), .B2(n120282), 
        .ZN(n5689) );
  OAI22_X1 U84498 ( .A1(n120290), .A2(n114515), .B1(n120808), .B2(n120282), 
        .ZN(n5690) );
  OAI22_X1 U84499 ( .A1(n120264), .A2(n114597), .B1(n120766), .B2(n120256), 
        .ZN(n5548) );
  OAI22_X1 U84500 ( .A1(n120264), .A2(n114596), .B1(n120769), .B2(n120256), 
        .ZN(n5549) );
  OAI22_X1 U84501 ( .A1(n120264), .A2(n114595), .B1(n120772), .B2(n120256), 
        .ZN(n5550) );
  OAI22_X1 U84502 ( .A1(n120264), .A2(n114594), .B1(n120775), .B2(n120257), 
        .ZN(n5551) );
  OAI22_X1 U84503 ( .A1(n120264), .A2(n114593), .B1(n120778), .B2(n120257), 
        .ZN(n5552) );
  OAI22_X1 U84504 ( .A1(n120264), .A2(n114592), .B1(n120781), .B2(n120257), 
        .ZN(n5553) );
  OAI22_X1 U84505 ( .A1(n120265), .A2(n114591), .B1(n120784), .B2(n120257), 
        .ZN(n5554) );
  OAI22_X1 U84506 ( .A1(n120265), .A2(n114590), .B1(n120787), .B2(n120257), 
        .ZN(n5555) );
  OAI22_X1 U84507 ( .A1(n120265), .A2(n114589), .B1(n120790), .B2(n120257), 
        .ZN(n5556) );
  OAI22_X1 U84508 ( .A1(n120265), .A2(n114588), .B1(n120793), .B2(n120257), 
        .ZN(n5557) );
  OAI22_X1 U84509 ( .A1(n120265), .A2(n114587), .B1(n120796), .B2(n120257), 
        .ZN(n5558) );
  OAI22_X1 U84510 ( .A1(n120265), .A2(n114586), .B1(n120799), .B2(n120257), 
        .ZN(n5559) );
  OAI22_X1 U84511 ( .A1(n120265), .A2(n114585), .B1(n120802), .B2(n120257), 
        .ZN(n5560) );
  OAI22_X1 U84512 ( .A1(n120265), .A2(n114584), .B1(n120805), .B2(n120257), 
        .ZN(n5561) );
  OAI22_X1 U84513 ( .A1(n120265), .A2(n114583), .B1(n120808), .B2(n120257), 
        .ZN(n5562) );
  OAI22_X1 U84514 ( .A1(n120312), .A2(n114442), .B1(n120631), .B2(n120304), 
        .ZN(n5759) );
  OAI22_X1 U84515 ( .A1(n120312), .A2(n114441), .B1(n120634), .B2(n120304), 
        .ZN(n5760) );
  OAI22_X1 U84516 ( .A1(n120312), .A2(n114440), .B1(n120637), .B2(n120304), 
        .ZN(n5761) );
  OAI22_X1 U84517 ( .A1(n120312), .A2(n114439), .B1(n120640), .B2(n120304), 
        .ZN(n5762) );
  OAI22_X1 U84518 ( .A1(n120312), .A2(n114438), .B1(n120643), .B2(n120304), 
        .ZN(n5763) );
  OAI22_X1 U84519 ( .A1(n120312), .A2(n114437), .B1(n120646), .B2(n120304), 
        .ZN(n5764) );
  OAI22_X1 U84520 ( .A1(n120312), .A2(n114436), .B1(n120649), .B2(n120304), 
        .ZN(n5765) );
  OAI22_X1 U84521 ( .A1(n120312), .A2(n114435), .B1(n120652), .B2(n120304), 
        .ZN(n5766) );
  OAI22_X1 U84522 ( .A1(n120312), .A2(n114434), .B1(n120655), .B2(n120304), 
        .ZN(n5767) );
  OAI22_X1 U84523 ( .A1(n120312), .A2(n114433), .B1(n120658), .B2(n120304), 
        .ZN(n5768) );
  OAI22_X1 U84524 ( .A1(n120312), .A2(n114432), .B1(n120661), .B2(n120304), 
        .ZN(n5769) );
  OAI22_X1 U84525 ( .A1(n120312), .A2(n114431), .B1(n120664), .B2(n120304), 
        .ZN(n5770) );
  OAI22_X1 U84526 ( .A1(n120313), .A2(n114430), .B1(n120667), .B2(n120305), 
        .ZN(n5771) );
  OAI22_X1 U84527 ( .A1(n120313), .A2(n114429), .B1(n120670), .B2(n120305), 
        .ZN(n5772) );
  OAI22_X1 U84528 ( .A1(n120313), .A2(n114428), .B1(n120673), .B2(n120305), 
        .ZN(n5773) );
  OAI22_X1 U84529 ( .A1(n120313), .A2(n114427), .B1(n120676), .B2(n120305), 
        .ZN(n5774) );
  OAI22_X1 U84530 ( .A1(n120313), .A2(n114426), .B1(n120679), .B2(n120305), 
        .ZN(n5775) );
  OAI22_X1 U84531 ( .A1(n120313), .A2(n114425), .B1(n120682), .B2(n120305), 
        .ZN(n5776) );
  OAI22_X1 U84532 ( .A1(n120313), .A2(n114424), .B1(n120685), .B2(n120305), 
        .ZN(n5777) );
  OAI22_X1 U84533 ( .A1(n120313), .A2(n114423), .B1(n120688), .B2(n120305), 
        .ZN(n5778) );
  OAI22_X1 U84534 ( .A1(n120313), .A2(n114422), .B1(n120691), .B2(n120305), 
        .ZN(n5779) );
  OAI22_X1 U84535 ( .A1(n120313), .A2(n114421), .B1(n120694), .B2(n120305), 
        .ZN(n5780) );
  OAI22_X1 U84536 ( .A1(n120313), .A2(n114420), .B1(n120697), .B2(n120305), 
        .ZN(n5781) );
  OAI22_X1 U84537 ( .A1(n120313), .A2(n114419), .B1(n120700), .B2(n120305), 
        .ZN(n5782) );
  OAI22_X1 U84538 ( .A1(n120313), .A2(n114418), .B1(n120703), .B2(n120306), 
        .ZN(n5783) );
  OAI22_X1 U84539 ( .A1(n120314), .A2(n114417), .B1(n120706), .B2(n120306), 
        .ZN(n5784) );
  OAI22_X1 U84540 ( .A1(n120314), .A2(n114416), .B1(n120709), .B2(n120306), 
        .ZN(n5785) );
  OAI22_X1 U84541 ( .A1(n120314), .A2(n114415), .B1(n120712), .B2(n120306), 
        .ZN(n5786) );
  OAI22_X1 U84542 ( .A1(n120314), .A2(n114414), .B1(n120715), .B2(n120306), 
        .ZN(n5787) );
  OAI22_X1 U84543 ( .A1(n120314), .A2(n114413), .B1(n120718), .B2(n120306), 
        .ZN(n5788) );
  OAI22_X1 U84544 ( .A1(n120314), .A2(n114412), .B1(n120721), .B2(n120306), 
        .ZN(n5789) );
  OAI22_X1 U84545 ( .A1(n120314), .A2(n114411), .B1(n120724), .B2(n120306), 
        .ZN(n5790) );
  OAI22_X1 U84546 ( .A1(n120314), .A2(n114410), .B1(n120727), .B2(n120306), 
        .ZN(n5791) );
  OAI22_X1 U84547 ( .A1(n120314), .A2(n114409), .B1(n120730), .B2(n120306), 
        .ZN(n5792) );
  OAI22_X1 U84548 ( .A1(n120314), .A2(n114408), .B1(n120733), .B2(n120306), 
        .ZN(n5793) );
  OAI22_X1 U84549 ( .A1(n120314), .A2(n114407), .B1(n120736), .B2(n120306), 
        .ZN(n5794) );
  OAI22_X1 U84550 ( .A1(n120314), .A2(n114406), .B1(n120739), .B2(n120307), 
        .ZN(n5795) );
  OAI22_X1 U84551 ( .A1(n120314), .A2(n114405), .B1(n120742), .B2(n120307), 
        .ZN(n5796) );
  OAI22_X1 U84552 ( .A1(n120315), .A2(n114404), .B1(n120745), .B2(n120307), 
        .ZN(n5797) );
  OAI22_X1 U84553 ( .A1(n120315), .A2(n114403), .B1(n120748), .B2(n120307), 
        .ZN(n5798) );
  OAI22_X1 U84554 ( .A1(n120315), .A2(n114402), .B1(n120751), .B2(n120307), 
        .ZN(n5799) );
  OAI22_X1 U84555 ( .A1(n120315), .A2(n114401), .B1(n120754), .B2(n120307), 
        .ZN(n5800) );
  OAI22_X1 U84556 ( .A1(n120315), .A2(n114400), .B1(n120757), .B2(n120307), 
        .ZN(n5801) );
  OAI22_X1 U84557 ( .A1(n120315), .A2(n114399), .B1(n120760), .B2(n120307), 
        .ZN(n5802) );
  OAI22_X1 U84558 ( .A1(n120315), .A2(n114398), .B1(n120763), .B2(n120307), 
        .ZN(n5803) );
  OAI22_X1 U84559 ( .A1(n120315), .A2(n114397), .B1(n120766), .B2(n120307), 
        .ZN(n5804) );
  OAI22_X1 U84560 ( .A1(n120315), .A2(n114396), .B1(n120769), .B2(n120307), 
        .ZN(n5805) );
  OAI22_X1 U84561 ( .A1(n120315), .A2(n114395), .B1(n120772), .B2(n120307), 
        .ZN(n5806) );
  OAI22_X1 U84562 ( .A1(n120315), .A2(n114394), .B1(n120775), .B2(n120308), 
        .ZN(n5807) );
  OAI22_X1 U84563 ( .A1(n120315), .A2(n114393), .B1(n120778), .B2(n120308), 
        .ZN(n5808) );
  OAI22_X1 U84564 ( .A1(n120315), .A2(n114392), .B1(n120781), .B2(n120308), 
        .ZN(n5809) );
  OAI22_X1 U84565 ( .A1(n120316), .A2(n114391), .B1(n120784), .B2(n120308), 
        .ZN(n5810) );
  OAI22_X1 U84566 ( .A1(n120316), .A2(n114390), .B1(n120787), .B2(n120308), 
        .ZN(n5811) );
  OAI22_X1 U84567 ( .A1(n120316), .A2(n114389), .B1(n120790), .B2(n120308), 
        .ZN(n5812) );
  OAI22_X1 U84568 ( .A1(n120316), .A2(n114388), .B1(n120793), .B2(n120308), 
        .ZN(n5813) );
  OAI22_X1 U84569 ( .A1(n120316), .A2(n114387), .B1(n120796), .B2(n120308), 
        .ZN(n5814) );
  OAI22_X1 U84570 ( .A1(n120316), .A2(n114386), .B1(n120799), .B2(n120308), 
        .ZN(n5815) );
  OAI22_X1 U84571 ( .A1(n120316), .A2(n114385), .B1(n120802), .B2(n120308), 
        .ZN(n5816) );
  OAI22_X1 U84572 ( .A1(n120316), .A2(n114384), .B1(n120805), .B2(n120308), 
        .ZN(n5817) );
  OAI22_X1 U84573 ( .A1(n120299), .A2(n114508), .B1(n120631), .B2(n120291), 
        .ZN(n5695) );
  OAI22_X1 U84574 ( .A1(n120299), .A2(n114507), .B1(n120634), .B2(n120291), 
        .ZN(n5696) );
  OAI22_X1 U84575 ( .A1(n120299), .A2(n114506), .B1(n120637), .B2(n120291), 
        .ZN(n5697) );
  OAI22_X1 U84576 ( .A1(n120299), .A2(n114505), .B1(n120640), .B2(n120291), 
        .ZN(n5698) );
  OAI22_X1 U84577 ( .A1(n120299), .A2(n114504), .B1(n120643), .B2(n120291), 
        .ZN(n5699) );
  OAI22_X1 U84578 ( .A1(n120299), .A2(n114503), .B1(n120646), .B2(n120291), 
        .ZN(n5700) );
  OAI22_X1 U84579 ( .A1(n120299), .A2(n114502), .B1(n120649), .B2(n120291), 
        .ZN(n5701) );
  OAI22_X1 U84580 ( .A1(n120299), .A2(n114501), .B1(n120652), .B2(n120291), 
        .ZN(n5702) );
  OAI22_X1 U84581 ( .A1(n120299), .A2(n114500), .B1(n120655), .B2(n120291), 
        .ZN(n5703) );
  OAI22_X1 U84582 ( .A1(n120299), .A2(n114499), .B1(n120658), .B2(n120291), 
        .ZN(n5704) );
  OAI22_X1 U84583 ( .A1(n120299), .A2(n114498), .B1(n120661), .B2(n120291), 
        .ZN(n5705) );
  OAI22_X1 U84584 ( .A1(n120299), .A2(n114497), .B1(n120664), .B2(n120291), 
        .ZN(n5706) );
  OAI22_X1 U84585 ( .A1(n120300), .A2(n114496), .B1(n120667), .B2(n120292), 
        .ZN(n5707) );
  OAI22_X1 U84586 ( .A1(n120300), .A2(n114495), .B1(n120670), .B2(n120292), 
        .ZN(n5708) );
  OAI22_X1 U84587 ( .A1(n120300), .A2(n114494), .B1(n120673), .B2(n120292), 
        .ZN(n5709) );
  OAI22_X1 U84588 ( .A1(n120300), .A2(n114493), .B1(n120676), .B2(n120292), 
        .ZN(n5710) );
  OAI22_X1 U84589 ( .A1(n120300), .A2(n114492), .B1(n120679), .B2(n120292), 
        .ZN(n5711) );
  OAI22_X1 U84590 ( .A1(n120300), .A2(n114491), .B1(n120682), .B2(n120292), 
        .ZN(n5712) );
  OAI22_X1 U84591 ( .A1(n120300), .A2(n114490), .B1(n120685), .B2(n120292), 
        .ZN(n5713) );
  OAI22_X1 U84592 ( .A1(n120300), .A2(n114489), .B1(n120688), .B2(n120292), 
        .ZN(n5714) );
  OAI22_X1 U84593 ( .A1(n120300), .A2(n114488), .B1(n120691), .B2(n120292), 
        .ZN(n5715) );
  OAI22_X1 U84594 ( .A1(n120300), .A2(n114487), .B1(n120694), .B2(n120292), 
        .ZN(n5716) );
  OAI22_X1 U84595 ( .A1(n120300), .A2(n114486), .B1(n120697), .B2(n120292), 
        .ZN(n5717) );
  OAI22_X1 U84596 ( .A1(n120300), .A2(n114485), .B1(n120700), .B2(n120292), 
        .ZN(n5718) );
  OAI22_X1 U84597 ( .A1(n120300), .A2(n114484), .B1(n120703), .B2(n120293), 
        .ZN(n5719) );
  OAI22_X1 U84598 ( .A1(n120301), .A2(n114483), .B1(n120706), .B2(n120293), 
        .ZN(n5720) );
  OAI22_X1 U84599 ( .A1(n120301), .A2(n114482), .B1(n120709), .B2(n120293), 
        .ZN(n5721) );
  OAI22_X1 U84600 ( .A1(n120301), .A2(n114481), .B1(n120712), .B2(n120293), 
        .ZN(n5722) );
  OAI22_X1 U84601 ( .A1(n120301), .A2(n114480), .B1(n120715), .B2(n120293), 
        .ZN(n5723) );
  OAI22_X1 U84602 ( .A1(n120301), .A2(n114479), .B1(n120718), .B2(n120293), 
        .ZN(n5724) );
  OAI22_X1 U84603 ( .A1(n120301), .A2(n114478), .B1(n120721), .B2(n120293), 
        .ZN(n5725) );
  OAI22_X1 U84604 ( .A1(n120301), .A2(n114477), .B1(n120724), .B2(n120293), 
        .ZN(n5726) );
  OAI22_X1 U84605 ( .A1(n120301), .A2(n114476), .B1(n120727), .B2(n120293), 
        .ZN(n5727) );
  OAI22_X1 U84606 ( .A1(n120301), .A2(n114475), .B1(n120730), .B2(n120293), 
        .ZN(n5728) );
  OAI22_X1 U84607 ( .A1(n120301), .A2(n114474), .B1(n120733), .B2(n120293), 
        .ZN(n5729) );
  OAI22_X1 U84608 ( .A1(n120301), .A2(n114473), .B1(n120736), .B2(n120293), 
        .ZN(n5730) );
  OAI22_X1 U84609 ( .A1(n120301), .A2(n114472), .B1(n120739), .B2(n120294), 
        .ZN(n5731) );
  OAI22_X1 U84610 ( .A1(n120301), .A2(n114471), .B1(n120742), .B2(n120294), 
        .ZN(n5732) );
  OAI22_X1 U84611 ( .A1(n120302), .A2(n114470), .B1(n120745), .B2(n120294), 
        .ZN(n5733) );
  OAI22_X1 U84612 ( .A1(n120302), .A2(n114469), .B1(n120748), .B2(n120294), 
        .ZN(n5734) );
  OAI22_X1 U84613 ( .A1(n120302), .A2(n114468), .B1(n120751), .B2(n120294), 
        .ZN(n5735) );
  OAI22_X1 U84614 ( .A1(n120302), .A2(n114467), .B1(n120754), .B2(n120294), 
        .ZN(n5736) );
  OAI22_X1 U84615 ( .A1(n120302), .A2(n114466), .B1(n120757), .B2(n120294), 
        .ZN(n5737) );
  OAI22_X1 U84616 ( .A1(n120302), .A2(n114465), .B1(n120760), .B2(n120294), 
        .ZN(n5738) );
  OAI22_X1 U84617 ( .A1(n120302), .A2(n114464), .B1(n120763), .B2(n120294), 
        .ZN(n5739) );
  OAI22_X1 U84618 ( .A1(n120302), .A2(n114463), .B1(n120766), .B2(n120294), 
        .ZN(n5740) );
  OAI22_X1 U84619 ( .A1(n120302), .A2(n114462), .B1(n120769), .B2(n120294), 
        .ZN(n5741) );
  OAI22_X1 U84620 ( .A1(n120302), .A2(n114461), .B1(n120772), .B2(n120294), 
        .ZN(n5742) );
  OAI22_X1 U84621 ( .A1(n120302), .A2(n114460), .B1(n120775), .B2(n120295), 
        .ZN(n5743) );
  OAI22_X1 U84622 ( .A1(n120302), .A2(n114459), .B1(n120778), .B2(n120295), 
        .ZN(n5744) );
  OAI22_X1 U84623 ( .A1(n120302), .A2(n114458), .B1(n120781), .B2(n120295), 
        .ZN(n5745) );
  OAI22_X1 U84624 ( .A1(n120303), .A2(n114457), .B1(n120784), .B2(n120295), 
        .ZN(n5746) );
  OAI22_X1 U84625 ( .A1(n120303), .A2(n114456), .B1(n120787), .B2(n120295), 
        .ZN(n5747) );
  OAI22_X1 U84626 ( .A1(n120303), .A2(n114455), .B1(n120790), .B2(n120295), 
        .ZN(n5748) );
  OAI22_X1 U84627 ( .A1(n120303), .A2(n114454), .B1(n120793), .B2(n120295), 
        .ZN(n5749) );
  OAI22_X1 U84628 ( .A1(n120303), .A2(n114453), .B1(n120796), .B2(n120295), 
        .ZN(n5750) );
  OAI22_X1 U84629 ( .A1(n120303), .A2(n114452), .B1(n120799), .B2(n120295), 
        .ZN(n5751) );
  OAI22_X1 U84630 ( .A1(n120303), .A2(n114451), .B1(n120802), .B2(n120295), 
        .ZN(n5752) );
  OAI22_X1 U84631 ( .A1(n120303), .A2(n114450), .B1(n120805), .B2(n120295), 
        .ZN(n5753) );
  OAI22_X1 U84632 ( .A1(n120303), .A2(n114449), .B1(n120808), .B2(n120295), 
        .ZN(n5754) );
  OAI22_X1 U84633 ( .A1(n120316), .A2(n114383), .B1(n120808), .B2(n120308), 
        .ZN(n5818) );
  OAI22_X1 U84634 ( .A1(n120545), .A2(n114051), .B1(n120629), .B2(n120537), 
        .ZN(n6975) );
  OAI22_X1 U84635 ( .A1(n120549), .A2(n114050), .B1(n120632), .B2(n120537), 
        .ZN(n6976) );
  OAI22_X1 U84636 ( .A1(n120549), .A2(n114049), .B1(n120635), .B2(n120537), 
        .ZN(n6977) );
  OAI22_X1 U84637 ( .A1(n120549), .A2(n114048), .B1(n120638), .B2(n120537), 
        .ZN(n6978) );
  OAI22_X1 U84638 ( .A1(n120549), .A2(n114047), .B1(n120641), .B2(n120537), 
        .ZN(n6979) );
  OAI22_X1 U84639 ( .A1(n120549), .A2(n114046), .B1(n120644), .B2(n120537), 
        .ZN(n6980) );
  OAI22_X1 U84640 ( .A1(n120549), .A2(n114045), .B1(n120647), .B2(n120537), 
        .ZN(n6981) );
  OAI22_X1 U84641 ( .A1(n120549), .A2(n114044), .B1(n120650), .B2(n120537), 
        .ZN(n6982) );
  OAI22_X1 U84642 ( .A1(n120549), .A2(n114043), .B1(n120653), .B2(n120537), 
        .ZN(n6983) );
  OAI22_X1 U84643 ( .A1(n120549), .A2(n114042), .B1(n120656), .B2(n120537), 
        .ZN(n6984) );
  OAI22_X1 U84644 ( .A1(n120549), .A2(n114041), .B1(n120659), .B2(n120537), 
        .ZN(n6985) );
  OAI22_X1 U84645 ( .A1(n120549), .A2(n114040), .B1(n120662), .B2(n120537), 
        .ZN(n6986) );
  OAI22_X1 U84646 ( .A1(n120549), .A2(n114039), .B1(n120665), .B2(n120538), 
        .ZN(n6987) );
  OAI22_X1 U84647 ( .A1(n120549), .A2(n114038), .B1(n120668), .B2(n120538), 
        .ZN(n6988) );
  OAI22_X1 U84648 ( .A1(n120548), .A2(n114037), .B1(n120671), .B2(n120538), 
        .ZN(n6989) );
  OAI22_X1 U84649 ( .A1(n120548), .A2(n114036), .B1(n120674), .B2(n120538), 
        .ZN(n6990) );
  OAI22_X1 U84650 ( .A1(n120548), .A2(n114035), .B1(n120677), .B2(n120538), 
        .ZN(n6991) );
  OAI22_X1 U84651 ( .A1(n120548), .A2(n114034), .B1(n120680), .B2(n120538), 
        .ZN(n6992) );
  OAI22_X1 U84652 ( .A1(n120548), .A2(n114033), .B1(n120683), .B2(n120538), 
        .ZN(n6993) );
  OAI22_X1 U84653 ( .A1(n120548), .A2(n114032), .B1(n120686), .B2(n120538), 
        .ZN(n6994) );
  OAI22_X1 U84654 ( .A1(n120548), .A2(n114031), .B1(n120689), .B2(n120538), 
        .ZN(n6995) );
  OAI22_X1 U84655 ( .A1(n120548), .A2(n114030), .B1(n120692), .B2(n120538), 
        .ZN(n6996) );
  OAI22_X1 U84656 ( .A1(n120548), .A2(n114029), .B1(n120695), .B2(n120538), 
        .ZN(n6997) );
  OAI22_X1 U84657 ( .A1(n120548), .A2(n114028), .B1(n120698), .B2(n120538), 
        .ZN(n6998) );
  OAI22_X1 U84658 ( .A1(n120548), .A2(n114027), .B1(n120701), .B2(n120539), 
        .ZN(n6999) );
  OAI22_X1 U84659 ( .A1(n120548), .A2(n114026), .B1(n120704), .B2(n120539), 
        .ZN(n7000) );
  OAI22_X1 U84660 ( .A1(n120548), .A2(n114025), .B1(n120707), .B2(n120539), 
        .ZN(n7001) );
  OAI22_X1 U84661 ( .A1(n120547), .A2(n114024), .B1(n120710), .B2(n120539), 
        .ZN(n7002) );
  OAI22_X1 U84662 ( .A1(n120547), .A2(n114023), .B1(n120713), .B2(n120539), 
        .ZN(n7003) );
  OAI22_X1 U84663 ( .A1(n120547), .A2(n114022), .B1(n120716), .B2(n120539), 
        .ZN(n7004) );
  OAI22_X1 U84664 ( .A1(n120547), .A2(n114021), .B1(n120719), .B2(n120539), 
        .ZN(n7005) );
  OAI22_X1 U84665 ( .A1(n120547), .A2(n114020), .B1(n120722), .B2(n120539), 
        .ZN(n7006) );
  OAI22_X1 U84666 ( .A1(n120547), .A2(n114019), .B1(n120725), .B2(n120539), 
        .ZN(n7007) );
  OAI22_X1 U84667 ( .A1(n120547), .A2(n114018), .B1(n120728), .B2(n120539), 
        .ZN(n7008) );
  OAI22_X1 U84668 ( .A1(n120547), .A2(n114017), .B1(n120731), .B2(n120539), 
        .ZN(n7009) );
  OAI22_X1 U84669 ( .A1(n120547), .A2(n114016), .B1(n120734), .B2(n120539), 
        .ZN(n7010) );
  OAI22_X1 U84670 ( .A1(n120547), .A2(n114015), .B1(n120737), .B2(n120540), 
        .ZN(n7011) );
  OAI22_X1 U84671 ( .A1(n120547), .A2(n114014), .B1(n120740), .B2(n120540), 
        .ZN(n7012) );
  OAI22_X1 U84672 ( .A1(n120547), .A2(n114013), .B1(n120743), .B2(n120540), 
        .ZN(n7013) );
  OAI22_X1 U84673 ( .A1(n120546), .A2(n114012), .B1(n120746), .B2(n120540), 
        .ZN(n7014) );
  OAI22_X1 U84674 ( .A1(n120546), .A2(n114011), .B1(n120749), .B2(n120540), 
        .ZN(n7015) );
  OAI22_X1 U84675 ( .A1(n120546), .A2(n114010), .B1(n120752), .B2(n120540), 
        .ZN(n7016) );
  OAI22_X1 U84676 ( .A1(n120546), .A2(n114009), .B1(n120755), .B2(n120540), 
        .ZN(n7017) );
  OAI22_X1 U84677 ( .A1(n120546), .A2(n114008), .B1(n120758), .B2(n120540), 
        .ZN(n7018) );
  OAI22_X1 U84678 ( .A1(n120546), .A2(n114007), .B1(n120761), .B2(n120540), 
        .ZN(n7019) );
  OAI22_X1 U84679 ( .A1(n120546), .A2(n114006), .B1(n120764), .B2(n120540), 
        .ZN(n7020) );
  OAI22_X1 U84680 ( .A1(n120546), .A2(n114005), .B1(n120767), .B2(n120540), 
        .ZN(n7021) );
  OAI22_X1 U84681 ( .A1(n120547), .A2(n114004), .B1(n120770), .B2(n120540), 
        .ZN(n7022) );
  OAI22_X1 U84682 ( .A1(n120546), .A2(n114003), .B1(n120773), .B2(n120541), 
        .ZN(n7023) );
  OAI22_X1 U84683 ( .A1(n120546), .A2(n114002), .B1(n120776), .B2(n120541), 
        .ZN(n7024) );
  OAI22_X1 U84684 ( .A1(n120546), .A2(n114001), .B1(n120779), .B2(n120541), 
        .ZN(n7025) );
  OAI22_X1 U84685 ( .A1(n120546), .A2(n114000), .B1(n120782), .B2(n120541), 
        .ZN(n7026) );
  OAI22_X1 U84686 ( .A1(n120546), .A2(n113999), .B1(n120785), .B2(n120541), 
        .ZN(n7027) );
  OAI22_X1 U84687 ( .A1(n120545), .A2(n113998), .B1(n120788), .B2(n120541), 
        .ZN(n7028) );
  OAI22_X1 U84688 ( .A1(n120545), .A2(n113997), .B1(n120791), .B2(n120541), 
        .ZN(n7029) );
  OAI22_X1 U84689 ( .A1(n120545), .A2(n113996), .B1(n120794), .B2(n120541), 
        .ZN(n7030) );
  OAI22_X1 U84690 ( .A1(n120545), .A2(n113995), .B1(n120797), .B2(n120541), 
        .ZN(n7031) );
  OAI22_X1 U84691 ( .A1(n120545), .A2(n113994), .B1(n120800), .B2(n120541), 
        .ZN(n7032) );
  OAI22_X1 U84692 ( .A1(n120545), .A2(n113993), .B1(n120803), .B2(n120541), 
        .ZN(n7033) );
  OAI22_X1 U84693 ( .A1(n120545), .A2(n113992), .B1(n120806), .B2(n120541), 
        .ZN(n7034) );
  OAI22_X1 U84694 ( .A1(n120829), .A2(n113890), .B1(n120821), .B2(n120629), 
        .ZN(n7423) );
  OAI22_X1 U84695 ( .A1(n120833), .A2(n113888), .B1(n120821), .B2(n120632), 
        .ZN(n7424) );
  OAI22_X1 U84696 ( .A1(n120833), .A2(n113886), .B1(n120821), .B2(n120635), 
        .ZN(n7425) );
  OAI22_X1 U84697 ( .A1(n120833), .A2(n113884), .B1(n120821), .B2(n120638), 
        .ZN(n7426) );
  OAI22_X1 U84698 ( .A1(n120833), .A2(n113882), .B1(n120821), .B2(n120641), 
        .ZN(n7427) );
  OAI22_X1 U84699 ( .A1(n120833), .A2(n113880), .B1(n120821), .B2(n120644), 
        .ZN(n7428) );
  OAI22_X1 U84700 ( .A1(n120833), .A2(n113878), .B1(n120821), .B2(n120647), 
        .ZN(n7429) );
  OAI22_X1 U84701 ( .A1(n120833), .A2(n113876), .B1(n120821), .B2(n120650), 
        .ZN(n7430) );
  OAI22_X1 U84702 ( .A1(n120833), .A2(n113874), .B1(n120821), .B2(n120653), 
        .ZN(n7431) );
  OAI22_X1 U84703 ( .A1(n120833), .A2(n113872), .B1(n120821), .B2(n120656), 
        .ZN(n7432) );
  OAI22_X1 U84704 ( .A1(n120833), .A2(n113870), .B1(n120821), .B2(n120659), 
        .ZN(n7433) );
  OAI22_X1 U84705 ( .A1(n120833), .A2(n113868), .B1(n120821), .B2(n120662), 
        .ZN(n7434) );
  OAI22_X1 U84706 ( .A1(n120390), .A2(n114233), .B1(n120630), .B2(n120379), 
        .ZN(n6143) );
  OAI22_X1 U84707 ( .A1(n120390), .A2(n114232), .B1(n120633), .B2(n120379), 
        .ZN(n6144) );
  OAI22_X1 U84708 ( .A1(n120390), .A2(n114231), .B1(n120636), .B2(n120379), 
        .ZN(n6145) );
  OAI22_X1 U84709 ( .A1(n120390), .A2(n114230), .B1(n120639), .B2(n120379), 
        .ZN(n6146) );
  OAI22_X1 U84710 ( .A1(n120389), .A2(n114229), .B1(n120642), .B2(n120379), 
        .ZN(n6147) );
  OAI22_X1 U84711 ( .A1(n120389), .A2(n114228), .B1(n120645), .B2(n120379), 
        .ZN(n6148) );
  OAI22_X1 U84712 ( .A1(n120389), .A2(n114227), .B1(n120648), .B2(n120379), 
        .ZN(n6149) );
  OAI22_X1 U84713 ( .A1(n120389), .A2(n114226), .B1(n120651), .B2(n120379), 
        .ZN(n6150) );
  OAI22_X1 U84714 ( .A1(n120389), .A2(n114225), .B1(n120654), .B2(n120379), 
        .ZN(n6151) );
  OAI22_X1 U84715 ( .A1(n120389), .A2(n114224), .B1(n120657), .B2(n120379), 
        .ZN(n6152) );
  OAI22_X1 U84716 ( .A1(n120389), .A2(n114223), .B1(n120660), .B2(n120379), 
        .ZN(n6153) );
  OAI22_X1 U84717 ( .A1(n120389), .A2(n114222), .B1(n120663), .B2(n120379), 
        .ZN(n6154) );
  OAI22_X1 U84718 ( .A1(n120389), .A2(n114221), .B1(n120666), .B2(n120380), 
        .ZN(n6155) );
  OAI22_X1 U84719 ( .A1(n120389), .A2(n114220), .B1(n120669), .B2(n120380), 
        .ZN(n6156) );
  OAI22_X1 U84720 ( .A1(n120389), .A2(n114219), .B1(n120672), .B2(n120380), 
        .ZN(n6157) );
  OAI22_X1 U84721 ( .A1(n120389), .A2(n114218), .B1(n120675), .B2(n120380), 
        .ZN(n6158) );
  OAI22_X1 U84722 ( .A1(n120389), .A2(n114217), .B1(n120678), .B2(n120380), 
        .ZN(n6159) );
  OAI22_X1 U84723 ( .A1(n120388), .A2(n114216), .B1(n120681), .B2(n120380), 
        .ZN(n6160) );
  OAI22_X1 U84724 ( .A1(n120388), .A2(n114215), .B1(n120684), .B2(n120380), 
        .ZN(n6161) );
  OAI22_X1 U84725 ( .A1(n120570), .A2(n113979), .B1(n120629), .B2(n120562), 
        .ZN(n7103) );
  OAI22_X1 U84726 ( .A1(n120570), .A2(n113978), .B1(n120632), .B2(n120562), 
        .ZN(n7104) );
  OAI22_X1 U84727 ( .A1(n120570), .A2(n113977), .B1(n120635), .B2(n120562), 
        .ZN(n7105) );
  OAI22_X1 U84728 ( .A1(n120570), .A2(n113976), .B1(n120638), .B2(n120562), 
        .ZN(n7106) );
  OAI22_X1 U84729 ( .A1(n120570), .A2(n113975), .B1(n120641), .B2(n120562), 
        .ZN(n7107) );
  OAI22_X1 U84730 ( .A1(n120570), .A2(n113974), .B1(n120644), .B2(n120562), 
        .ZN(n7108) );
  OAI22_X1 U84731 ( .A1(n120570), .A2(n113973), .B1(n120647), .B2(n120562), 
        .ZN(n7109) );
  OAI22_X1 U84732 ( .A1(n120570), .A2(n113972), .B1(n120650), .B2(n120562), 
        .ZN(n7110) );
  OAI22_X1 U84733 ( .A1(n120570), .A2(n113971), .B1(n120653), .B2(n120562), 
        .ZN(n7111) );
  OAI22_X1 U84734 ( .A1(n120570), .A2(n113970), .B1(n120656), .B2(n120562), 
        .ZN(n7112) );
  OAI22_X1 U84735 ( .A1(n120570), .A2(n113969), .B1(n120659), .B2(n120562), 
        .ZN(n7113) );
  OAI22_X1 U84736 ( .A1(n120570), .A2(n113968), .B1(n120662), .B2(n120562), 
        .ZN(n7114) );
  OAI22_X1 U84737 ( .A1(n120571), .A2(n113967), .B1(n120665), .B2(n120563), 
        .ZN(n7115) );
  OAI22_X1 U84738 ( .A1(n120571), .A2(n113966), .B1(n120668), .B2(n120563), 
        .ZN(n7116) );
  OAI22_X1 U84739 ( .A1(n120571), .A2(n113965), .B1(n120671), .B2(n120563), 
        .ZN(n7117) );
  OAI22_X1 U84740 ( .A1(n120571), .A2(n113964), .B1(n120674), .B2(n120563), 
        .ZN(n7118) );
  OAI22_X1 U84741 ( .A1(n120571), .A2(n113963), .B1(n120677), .B2(n120563), 
        .ZN(n7119) );
  OAI22_X1 U84742 ( .A1(n120571), .A2(n113962), .B1(n120680), .B2(n120563), 
        .ZN(n7120) );
  OAI22_X1 U84743 ( .A1(n120571), .A2(n113961), .B1(n120683), .B2(n120563), 
        .ZN(n7121) );
  OAI22_X1 U84744 ( .A1(n120571), .A2(n113960), .B1(n120686), .B2(n120563), 
        .ZN(n7122) );
  OAI22_X1 U84745 ( .A1(n120571), .A2(n113959), .B1(n120689), .B2(n120563), 
        .ZN(n7123) );
  OAI22_X1 U84746 ( .A1(n120571), .A2(n113958), .B1(n120692), .B2(n120563), 
        .ZN(n7124) );
  OAI22_X1 U84747 ( .A1(n120571), .A2(n113957), .B1(n120695), .B2(n120563), 
        .ZN(n7125) );
  OAI22_X1 U84748 ( .A1(n120571), .A2(n113956), .B1(n120698), .B2(n120563), 
        .ZN(n7126) );
  OAI22_X1 U84749 ( .A1(n120571), .A2(n113955), .B1(n120701), .B2(n120564), 
        .ZN(n7127) );
  OAI22_X1 U84750 ( .A1(n120572), .A2(n113954), .B1(n120704), .B2(n120564), 
        .ZN(n7128) );
  OAI22_X1 U84751 ( .A1(n120572), .A2(n113953), .B1(n120707), .B2(n120564), 
        .ZN(n7129) );
  OAI22_X1 U84752 ( .A1(n120572), .A2(n113952), .B1(n120710), .B2(n120564), 
        .ZN(n7130) );
  OAI22_X1 U84753 ( .A1(n120572), .A2(n113951), .B1(n120713), .B2(n120564), 
        .ZN(n7131) );
  OAI22_X1 U84754 ( .A1(n120572), .A2(n113950), .B1(n120716), .B2(n120564), 
        .ZN(n7132) );
  OAI22_X1 U84755 ( .A1(n120572), .A2(n113949), .B1(n120719), .B2(n120564), 
        .ZN(n7133) );
  OAI22_X1 U84756 ( .A1(n120572), .A2(n113948), .B1(n120722), .B2(n120564), 
        .ZN(n7134) );
  OAI22_X1 U84757 ( .A1(n120572), .A2(n113947), .B1(n120725), .B2(n120564), 
        .ZN(n7135) );
  OAI22_X1 U84758 ( .A1(n120572), .A2(n113946), .B1(n120728), .B2(n120564), 
        .ZN(n7136) );
  OAI22_X1 U84759 ( .A1(n120572), .A2(n113945), .B1(n120731), .B2(n120564), 
        .ZN(n7137) );
  OAI22_X1 U84760 ( .A1(n120572), .A2(n113944), .B1(n120734), .B2(n120564), 
        .ZN(n7138) );
  OAI22_X1 U84761 ( .A1(n120572), .A2(n113943), .B1(n120737), .B2(n120565), 
        .ZN(n7139) );
  OAI22_X1 U84762 ( .A1(n120572), .A2(n113942), .B1(n120740), .B2(n120565), 
        .ZN(n7140) );
  OAI22_X1 U84763 ( .A1(n120573), .A2(n113941), .B1(n120743), .B2(n120565), 
        .ZN(n7141) );
  OAI22_X1 U84764 ( .A1(n120573), .A2(n113940), .B1(n120746), .B2(n120565), 
        .ZN(n7142) );
  OAI22_X1 U84765 ( .A1(n120573), .A2(n113939), .B1(n120749), .B2(n120565), 
        .ZN(n7143) );
  OAI22_X1 U84766 ( .A1(n120573), .A2(n113938), .B1(n120752), .B2(n120565), 
        .ZN(n7144) );
  OAI22_X1 U84767 ( .A1(n120573), .A2(n113937), .B1(n120755), .B2(n120565), 
        .ZN(n7145) );
  OAI22_X1 U84768 ( .A1(n120573), .A2(n113936), .B1(n120758), .B2(n120565), 
        .ZN(n7146) );
  OAI22_X1 U84769 ( .A1(n120573), .A2(n113935), .B1(n120761), .B2(n120565), 
        .ZN(n7147) );
  OAI22_X1 U84770 ( .A1(n120573), .A2(n113934), .B1(n120764), .B2(n120565), 
        .ZN(n7148) );
  OAI22_X1 U84771 ( .A1(n120573), .A2(n113933), .B1(n120767), .B2(n120565), 
        .ZN(n7149) );
  OAI22_X1 U84772 ( .A1(n120573), .A2(n113932), .B1(n120770), .B2(n120565), 
        .ZN(n7150) );
  OAI22_X1 U84773 ( .A1(n120573), .A2(n113931), .B1(n120773), .B2(n120566), 
        .ZN(n7151) );
  OAI22_X1 U84774 ( .A1(n120573), .A2(n113930), .B1(n120776), .B2(n120566), 
        .ZN(n7152) );
  OAI22_X1 U84775 ( .A1(n120573), .A2(n113929), .B1(n120779), .B2(n120566), 
        .ZN(n7153) );
  OAI22_X1 U84776 ( .A1(n120574), .A2(n113928), .B1(n120782), .B2(n120566), 
        .ZN(n7154) );
  OAI22_X1 U84777 ( .A1(n120574), .A2(n113927), .B1(n120785), .B2(n120566), 
        .ZN(n7155) );
  OAI22_X1 U84778 ( .A1(n120574), .A2(n113926), .B1(n120788), .B2(n120566), 
        .ZN(n7156) );
  OAI22_X1 U84779 ( .A1(n120574), .A2(n113925), .B1(n120791), .B2(n120566), 
        .ZN(n7157) );
  OAI22_X1 U84780 ( .A1(n120574), .A2(n113924), .B1(n120794), .B2(n120566), 
        .ZN(n7158) );
  OAI22_X1 U84781 ( .A1(n120574), .A2(n113923), .B1(n120797), .B2(n120566), 
        .ZN(n7159) );
  OAI22_X1 U84782 ( .A1(n120574), .A2(n113922), .B1(n120800), .B2(n120566), 
        .ZN(n7160) );
  OAI22_X1 U84783 ( .A1(n120574), .A2(n113921), .B1(n120803), .B2(n120566), 
        .ZN(n7161) );
  OAI22_X1 U84784 ( .A1(n120574), .A2(n113920), .B1(n120806), .B2(n120566), 
        .ZN(n7162) );
  OAI22_X1 U84785 ( .A1(n120374), .A2(n114299), .B1(n120630), .B2(n120366), 
        .ZN(n6079) );
  OAI22_X1 U84786 ( .A1(n120374), .A2(n114298), .B1(n120633), .B2(n120366), 
        .ZN(n6080) );
  OAI22_X1 U84787 ( .A1(n120374), .A2(n114297), .B1(n120636), .B2(n120366), 
        .ZN(n6081) );
  OAI22_X1 U84788 ( .A1(n120374), .A2(n114296), .B1(n120639), .B2(n120366), 
        .ZN(n6082) );
  OAI22_X1 U84789 ( .A1(n120374), .A2(n114295), .B1(n120642), .B2(n120366), 
        .ZN(n6083) );
  OAI22_X1 U84790 ( .A1(n120374), .A2(n114294), .B1(n120645), .B2(n120366), 
        .ZN(n6084) );
  OAI22_X1 U84791 ( .A1(n120374), .A2(n114293), .B1(n120648), .B2(n120366), 
        .ZN(n6085) );
  OAI22_X1 U84792 ( .A1(n120374), .A2(n114292), .B1(n120651), .B2(n120366), 
        .ZN(n6086) );
  OAI22_X1 U84793 ( .A1(n120374), .A2(n114291), .B1(n120654), .B2(n120366), 
        .ZN(n6087) );
  OAI22_X1 U84794 ( .A1(n120374), .A2(n114290), .B1(n120657), .B2(n120366), 
        .ZN(n6088) );
  OAI22_X1 U84795 ( .A1(n120374), .A2(n114289), .B1(n120660), .B2(n120366), 
        .ZN(n6089) );
  OAI22_X1 U84796 ( .A1(n120374), .A2(n114288), .B1(n120663), .B2(n120366), 
        .ZN(n6090) );
  OAI22_X1 U84797 ( .A1(n120375), .A2(n114287), .B1(n120666), .B2(n120367), 
        .ZN(n6091) );
  OAI22_X1 U84798 ( .A1(n120375), .A2(n114286), .B1(n120669), .B2(n120367), 
        .ZN(n6092) );
  OAI22_X1 U84799 ( .A1(n120375), .A2(n114285), .B1(n120672), .B2(n120367), 
        .ZN(n6093) );
  OAI22_X1 U84800 ( .A1(n120375), .A2(n114284), .B1(n120675), .B2(n120367), 
        .ZN(n6094) );
  OAI22_X1 U84801 ( .A1(n120375), .A2(n114283), .B1(n120678), .B2(n120367), 
        .ZN(n6095) );
  OAI22_X1 U84802 ( .A1(n120375), .A2(n114282), .B1(n120681), .B2(n120367), 
        .ZN(n6096) );
  OAI22_X1 U84803 ( .A1(n120375), .A2(n114281), .B1(n120684), .B2(n120367), 
        .ZN(n6097) );
  OAI22_X1 U84804 ( .A1(n120375), .A2(n114280), .B1(n120687), .B2(n120367), 
        .ZN(n6098) );
  OAI22_X1 U84805 ( .A1(n120375), .A2(n114279), .B1(n120690), .B2(n120367), 
        .ZN(n6099) );
  OAI22_X1 U84806 ( .A1(n120375), .A2(n114278), .B1(n120693), .B2(n120367), 
        .ZN(n6100) );
  OAI22_X1 U84807 ( .A1(n120375), .A2(n114277), .B1(n120696), .B2(n120367), 
        .ZN(n6101) );
  OAI22_X1 U84808 ( .A1(n120375), .A2(n114276), .B1(n120699), .B2(n120367), 
        .ZN(n6102) );
  OAI22_X1 U84809 ( .A1(n120375), .A2(n114275), .B1(n120702), .B2(n120368), 
        .ZN(n6103) );
  OAI22_X1 U84810 ( .A1(n120376), .A2(n114274), .B1(n120705), .B2(n120368), 
        .ZN(n6104) );
  OAI22_X1 U84811 ( .A1(n120376), .A2(n114273), .B1(n120708), .B2(n120368), 
        .ZN(n6105) );
  OAI22_X1 U84812 ( .A1(n120376), .A2(n114272), .B1(n120711), .B2(n120368), 
        .ZN(n6106) );
  OAI22_X1 U84813 ( .A1(n120376), .A2(n114271), .B1(n120714), .B2(n120368), 
        .ZN(n6107) );
  OAI22_X1 U84814 ( .A1(n120376), .A2(n114270), .B1(n120717), .B2(n120368), 
        .ZN(n6108) );
  OAI22_X1 U84815 ( .A1(n120376), .A2(n114269), .B1(n120720), .B2(n120368), 
        .ZN(n6109) );
  OAI22_X1 U84816 ( .A1(n120376), .A2(n114268), .B1(n120723), .B2(n120368), 
        .ZN(n6110) );
  OAI22_X1 U84817 ( .A1(n120376), .A2(n114267), .B1(n120726), .B2(n120368), 
        .ZN(n6111) );
  OAI22_X1 U84818 ( .A1(n120376), .A2(n114266), .B1(n120729), .B2(n120368), 
        .ZN(n6112) );
  OAI22_X1 U84819 ( .A1(n120376), .A2(n114265), .B1(n120732), .B2(n120368), 
        .ZN(n6113) );
  OAI22_X1 U84820 ( .A1(n120376), .A2(n114264), .B1(n120735), .B2(n120368), 
        .ZN(n6114) );
  OAI22_X1 U84821 ( .A1(n120376), .A2(n114263), .B1(n120738), .B2(n120369), 
        .ZN(n6115) );
  OAI22_X1 U84822 ( .A1(n120376), .A2(n114262), .B1(n120741), .B2(n120369), 
        .ZN(n6116) );
  OAI22_X1 U84823 ( .A1(n120377), .A2(n114261), .B1(n120744), .B2(n120369), 
        .ZN(n6117) );
  OAI22_X1 U84824 ( .A1(n120377), .A2(n114260), .B1(n120747), .B2(n120369), 
        .ZN(n6118) );
  OAI22_X1 U84825 ( .A1(n120377), .A2(n114259), .B1(n120750), .B2(n120369), 
        .ZN(n6119) );
  OAI22_X1 U84826 ( .A1(n120377), .A2(n114258), .B1(n120753), .B2(n120369), 
        .ZN(n6120) );
  OAI22_X1 U84827 ( .A1(n120377), .A2(n114257), .B1(n120756), .B2(n120369), 
        .ZN(n6121) );
  OAI22_X1 U84828 ( .A1(n120377), .A2(n114256), .B1(n120759), .B2(n120369), 
        .ZN(n6122) );
  OAI22_X1 U84829 ( .A1(n120377), .A2(n114255), .B1(n120762), .B2(n120369), 
        .ZN(n6123) );
  OAI22_X1 U84830 ( .A1(n120377), .A2(n114254), .B1(n120765), .B2(n120369), 
        .ZN(n6124) );
  OAI22_X1 U84831 ( .A1(n120377), .A2(n114253), .B1(n120768), .B2(n120369), 
        .ZN(n6125) );
  OAI22_X1 U84832 ( .A1(n120377), .A2(n114252), .B1(n120771), .B2(n120369), 
        .ZN(n6126) );
  OAI22_X1 U84833 ( .A1(n120377), .A2(n114251), .B1(n120774), .B2(n120370), 
        .ZN(n6127) );
  OAI22_X1 U84834 ( .A1(n120377), .A2(n114250), .B1(n120777), .B2(n120370), 
        .ZN(n6128) );
  OAI22_X1 U84835 ( .A1(n120377), .A2(n114249), .B1(n120780), .B2(n120370), 
        .ZN(n6129) );
  OAI22_X1 U84836 ( .A1(n120378), .A2(n114248), .B1(n120783), .B2(n120370), 
        .ZN(n6130) );
  OAI22_X1 U84837 ( .A1(n120378), .A2(n114247), .B1(n120786), .B2(n120370), 
        .ZN(n6131) );
  OAI22_X1 U84838 ( .A1(n120378), .A2(n114246), .B1(n120789), .B2(n120370), 
        .ZN(n6132) );
  OAI22_X1 U84839 ( .A1(n120378), .A2(n114245), .B1(n120792), .B2(n120370), 
        .ZN(n6133) );
  OAI22_X1 U84840 ( .A1(n120378), .A2(n114244), .B1(n120795), .B2(n120370), 
        .ZN(n6134) );
  OAI22_X1 U84841 ( .A1(n120378), .A2(n114243), .B1(n120798), .B2(n120370), 
        .ZN(n6135) );
  OAI22_X1 U84842 ( .A1(n120378), .A2(n114242), .B1(n120801), .B2(n120370), 
        .ZN(n6136) );
  OAI22_X1 U84843 ( .A1(n120378), .A2(n114241), .B1(n120804), .B2(n120370), 
        .ZN(n6137) );
  OAI22_X1 U84844 ( .A1(n120378), .A2(n114240), .B1(n120807), .B2(n120370), 
        .ZN(n6138) );
  OAI22_X1 U84845 ( .A1(n120411), .A2(n114210), .B1(n120630), .B2(n120403), 
        .ZN(n6271) );
  OAI22_X1 U84846 ( .A1(n120411), .A2(n114209), .B1(n120633), .B2(n120403), 
        .ZN(n6272) );
  OAI22_X1 U84847 ( .A1(n120411), .A2(n114208), .B1(n120636), .B2(n120403), 
        .ZN(n6273) );
  OAI22_X1 U84848 ( .A1(n120411), .A2(n114207), .B1(n120639), .B2(n120403), 
        .ZN(n6274) );
  OAI22_X1 U84849 ( .A1(n120411), .A2(n114206), .B1(n120642), .B2(n120403), 
        .ZN(n6275) );
  OAI22_X1 U84850 ( .A1(n120411), .A2(n114205), .B1(n120645), .B2(n120403), 
        .ZN(n6276) );
  OAI22_X1 U84851 ( .A1(n120411), .A2(n114204), .B1(n120648), .B2(n120403), 
        .ZN(n6277) );
  OAI22_X1 U84852 ( .A1(n120411), .A2(n114203), .B1(n120651), .B2(n120403), 
        .ZN(n6278) );
  OAI22_X1 U84853 ( .A1(n120411), .A2(n114202), .B1(n120654), .B2(n120403), 
        .ZN(n6279) );
  OAI22_X1 U84854 ( .A1(n120411), .A2(n114201), .B1(n120657), .B2(n120403), 
        .ZN(n6280) );
  OAI22_X1 U84855 ( .A1(n120411), .A2(n114200), .B1(n120660), .B2(n120403), 
        .ZN(n6281) );
  OAI22_X1 U84856 ( .A1(n120411), .A2(n114199), .B1(n120663), .B2(n120403), 
        .ZN(n6282) );
  OAI22_X1 U84857 ( .A1(n120412), .A2(n114198), .B1(n120666), .B2(n120404), 
        .ZN(n6283) );
  OAI22_X1 U84858 ( .A1(n120412), .A2(n114197), .B1(n120669), .B2(n120404), 
        .ZN(n6284) );
  OAI22_X1 U84859 ( .A1(n120412), .A2(n114196), .B1(n120672), .B2(n120404), 
        .ZN(n6285) );
  OAI22_X1 U84860 ( .A1(n120412), .A2(n114195), .B1(n120675), .B2(n120404), 
        .ZN(n6286) );
  OAI22_X1 U84861 ( .A1(n120412), .A2(n114194), .B1(n120678), .B2(n120404), 
        .ZN(n6287) );
  OAI22_X1 U84862 ( .A1(n120412), .A2(n114193), .B1(n120681), .B2(n120404), 
        .ZN(n6288) );
  OAI22_X1 U84863 ( .A1(n120412), .A2(n114192), .B1(n120684), .B2(n120404), 
        .ZN(n6289) );
  OAI22_X1 U84864 ( .A1(n120412), .A2(n114191), .B1(n120687), .B2(n120404), 
        .ZN(n6290) );
  OAI22_X1 U84865 ( .A1(n120412), .A2(n114190), .B1(n120690), .B2(n120404), 
        .ZN(n6291) );
  OAI22_X1 U84866 ( .A1(n120412), .A2(n114189), .B1(n120693), .B2(n120404), 
        .ZN(n6292) );
  OAI22_X1 U84867 ( .A1(n120412), .A2(n114188), .B1(n120696), .B2(n120404), 
        .ZN(n6293) );
  OAI22_X1 U84868 ( .A1(n120412), .A2(n114187), .B1(n120699), .B2(n120404), 
        .ZN(n6294) );
  OAI22_X1 U84869 ( .A1(n120412), .A2(n114186), .B1(n120702), .B2(n120405), 
        .ZN(n6295) );
  OAI22_X1 U84870 ( .A1(n120413), .A2(n114185), .B1(n120705), .B2(n120405), 
        .ZN(n6296) );
  OAI22_X1 U84871 ( .A1(n120413), .A2(n114184), .B1(n120708), .B2(n120405), 
        .ZN(n6297) );
  OAI22_X1 U84872 ( .A1(n120413), .A2(n114183), .B1(n120711), .B2(n120405), 
        .ZN(n6298) );
  OAI22_X1 U84873 ( .A1(n120413), .A2(n114182), .B1(n120714), .B2(n120405), 
        .ZN(n6299) );
  OAI22_X1 U84874 ( .A1(n120413), .A2(n114181), .B1(n120717), .B2(n120405), 
        .ZN(n6300) );
  OAI22_X1 U84875 ( .A1(n120413), .A2(n114180), .B1(n120720), .B2(n120405), 
        .ZN(n6301) );
  OAI22_X1 U84876 ( .A1(n120413), .A2(n114179), .B1(n120723), .B2(n120405), 
        .ZN(n6302) );
  OAI22_X1 U84877 ( .A1(n120413), .A2(n114178), .B1(n120726), .B2(n120405), 
        .ZN(n6303) );
  OAI22_X1 U84878 ( .A1(n120413), .A2(n114177), .B1(n120729), .B2(n120405), 
        .ZN(n6304) );
  OAI22_X1 U84879 ( .A1(n120413), .A2(n114176), .B1(n120732), .B2(n120405), 
        .ZN(n6305) );
  OAI22_X1 U84880 ( .A1(n120413), .A2(n114175), .B1(n120735), .B2(n120405), 
        .ZN(n6306) );
  OAI22_X1 U84881 ( .A1(n120413), .A2(n114174), .B1(n120738), .B2(n120406), 
        .ZN(n6307) );
  OAI22_X1 U84882 ( .A1(n120413), .A2(n114173), .B1(n120741), .B2(n120406), 
        .ZN(n6308) );
  OAI22_X1 U84883 ( .A1(n120414), .A2(n114172), .B1(n120744), .B2(n120406), 
        .ZN(n6309) );
  OAI22_X1 U84884 ( .A1(n120414), .A2(n114171), .B1(n120747), .B2(n120406), 
        .ZN(n6310) );
  OAI22_X1 U84885 ( .A1(n120414), .A2(n114170), .B1(n120750), .B2(n120406), 
        .ZN(n6311) );
  OAI22_X1 U84886 ( .A1(n120414), .A2(n114169), .B1(n120753), .B2(n120406), 
        .ZN(n6312) );
  OAI22_X1 U84887 ( .A1(n120414), .A2(n114168), .B1(n120756), .B2(n120406), 
        .ZN(n6313) );
  OAI22_X1 U84888 ( .A1(n120414), .A2(n114167), .B1(n120759), .B2(n120406), 
        .ZN(n6314) );
  OAI22_X1 U84889 ( .A1(n120414), .A2(n114166), .B1(n120762), .B2(n120406), 
        .ZN(n6315) );
  OAI22_X1 U84890 ( .A1(n120414), .A2(n114165), .B1(n120765), .B2(n120406), 
        .ZN(n6316) );
  OAI22_X1 U84891 ( .A1(n120414), .A2(n114164), .B1(n120768), .B2(n120406), 
        .ZN(n6317) );
  OAI22_X1 U84892 ( .A1(n120414), .A2(n114163), .B1(n120771), .B2(n120406), 
        .ZN(n6318) );
  OAI22_X1 U84893 ( .A1(n120414), .A2(n114162), .B1(n120774), .B2(n120407), 
        .ZN(n6319) );
  OAI22_X1 U84894 ( .A1(n120414), .A2(n114161), .B1(n120777), .B2(n120407), 
        .ZN(n6320) );
  OAI22_X1 U84895 ( .A1(n120414), .A2(n114160), .B1(n120780), .B2(n120407), 
        .ZN(n6321) );
  OAI22_X1 U84896 ( .A1(n120415), .A2(n114159), .B1(n120783), .B2(n120407), 
        .ZN(n6322) );
  OAI22_X1 U84897 ( .A1(n120415), .A2(n114158), .B1(n120786), .B2(n120407), 
        .ZN(n6323) );
  OAI22_X1 U84898 ( .A1(n120415), .A2(n114157), .B1(n120789), .B2(n120407), 
        .ZN(n6324) );
  OAI22_X1 U84899 ( .A1(n120415), .A2(n114156), .B1(n120792), .B2(n120407), 
        .ZN(n6325) );
  OAI22_X1 U84900 ( .A1(n120415), .A2(n114155), .B1(n120795), .B2(n120407), 
        .ZN(n6326) );
  OAI22_X1 U84901 ( .A1(n120415), .A2(n114154), .B1(n120798), .B2(n120407), 
        .ZN(n6327) );
  OAI22_X1 U84902 ( .A1(n120415), .A2(n114153), .B1(n120801), .B2(n120407), 
        .ZN(n6328) );
  OAI22_X1 U84903 ( .A1(n120415), .A2(n114152), .B1(n120804), .B2(n120407), 
        .ZN(n6329) );
  OAI22_X1 U84904 ( .A1(n120415), .A2(n114151), .B1(n120807), .B2(n120407), 
        .ZN(n6330) );
  OAI21_X1 U84905 ( .B1(n113901), .B2(n113913), .A(n120623), .ZN(n113914) );
  OAI21_X1 U84906 ( .B1(n113901), .B2(n113986), .A(n120623), .ZN(n113990) );
  BUF_X1 U84907 ( .A(n113891), .Z(n120631) );
  BUF_X1 U84908 ( .A(n113889), .Z(n120634) );
  BUF_X1 U84909 ( .A(n113887), .Z(n120637) );
  BUF_X1 U84910 ( .A(n113885), .Z(n120640) );
  BUF_X1 U84911 ( .A(n113883), .Z(n120643) );
  BUF_X1 U84912 ( .A(n113881), .Z(n120646) );
  BUF_X1 U84913 ( .A(n113879), .Z(n120649) );
  BUF_X1 U84914 ( .A(n113877), .Z(n120652) );
  BUF_X1 U84915 ( .A(n113875), .Z(n120655) );
  BUF_X1 U84916 ( .A(n113873), .Z(n120658) );
  BUF_X1 U84917 ( .A(n113871), .Z(n120661) );
  BUF_X1 U84918 ( .A(n113869), .Z(n120664) );
  BUF_X1 U84919 ( .A(n113867), .Z(n120667) );
  BUF_X1 U84920 ( .A(n113865), .Z(n120670) );
  BUF_X1 U84921 ( .A(n113863), .Z(n120673) );
  BUF_X1 U84922 ( .A(n113861), .Z(n120676) );
  BUF_X1 U84923 ( .A(n113859), .Z(n120679) );
  BUF_X1 U84924 ( .A(n113857), .Z(n120682) );
  BUF_X1 U84925 ( .A(n113855), .Z(n120685) );
  BUF_X1 U84926 ( .A(n113853), .Z(n120688) );
  BUF_X1 U84927 ( .A(n113851), .Z(n120691) );
  BUF_X1 U84928 ( .A(n113849), .Z(n120694) );
  BUF_X1 U84929 ( .A(n113847), .Z(n120697) );
  BUF_X1 U84930 ( .A(n113845), .Z(n120700) );
  BUF_X1 U84931 ( .A(n113843), .Z(n120703) );
  BUF_X1 U84932 ( .A(n113841), .Z(n120706) );
  BUF_X1 U84933 ( .A(n113839), .Z(n120709) );
  BUF_X1 U84934 ( .A(n113837), .Z(n120712) );
  BUF_X1 U84935 ( .A(n113835), .Z(n120715) );
  BUF_X1 U84936 ( .A(n113833), .Z(n120718) );
  BUF_X1 U84937 ( .A(n113831), .Z(n120721) );
  BUF_X1 U84938 ( .A(n113829), .Z(n120724) );
  BUF_X1 U84939 ( .A(n113827), .Z(n120727) );
  BUF_X1 U84940 ( .A(n113825), .Z(n120730) );
  BUF_X1 U84941 ( .A(n113823), .Z(n120733) );
  BUF_X1 U84942 ( .A(n113821), .Z(n120736) );
  BUF_X1 U84943 ( .A(n113819), .Z(n120739) );
  BUF_X1 U84944 ( .A(n113817), .Z(n120742) );
  BUF_X1 U84945 ( .A(n113815), .Z(n120745) );
  BUF_X1 U84946 ( .A(n113813), .Z(n120748) );
  BUF_X1 U84947 ( .A(n113811), .Z(n120751) );
  BUF_X1 U84948 ( .A(n113809), .Z(n120754) );
  BUF_X1 U84949 ( .A(n113807), .Z(n120757) );
  BUF_X1 U84950 ( .A(n113805), .Z(n120760) );
  BUF_X1 U84951 ( .A(n113803), .Z(n120763) );
  BUF_X1 U84952 ( .A(n113801), .Z(n120766) );
  BUF_X1 U84953 ( .A(n113799), .Z(n120769) );
  BUF_X1 U84954 ( .A(n113797), .Z(n120772) );
  BUF_X1 U84955 ( .A(n113795), .Z(n120775) );
  BUF_X1 U84956 ( .A(n113793), .Z(n120778) );
  BUF_X1 U84957 ( .A(n113791), .Z(n120781) );
  BUF_X1 U84958 ( .A(n113789), .Z(n120784) );
  BUF_X1 U84959 ( .A(n113787), .Z(n120787) );
  BUF_X1 U84960 ( .A(n113785), .Z(n120790) );
  BUF_X1 U84961 ( .A(n113783), .Z(n120793) );
  BUF_X1 U84962 ( .A(n113781), .Z(n120796) );
  BUF_X1 U84963 ( .A(n113779), .Z(n120799) );
  BUF_X1 U84964 ( .A(n113777), .Z(n120802) );
  BUF_X1 U84965 ( .A(n113775), .Z(n120805) );
  BUF_X1 U84966 ( .A(n113771), .Z(n120811) );
  BUF_X1 U84967 ( .A(n113770), .Z(n120814) );
  BUF_X1 U84968 ( .A(n113769), .Z(n120817) );
  BUF_X1 U84969 ( .A(n113768), .Z(n120820) );
  BUF_X1 U84970 ( .A(n113773), .Z(n120808) );
  OAI21_X1 U84971 ( .B1(n113986), .B2(n114374), .A(n120624), .ZN(n114643) );
  OAI21_X1 U84972 ( .B1(n113908), .B2(n114141), .A(n120624), .ZN(n114145) );
  OAI21_X1 U84973 ( .B1(n113908), .B2(n114374), .A(n120625), .ZN(n114443) );
  OAI21_X1 U84974 ( .B1(n113894), .B2(n114121), .A(n120623), .ZN(n114055) );
  OAI21_X1 U84975 ( .B1(n113913), .B2(n114144), .A(n120624), .ZN(n114234) );
  OAI21_X1 U84976 ( .B1(n113894), .B2(n114371), .A(n120625), .ZN(n114305) );
  OAI21_X1 U84977 ( .B1(n113913), .B2(n114371), .A(n120625), .ZN(n114509) );
  OAI21_X1 U84978 ( .B1(n113986), .B2(n114371), .A(n120625), .ZN(n114577) );
  OAI21_X1 U84979 ( .B1(n113908), .B2(n114371), .A(n120625), .ZN(n114377) );
  AND2_X1 U84980 ( .A1(n116453), .A2(n116454), .ZN(n114662) );
  AND2_X1 U84981 ( .A1(n117945), .A2(n117946), .ZN(n116490) );
  AND2_X1 U84982 ( .A1(n117953), .A2(n117959), .ZN(n116523) );
  AND2_X1 U84983 ( .A1(n116445), .A2(n116446), .ZN(n114657) );
  AND2_X1 U84984 ( .A1(n116445), .A2(n116463), .ZN(n114676) );
  AND2_X1 U84985 ( .A1(n116452), .A2(n116457), .ZN(n114670) );
  AND2_X1 U84986 ( .A1(n117955), .A2(n117948), .ZN(n116503) );
  AND2_X1 U84987 ( .A1(n117947), .A2(n117945), .ZN(n116502) );
  AND2_X1 U84988 ( .A1(n117947), .A2(n117953), .ZN(n116497) );
  AND2_X1 U84989 ( .A1(n117962), .A2(n117953), .ZN(n116507) );
  AND2_X1 U84990 ( .A1(n117947), .A2(n117954), .ZN(n116495) );
  AND2_X1 U84991 ( .A1(n117961), .A2(n117954), .ZN(n116508) );
  AND2_X1 U84992 ( .A1(n116452), .A2(n116447), .ZN(n114664) );
  AND2_X1 U84993 ( .A1(n116464), .A2(n116447), .ZN(n114675) );
  AND2_X1 U84994 ( .A1(n117955), .A2(n117954), .ZN(n116529) );
  AND2_X1 U84995 ( .A1(n117968), .A2(n117954), .ZN(n116522) );
  AND2_X1 U84996 ( .A1(n116454), .A2(n116447), .ZN(n114691) );
  AND2_X1 U84997 ( .A1(n116459), .A2(n116447), .ZN(n114698) );
  AND2_X1 U84998 ( .A1(n116452), .A2(n116445), .ZN(n114669) );
  AND2_X1 U84999 ( .A1(n116454), .A2(n116445), .ZN(n114693) );
  AND2_X1 U85000 ( .A1(n116458), .A2(n116445), .ZN(n114700) );
  NOR3_X1 U85001 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n116471), .ZN(n116448) );
  NOR3_X1 U85002 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n117970), .ZN(n117959) );
  NOR3_X1 U85003 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n117967), .ZN(n117968) );
  NOR3_X1 U85004 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n116470), .ZN(n116459) );
  NOR3_X1 U85005 ( .A1(n117967), .A2(ADD_RD2[4]), .A3(n117958), .ZN(n117961)
         );
  NOR3_X1 U85006 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n116469), .ZN(n116446) );
  NOR3_X1 U85007 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(
        n116464) );
  NOR3_X1 U85008 ( .A1(n117970), .A2(ADD_RD2[3]), .A3(n117967), .ZN(n117962)
         );
  NOR3_X1 U85009 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(
        n117946) );
  NOR3_X1 U85010 ( .A1(n116470), .A2(ADD_RD1[0]), .A3(n116471), .ZN(n116458)
         );
  NOR3_X1 U85011 ( .A1(n117970), .A2(ADD_RD2[0]), .A3(n117958), .ZN(n117955)
         );
  NOR3_X1 U85012 ( .A1(n116469), .A2(ADD_RD1[3]), .A3(n116471), .ZN(n116454)
         );
  NOR3_X1 U85013 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n117958), .ZN(n117947) );
  NOR3_X1 U85014 ( .A1(n116469), .A2(ADD_RD1[4]), .A3(n116470), .ZN(n116452)
         );
  OAI222_X1 U85015 ( .A1(n113968), .A2(n119904), .B1(n90359), .B2(n119898), 
        .C1(n99364), .C2(n119892), .ZN(n117709) );
  OAI222_X1 U85016 ( .A1(n113967), .A2(n119905), .B1(n90358), .B2(n119899), 
        .C1(n99363), .C2(n119893), .ZN(n117687) );
  OAI222_X1 U85017 ( .A1(n113966), .A2(n119905), .B1(n90357), .B2(n119899), 
        .C1(n99362), .C2(n119893), .ZN(n117665) );
  OAI222_X1 U85018 ( .A1(n113965), .A2(n119905), .B1(n90356), .B2(n119899), 
        .C1(n99361), .C2(n119893), .ZN(n117643) );
  OAI222_X1 U85019 ( .A1(n113964), .A2(n119905), .B1(n90355), .B2(n119899), 
        .C1(n99360), .C2(n119893), .ZN(n117621) );
  OAI222_X1 U85020 ( .A1(n113963), .A2(n119905), .B1(n90354), .B2(n119899), 
        .C1(n99359), .C2(n119893), .ZN(n117599) );
  OAI222_X1 U85021 ( .A1(n113962), .A2(n119905), .B1(n90353), .B2(n119899), 
        .C1(n99358), .C2(n119893), .ZN(n117577) );
  OAI222_X1 U85022 ( .A1(n113961), .A2(n119905), .B1(n90352), .B2(n119899), 
        .C1(n99357), .C2(n119893), .ZN(n117555) );
  OAI222_X1 U85023 ( .A1(n113960), .A2(n119905), .B1(n90351), .B2(n119899), 
        .C1(n99356), .C2(n119893), .ZN(n117532) );
  OAI222_X1 U85024 ( .A1(n113959), .A2(n119905), .B1(n90350), .B2(n119899), 
        .C1(n99355), .C2(n119893), .ZN(n117509) );
  OAI222_X1 U85025 ( .A1(n113958), .A2(n119905), .B1(n90349), .B2(n119899), 
        .C1(n99354), .C2(n119893), .ZN(n117486) );
  OAI222_X1 U85026 ( .A1(n113957), .A2(n119905), .B1(n90348), .B2(n119899), 
        .C1(n99353), .C2(n119893), .ZN(n117463) );
  OAI222_X1 U85027 ( .A1(n113956), .A2(n119905), .B1(n90347), .B2(n119899), 
        .C1(n99352), .C2(n119893), .ZN(n117440) );
  OAI222_X1 U85028 ( .A1(n113955), .A2(n119906), .B1(n90346), .B2(n119900), 
        .C1(n99351), .C2(n119894), .ZN(n117417) );
  OAI222_X1 U85029 ( .A1(n113954), .A2(n119906), .B1(n90345), .B2(n119900), 
        .C1(n99350), .C2(n119894), .ZN(n117394) );
  OAI222_X1 U85030 ( .A1(n113953), .A2(n119906), .B1(n90344), .B2(n119900), 
        .C1(n99349), .C2(n119894), .ZN(n117371) );
  OAI222_X1 U85031 ( .A1(n113952), .A2(n119906), .B1(n90343), .B2(n119900), 
        .C1(n99348), .C2(n119894), .ZN(n117348) );
  OAI222_X1 U85032 ( .A1(n113951), .A2(n119906), .B1(n90342), .B2(n119900), 
        .C1(n99347), .C2(n119894), .ZN(n117325) );
  OAI222_X1 U85033 ( .A1(n113950), .A2(n119906), .B1(n90341), .B2(n119900), 
        .C1(n99346), .C2(n119894), .ZN(n117302) );
  OAI222_X1 U85034 ( .A1(n113949), .A2(n119906), .B1(n90340), .B2(n119900), 
        .C1(n99345), .C2(n119894), .ZN(n117279) );
  OAI222_X1 U85035 ( .A1(n113948), .A2(n119906), .B1(n90339), .B2(n119900), 
        .C1(n99344), .C2(n119894), .ZN(n117256) );
  OAI222_X1 U85036 ( .A1(n113947), .A2(n119906), .B1(n90338), .B2(n119900), 
        .C1(n99343), .C2(n119894), .ZN(n117233) );
  OAI222_X1 U85037 ( .A1(n113946), .A2(n119906), .B1(n90337), .B2(n119900), 
        .C1(n99342), .C2(n119894), .ZN(n117210) );
  OAI222_X1 U85038 ( .A1(n113945), .A2(n119906), .B1(n90336), .B2(n119900), 
        .C1(n99341), .C2(n119894), .ZN(n117187) );
  OAI222_X1 U85039 ( .A1(n113944), .A2(n119906), .B1(n90335), .B2(n119900), 
        .C1(n99340), .C2(n119894), .ZN(n117164) );
  OAI222_X1 U85040 ( .A1(n113943), .A2(n119907), .B1(n90334), .B2(n119901), 
        .C1(n99339), .C2(n119895), .ZN(n117141) );
  OAI222_X1 U85041 ( .A1(n113942), .A2(n119907), .B1(n90333), .B2(n119901), 
        .C1(n99338), .C2(n119895), .ZN(n117118) );
  OAI222_X1 U85042 ( .A1(n113941), .A2(n119907), .B1(n90332), .B2(n119901), 
        .C1(n99337), .C2(n119895), .ZN(n117095) );
  OAI222_X1 U85043 ( .A1(n113940), .A2(n119907), .B1(n90331), .B2(n119901), 
        .C1(n99336), .C2(n119895), .ZN(n117072) );
  OAI222_X1 U85044 ( .A1(n113939), .A2(n119907), .B1(n90330), .B2(n119901), 
        .C1(n99335), .C2(n119895), .ZN(n117049) );
  OAI222_X1 U85045 ( .A1(n113938), .A2(n119907), .B1(n90329), .B2(n119901), 
        .C1(n99334), .C2(n119895), .ZN(n117026) );
  OAI222_X1 U85046 ( .A1(n113937), .A2(n119907), .B1(n90328), .B2(n119901), 
        .C1(n99333), .C2(n119895), .ZN(n117003) );
  OAI222_X1 U85047 ( .A1(n113936), .A2(n119907), .B1(n90327), .B2(n119901), 
        .C1(n99332), .C2(n119895), .ZN(n116980) );
  OAI222_X1 U85048 ( .A1(n113935), .A2(n119907), .B1(n90326), .B2(n119901), 
        .C1(n99331), .C2(n119895), .ZN(n116957) );
  OAI222_X1 U85049 ( .A1(n113934), .A2(n119907), .B1(n90325), .B2(n119901), 
        .C1(n99330), .C2(n119895), .ZN(n116934) );
  OAI222_X1 U85050 ( .A1(n113933), .A2(n119907), .B1(n90324), .B2(n119901), 
        .C1(n99329), .C2(n119895), .ZN(n116911) );
  OAI222_X1 U85051 ( .A1(n113932), .A2(n119907), .B1(n90323), .B2(n119901), 
        .C1(n99328), .C2(n119895), .ZN(n116888) );
  OAI222_X1 U85052 ( .A1(n113931), .A2(n119908), .B1(n90322), .B2(n119902), 
        .C1(n99327), .C2(n119896), .ZN(n116865) );
  OAI222_X1 U85053 ( .A1(n113930), .A2(n119908), .B1(n90321), .B2(n119902), 
        .C1(n99326), .C2(n119896), .ZN(n116842) );
  OAI222_X1 U85054 ( .A1(n113929), .A2(n119908), .B1(n90320), .B2(n119902), 
        .C1(n99325), .C2(n119896), .ZN(n116819) );
  OAI222_X1 U85055 ( .A1(n113928), .A2(n119908), .B1(n90319), .B2(n119902), 
        .C1(n99324), .C2(n119896), .ZN(n116796) );
  OAI222_X1 U85056 ( .A1(n113927), .A2(n119908), .B1(n90318), .B2(n119902), 
        .C1(n99323), .C2(n119896), .ZN(n116773) );
  OAI222_X1 U85057 ( .A1(n113926), .A2(n119908), .B1(n90317), .B2(n119902), 
        .C1(n99322), .C2(n119896), .ZN(n116750) );
  OAI222_X1 U85058 ( .A1(n113925), .A2(n119908), .B1(n90316), .B2(n119902), 
        .C1(n99321), .C2(n119896), .ZN(n116727) );
  OAI222_X1 U85059 ( .A1(n113924), .A2(n119908), .B1(n90315), .B2(n119902), 
        .C1(n99320), .C2(n119896), .ZN(n116704) );
  OAI222_X1 U85060 ( .A1(n113923), .A2(n119908), .B1(n90314), .B2(n119902), 
        .C1(n99319), .C2(n119896), .ZN(n116681) );
  OAI222_X1 U85061 ( .A1(n113922), .A2(n119908), .B1(n90313), .B2(n119902), 
        .C1(n99318), .C2(n119896), .ZN(n116658) );
  OAI222_X1 U85062 ( .A1(n113921), .A2(n119908), .B1(n90312), .B2(n119902), 
        .C1(n99317), .C2(n119896), .ZN(n116635) );
  OAI222_X1 U85063 ( .A1(n113920), .A2(n119908), .B1(n90311), .B2(n119902), 
        .C1(n99316), .C2(n119896), .ZN(n116612) );
  OAI222_X1 U85064 ( .A1(n99131), .A2(n120105), .B1(n120099), .B2(n115146), 
        .C1(n113933), .C2(n120093), .ZN(n115165) );
  OAI222_X1 U85065 ( .A1(n99130), .A2(n120105), .B1(n120099), .B2(n115118), 
        .C1(n113932), .C2(n120093), .ZN(n115137) );
  OAI222_X1 U85066 ( .A1(n99129), .A2(n120106), .B1(n120100), .B2(n115090), 
        .C1(n113931), .C2(n120094), .ZN(n115109) );
  OAI222_X1 U85067 ( .A1(n99128), .A2(n120106), .B1(n120100), .B2(n115062), 
        .C1(n113930), .C2(n120094), .ZN(n115081) );
  OAI222_X1 U85068 ( .A1(n99127), .A2(n120106), .B1(n120100), .B2(n115034), 
        .C1(n113929), .C2(n120094), .ZN(n115053) );
  OAI222_X1 U85069 ( .A1(n99126), .A2(n120106), .B1(n120100), .B2(n115006), 
        .C1(n113928), .C2(n120094), .ZN(n115025) );
  OAI222_X1 U85070 ( .A1(n99125), .A2(n120106), .B1(n120100), .B2(n114978), 
        .C1(n113927), .C2(n120094), .ZN(n114997) );
  OAI222_X1 U85071 ( .A1(n99124), .A2(n120106), .B1(n120100), .B2(n114950), 
        .C1(n113926), .C2(n120094), .ZN(n114969) );
  OAI222_X1 U85072 ( .A1(n99123), .A2(n120106), .B1(n120100), .B2(n114922), 
        .C1(n113925), .C2(n120094), .ZN(n114941) );
  OAI222_X1 U85073 ( .A1(n99122), .A2(n120106), .B1(n120100), .B2(n114894), 
        .C1(n113924), .C2(n120094), .ZN(n114913) );
  OAI222_X1 U85074 ( .A1(n99121), .A2(n120106), .B1(n120100), .B2(n114866), 
        .C1(n113923), .C2(n120094), .ZN(n114885) );
  OAI222_X1 U85075 ( .A1(n99120), .A2(n120106), .B1(n120100), .B2(n114838), 
        .C1(n113922), .C2(n120094), .ZN(n114857) );
  OAI222_X1 U85076 ( .A1(n99119), .A2(n120106), .B1(n120100), .B2(n114810), 
        .C1(n113921), .C2(n120094), .ZN(n114829) );
  OAI222_X1 U85077 ( .A1(n99118), .A2(n120106), .B1(n120100), .B2(n114782), 
        .C1(n113920), .C2(n120094), .ZN(n114801) );
  OAI222_X1 U85078 ( .A1(n99177), .A2(n120102), .B1(n120096), .B2(n116434), 
        .C1(n113979), .C2(n120090), .ZN(n116465) );
  OAI222_X1 U85079 ( .A1(n99176), .A2(n120102), .B1(n120096), .B2(n116406), 
        .C1(n113978), .C2(n120090), .ZN(n116425) );
  OAI222_X1 U85080 ( .A1(n99175), .A2(n120102), .B1(n120096), .B2(n116378), 
        .C1(n113977), .C2(n120090), .ZN(n116397) );
  OAI222_X1 U85081 ( .A1(n99174), .A2(n120102), .B1(n120096), .B2(n116350), 
        .C1(n113976), .C2(n120090), .ZN(n116369) );
  OAI222_X1 U85082 ( .A1(n113972), .A2(n119904), .B1(n90363), .B2(n119898), 
        .C1(n99368), .C2(n119892), .ZN(n117797) );
  OAI222_X1 U85083 ( .A1(n113971), .A2(n119904), .B1(n90362), .B2(n119898), 
        .C1(n99367), .C2(n119892), .ZN(n117775) );
  OAI222_X1 U85084 ( .A1(n113970), .A2(n119904), .B1(n90361), .B2(n119898), 
        .C1(n99366), .C2(n119892), .ZN(n117753) );
  OAI222_X1 U85085 ( .A1(n113969), .A2(n119904), .B1(n90360), .B2(n119898), 
        .C1(n99365), .C2(n119892), .ZN(n117731) );
  OAI222_X1 U85086 ( .A1(n113979), .A2(n119904), .B1(n90370), .B2(n119898), 
        .C1(n99375), .C2(n119892), .ZN(n117963) );
  OAI222_X1 U85087 ( .A1(n113978), .A2(n119904), .B1(n90369), .B2(n119898), 
        .C1(n99374), .C2(n119892), .ZN(n117929) );
  OAI222_X1 U85088 ( .A1(n113977), .A2(n119904), .B1(n90368), .B2(n119898), 
        .C1(n99373), .C2(n119892), .ZN(n117907) );
  OAI222_X1 U85089 ( .A1(n113976), .A2(n119904), .B1(n90367), .B2(n119898), 
        .C1(n99372), .C2(n119892), .ZN(n117885) );
  OAI222_X1 U85090 ( .A1(n113975), .A2(n119904), .B1(n90366), .B2(n119898), 
        .C1(n99371), .C2(n119892), .ZN(n117863) );
  OAI222_X1 U85091 ( .A1(n113974), .A2(n119904), .B1(n90365), .B2(n119898), 
        .C1(n99370), .C2(n119892), .ZN(n117841) );
  OAI222_X1 U85092 ( .A1(n113973), .A2(n119904), .B1(n90364), .B2(n119898), 
        .C1(n99369), .C2(n119892), .ZN(n117819) );
  OAI222_X1 U85093 ( .A1(n99173), .A2(n120102), .B1(n120096), .B2(n116322), 
        .C1(n113975), .C2(n120090), .ZN(n116341) );
  OAI222_X1 U85094 ( .A1(n99172), .A2(n120102), .B1(n120096), .B2(n116294), 
        .C1(n113974), .C2(n120090), .ZN(n116313) );
  OAI222_X1 U85095 ( .A1(n99171), .A2(n120102), .B1(n120096), .B2(n116266), 
        .C1(n113973), .C2(n120090), .ZN(n116285) );
  OAI222_X1 U85096 ( .A1(n99170), .A2(n120102), .B1(n120096), .B2(n116238), 
        .C1(n113972), .C2(n120090), .ZN(n116257) );
  OAI222_X1 U85097 ( .A1(n99169), .A2(n120102), .B1(n120096), .B2(n116210), 
        .C1(n113971), .C2(n120090), .ZN(n116229) );
  OAI222_X1 U85098 ( .A1(n99168), .A2(n120102), .B1(n120096), .B2(n116182), 
        .C1(n113970), .C2(n120090), .ZN(n116201) );
  OAI222_X1 U85099 ( .A1(n99167), .A2(n120102), .B1(n120096), .B2(n116154), 
        .C1(n113969), .C2(n120090), .ZN(n116173) );
  OAI222_X1 U85100 ( .A1(n99166), .A2(n120102), .B1(n120096), .B2(n116126), 
        .C1(n113968), .C2(n120090), .ZN(n116145) );
  OAI222_X1 U85101 ( .A1(n99165), .A2(n120103), .B1(n120097), .B2(n116098), 
        .C1(n113967), .C2(n120091), .ZN(n116117) );
  OAI222_X1 U85102 ( .A1(n99164), .A2(n120103), .B1(n120097), .B2(n116070), 
        .C1(n113966), .C2(n120091), .ZN(n116089) );
  OAI222_X1 U85103 ( .A1(n99163), .A2(n120103), .B1(n120097), .B2(n116042), 
        .C1(n113965), .C2(n120091), .ZN(n116061) );
  OAI222_X1 U85104 ( .A1(n99162), .A2(n120103), .B1(n120097), .B2(n116014), 
        .C1(n113964), .C2(n120091), .ZN(n116033) );
  OAI222_X1 U85105 ( .A1(n99161), .A2(n120103), .B1(n120097), .B2(n115986), 
        .C1(n113963), .C2(n120091), .ZN(n116005) );
  OAI222_X1 U85106 ( .A1(n99160), .A2(n120103), .B1(n120097), .B2(n115958), 
        .C1(n113962), .C2(n120091), .ZN(n115977) );
  OAI222_X1 U85107 ( .A1(n99159), .A2(n120103), .B1(n120097), .B2(n115930), 
        .C1(n113961), .C2(n120091), .ZN(n115949) );
  OAI222_X1 U85108 ( .A1(n99158), .A2(n120103), .B1(n120097), .B2(n115902), 
        .C1(n113960), .C2(n120091), .ZN(n115921) );
  OAI222_X1 U85109 ( .A1(n99157), .A2(n120103), .B1(n120097), .B2(n115874), 
        .C1(n113959), .C2(n120091), .ZN(n115893) );
  OAI222_X1 U85110 ( .A1(n99156), .A2(n120103), .B1(n120097), .B2(n115846), 
        .C1(n113958), .C2(n120091), .ZN(n115865) );
  OAI222_X1 U85111 ( .A1(n99155), .A2(n120103), .B1(n120097), .B2(n115818), 
        .C1(n113957), .C2(n120091), .ZN(n115837) );
  OAI222_X1 U85112 ( .A1(n99154), .A2(n120103), .B1(n120097), .B2(n115790), 
        .C1(n113956), .C2(n120091), .ZN(n115809) );
  OAI222_X1 U85113 ( .A1(n99153), .A2(n120104), .B1(n120098), .B2(n115762), 
        .C1(n113955), .C2(n120092), .ZN(n115781) );
  OAI222_X1 U85114 ( .A1(n99152), .A2(n120104), .B1(n120098), .B2(n115734), 
        .C1(n113954), .C2(n120092), .ZN(n115753) );
  OAI222_X1 U85115 ( .A1(n99151), .A2(n120104), .B1(n120098), .B2(n115706), 
        .C1(n113953), .C2(n120092), .ZN(n115725) );
  OAI222_X1 U85116 ( .A1(n99150), .A2(n120104), .B1(n120098), .B2(n115678), 
        .C1(n113952), .C2(n120092), .ZN(n115697) );
  OAI222_X1 U85117 ( .A1(n99149), .A2(n120104), .B1(n120098), .B2(n115650), 
        .C1(n113951), .C2(n120092), .ZN(n115669) );
  OAI222_X1 U85118 ( .A1(n99148), .A2(n120104), .B1(n120098), .B2(n115622), 
        .C1(n113950), .C2(n120092), .ZN(n115641) );
  OAI222_X1 U85119 ( .A1(n99147), .A2(n120104), .B1(n120098), .B2(n115594), 
        .C1(n113949), .C2(n120092), .ZN(n115613) );
  OAI222_X1 U85120 ( .A1(n99146), .A2(n120104), .B1(n120098), .B2(n115566), 
        .C1(n113948), .C2(n120092), .ZN(n115585) );
  OAI222_X1 U85121 ( .A1(n99145), .A2(n120104), .B1(n120098), .B2(n115538), 
        .C1(n113947), .C2(n120092), .ZN(n115557) );
  OAI222_X1 U85122 ( .A1(n99144), .A2(n120104), .B1(n120098), .B2(n115510), 
        .C1(n113946), .C2(n120092), .ZN(n115529) );
  OAI222_X1 U85123 ( .A1(n99143), .A2(n120104), .B1(n120098), .B2(n115482), 
        .C1(n113945), .C2(n120092), .ZN(n115501) );
  OAI222_X1 U85124 ( .A1(n99142), .A2(n120104), .B1(n120098), .B2(n115454), 
        .C1(n113944), .C2(n120092), .ZN(n115473) );
  OAI222_X1 U85125 ( .A1(n99141), .A2(n120105), .B1(n120099), .B2(n115426), 
        .C1(n113943), .C2(n120093), .ZN(n115445) );
  OAI222_X1 U85126 ( .A1(n99140), .A2(n120105), .B1(n120099), .B2(n115398), 
        .C1(n113942), .C2(n120093), .ZN(n115417) );
  OAI222_X1 U85127 ( .A1(n99139), .A2(n120105), .B1(n120099), .B2(n115370), 
        .C1(n113941), .C2(n120093), .ZN(n115389) );
  OAI222_X1 U85128 ( .A1(n99138), .A2(n120105), .B1(n120099), .B2(n115342), 
        .C1(n113940), .C2(n120093), .ZN(n115361) );
  OAI222_X1 U85129 ( .A1(n99137), .A2(n120105), .B1(n120099), .B2(n115314), 
        .C1(n113939), .C2(n120093), .ZN(n115333) );
  OAI222_X1 U85130 ( .A1(n99136), .A2(n120105), .B1(n120099), .B2(n115286), 
        .C1(n113938), .C2(n120093), .ZN(n115305) );
  OAI222_X1 U85131 ( .A1(n99135), .A2(n120105), .B1(n120099), .B2(n115258), 
        .C1(n113937), .C2(n120093), .ZN(n115277) );
  OAI222_X1 U85132 ( .A1(n99134), .A2(n120105), .B1(n120099), .B2(n115230), 
        .C1(n113936), .C2(n120093), .ZN(n115249) );
  OAI222_X1 U85133 ( .A1(n99133), .A2(n120105), .B1(n120099), .B2(n115202), 
        .C1(n113935), .C2(n120093), .ZN(n115221) );
  OAI222_X1 U85134 ( .A1(n99132), .A2(n120105), .B1(n120099), .B2(n115174), 
        .C1(n113934), .C2(n120093), .ZN(n115193) );
  OAI222_X1 U85135 ( .A1(n99117), .A2(n120107), .B1(n120101), .B2(n114756), 
        .C1(n113919), .C2(n120095), .ZN(n114773) );
  OAI222_X1 U85136 ( .A1(n99116), .A2(n120107), .B1(n120101), .B2(n114730), 
        .C1(n113918), .C2(n120095), .ZN(n114747) );
  OAI222_X1 U85137 ( .A1(n99115), .A2(n120107), .B1(n120101), .B2(n114704), 
        .C1(n113917), .C2(n120095), .ZN(n114721) );
  OAI222_X1 U85138 ( .A1(n99113), .A2(n120107), .B1(n114644), .B2(n120101), 
        .C1(n113915), .C2(n120095), .ZN(n114678) );
  OAI222_X1 U85139 ( .A1(n113919), .A2(n119909), .B1(n90310), .B2(n119903), 
        .C1(n99315), .C2(n119897), .ZN(n116589) );
  OAI222_X1 U85140 ( .A1(n113918), .A2(n119909), .B1(n90309), .B2(n119903), 
        .C1(n99314), .C2(n119897), .ZN(n116568) );
  OAI222_X1 U85141 ( .A1(n113917), .A2(n119909), .B1(n90308), .B2(n119903), 
        .C1(n99313), .C2(n119897), .ZN(n116547) );
  OAI222_X1 U85142 ( .A1(n113915), .A2(n119909), .B1(n90306), .B2(n119903), 
        .C1(n99311), .C2(n119897), .ZN(n116509) );
  NOR4_X1 U85143 ( .A1(n117697), .A2(n117698), .A3(n117699), .A4(n117700), 
        .ZN(n117696) );
  OAI221_X1 U85144 ( .B1(n99232), .B2(n119964), .C1(n98896), .C2(n119958), .A(
        n117708), .ZN(n117697) );
  OAI221_X1 U85145 ( .B1(n114497), .B2(n120036), .C1(n99298), .C2(n120030), 
        .A(n117701), .ZN(n117700) );
  OAI221_X1 U85146 ( .B1(n114563), .B2(n119988), .C1(n114199), .C2(n119982), 
        .A(n117706), .ZN(n117698) );
  NOR4_X1 U85147 ( .A1(n117675), .A2(n117676), .A3(n117677), .A4(n117678), 
        .ZN(n117674) );
  OAI221_X1 U85148 ( .B1(n99231), .B2(n119965), .C1(n98895), .C2(n119959), .A(
        n117686), .ZN(n117675) );
  OAI221_X1 U85149 ( .B1(n114496), .B2(n120037), .C1(n99297), .C2(n120031), 
        .A(n117679), .ZN(n117678) );
  OAI221_X1 U85150 ( .B1(n114562), .B2(n119989), .C1(n114198), .C2(n119983), 
        .A(n117684), .ZN(n117676) );
  NOR4_X1 U85151 ( .A1(n117653), .A2(n117654), .A3(n117655), .A4(n117656), 
        .ZN(n117652) );
  OAI221_X1 U85152 ( .B1(n99230), .B2(n119965), .C1(n98894), .C2(n119959), .A(
        n117664), .ZN(n117653) );
  OAI221_X1 U85153 ( .B1(n114495), .B2(n120037), .C1(n99296), .C2(n120031), 
        .A(n117657), .ZN(n117656) );
  OAI221_X1 U85154 ( .B1(n114561), .B2(n119989), .C1(n114197), .C2(n119983), 
        .A(n117662), .ZN(n117654) );
  NOR4_X1 U85155 ( .A1(n117631), .A2(n117632), .A3(n117633), .A4(n117634), 
        .ZN(n117630) );
  OAI221_X1 U85156 ( .B1(n99229), .B2(n119965), .C1(n98893), .C2(n119959), .A(
        n117642), .ZN(n117631) );
  OAI221_X1 U85157 ( .B1(n114494), .B2(n120037), .C1(n99295), .C2(n120031), 
        .A(n117635), .ZN(n117634) );
  OAI221_X1 U85158 ( .B1(n114560), .B2(n119989), .C1(n114196), .C2(n119983), 
        .A(n117640), .ZN(n117632) );
  NOR4_X1 U85159 ( .A1(n117609), .A2(n117610), .A3(n117611), .A4(n117612), 
        .ZN(n117608) );
  OAI221_X1 U85160 ( .B1(n99228), .B2(n119965), .C1(n98892), .C2(n119959), .A(
        n117620), .ZN(n117609) );
  OAI221_X1 U85161 ( .B1(n114493), .B2(n120037), .C1(n99294), .C2(n120031), 
        .A(n117613), .ZN(n117612) );
  OAI221_X1 U85162 ( .B1(n114559), .B2(n119989), .C1(n114195), .C2(n119983), 
        .A(n117618), .ZN(n117610) );
  NOR4_X1 U85163 ( .A1(n117587), .A2(n117588), .A3(n117589), .A4(n117590), 
        .ZN(n117586) );
  OAI221_X1 U85164 ( .B1(n99227), .B2(n119965), .C1(n98891), .C2(n119959), .A(
        n117598), .ZN(n117587) );
  OAI221_X1 U85165 ( .B1(n114492), .B2(n120037), .C1(n99293), .C2(n120031), 
        .A(n117591), .ZN(n117590) );
  OAI221_X1 U85166 ( .B1(n114558), .B2(n119989), .C1(n114194), .C2(n119983), 
        .A(n117596), .ZN(n117588) );
  NOR4_X1 U85167 ( .A1(n117565), .A2(n117566), .A3(n117567), .A4(n117568), 
        .ZN(n117564) );
  OAI221_X1 U85168 ( .B1(n99226), .B2(n119965), .C1(n98890), .C2(n119959), .A(
        n117576), .ZN(n117565) );
  OAI221_X1 U85169 ( .B1(n114491), .B2(n120037), .C1(n99292), .C2(n120031), 
        .A(n117569), .ZN(n117568) );
  OAI221_X1 U85170 ( .B1(n114557), .B2(n119989), .C1(n114193), .C2(n119983), 
        .A(n117574), .ZN(n117566) );
  NOR4_X1 U85171 ( .A1(n117543), .A2(n117544), .A3(n117545), .A4(n117546), 
        .ZN(n117542) );
  OAI221_X1 U85172 ( .B1(n99225), .B2(n119965), .C1(n98889), .C2(n119959), .A(
        n117554), .ZN(n117543) );
  OAI221_X1 U85173 ( .B1(n114490), .B2(n120037), .C1(n99291), .C2(n120031), 
        .A(n117547), .ZN(n117546) );
  OAI221_X1 U85174 ( .B1(n114556), .B2(n119989), .C1(n114192), .C2(n119983), 
        .A(n117552), .ZN(n117544) );
  NOR4_X1 U85175 ( .A1(n117520), .A2(n117521), .A3(n117522), .A4(n117523), 
        .ZN(n117519) );
  OAI221_X1 U85176 ( .B1(n99224), .B2(n119965), .C1(n98888), .C2(n119959), .A(
        n117531), .ZN(n117520) );
  OAI221_X1 U85177 ( .B1(n114489), .B2(n120037), .C1(n99290), .C2(n120031), 
        .A(n117524), .ZN(n117523) );
  OAI221_X1 U85178 ( .B1(n114555), .B2(n119989), .C1(n114191), .C2(n119983), 
        .A(n117529), .ZN(n117521) );
  NOR4_X1 U85179 ( .A1(n117497), .A2(n117498), .A3(n117499), .A4(n117500), 
        .ZN(n117496) );
  OAI221_X1 U85180 ( .B1(n99223), .B2(n119965), .C1(n98887), .C2(n119959), .A(
        n117508), .ZN(n117497) );
  OAI221_X1 U85181 ( .B1(n114488), .B2(n120037), .C1(n99289), .C2(n120031), 
        .A(n117501), .ZN(n117500) );
  OAI221_X1 U85182 ( .B1(n114554), .B2(n119989), .C1(n114190), .C2(n119983), 
        .A(n117506), .ZN(n117498) );
  NOR4_X1 U85183 ( .A1(n117474), .A2(n117475), .A3(n117476), .A4(n117477), 
        .ZN(n117473) );
  OAI221_X1 U85184 ( .B1(n99222), .B2(n119965), .C1(n98886), .C2(n119959), .A(
        n117485), .ZN(n117474) );
  OAI221_X1 U85185 ( .B1(n114487), .B2(n120037), .C1(n99288), .C2(n120031), 
        .A(n117478), .ZN(n117477) );
  OAI221_X1 U85186 ( .B1(n114553), .B2(n119989), .C1(n114189), .C2(n119983), 
        .A(n117483), .ZN(n117475) );
  NOR4_X1 U85187 ( .A1(n117451), .A2(n117452), .A3(n117453), .A4(n117454), 
        .ZN(n117450) );
  OAI221_X1 U85188 ( .B1(n99221), .B2(n119965), .C1(n98885), .C2(n119959), .A(
        n117462), .ZN(n117451) );
  OAI221_X1 U85189 ( .B1(n114486), .B2(n120037), .C1(n99287), .C2(n120031), 
        .A(n117455), .ZN(n117454) );
  OAI221_X1 U85190 ( .B1(n114552), .B2(n119989), .C1(n114188), .C2(n119983), 
        .A(n117460), .ZN(n117452) );
  NOR4_X1 U85191 ( .A1(n117428), .A2(n117429), .A3(n117430), .A4(n117431), 
        .ZN(n117427) );
  OAI221_X1 U85192 ( .B1(n99220), .B2(n119965), .C1(n98884), .C2(n119959), .A(
        n117439), .ZN(n117428) );
  OAI221_X1 U85193 ( .B1(n114485), .B2(n120037), .C1(n99286), .C2(n120031), 
        .A(n117432), .ZN(n117431) );
  OAI221_X1 U85194 ( .B1(n114551), .B2(n119989), .C1(n114187), .C2(n119983), 
        .A(n117437), .ZN(n117429) );
  NOR4_X1 U85195 ( .A1(n117405), .A2(n117406), .A3(n117407), .A4(n117408), 
        .ZN(n117404) );
  OAI221_X1 U85196 ( .B1(n99219), .B2(n119966), .C1(n98883), .C2(n119960), .A(
        n117416), .ZN(n117405) );
  OAI221_X1 U85197 ( .B1(n114484), .B2(n120038), .C1(n99285), .C2(n120032), 
        .A(n117409), .ZN(n117408) );
  OAI221_X1 U85198 ( .B1(n114550), .B2(n119990), .C1(n114186), .C2(n119984), 
        .A(n117414), .ZN(n117406) );
  NOR4_X1 U85199 ( .A1(n117382), .A2(n117383), .A3(n117384), .A4(n117385), 
        .ZN(n117381) );
  OAI221_X1 U85200 ( .B1(n99218), .B2(n119966), .C1(n98882), .C2(n119960), .A(
        n117393), .ZN(n117382) );
  OAI221_X1 U85201 ( .B1(n114483), .B2(n120038), .C1(n99284), .C2(n120032), 
        .A(n117386), .ZN(n117385) );
  OAI221_X1 U85202 ( .B1(n114549), .B2(n119990), .C1(n114185), .C2(n119984), 
        .A(n117391), .ZN(n117383) );
  NOR4_X1 U85203 ( .A1(n117359), .A2(n117360), .A3(n117361), .A4(n117362), 
        .ZN(n117358) );
  OAI221_X1 U85204 ( .B1(n99217), .B2(n119966), .C1(n98881), .C2(n119960), .A(
        n117370), .ZN(n117359) );
  OAI221_X1 U85205 ( .B1(n114482), .B2(n120038), .C1(n99283), .C2(n120032), 
        .A(n117363), .ZN(n117362) );
  OAI221_X1 U85206 ( .B1(n114548), .B2(n119990), .C1(n114184), .C2(n119984), 
        .A(n117368), .ZN(n117360) );
  NOR4_X1 U85207 ( .A1(n117336), .A2(n117337), .A3(n117338), .A4(n117339), 
        .ZN(n117335) );
  OAI221_X1 U85208 ( .B1(n99216), .B2(n119966), .C1(n98880), .C2(n119960), .A(
        n117347), .ZN(n117336) );
  OAI221_X1 U85209 ( .B1(n114481), .B2(n120038), .C1(n99282), .C2(n120032), 
        .A(n117340), .ZN(n117339) );
  OAI221_X1 U85210 ( .B1(n114547), .B2(n119990), .C1(n114183), .C2(n119984), 
        .A(n117345), .ZN(n117337) );
  NOR4_X1 U85211 ( .A1(n117313), .A2(n117314), .A3(n117315), .A4(n117316), 
        .ZN(n117312) );
  OAI221_X1 U85212 ( .B1(n99215), .B2(n119966), .C1(n98879), .C2(n119960), .A(
        n117324), .ZN(n117313) );
  OAI221_X1 U85213 ( .B1(n114480), .B2(n120038), .C1(n99281), .C2(n120032), 
        .A(n117317), .ZN(n117316) );
  OAI221_X1 U85214 ( .B1(n114546), .B2(n119990), .C1(n114182), .C2(n119984), 
        .A(n117322), .ZN(n117314) );
  NOR4_X1 U85215 ( .A1(n117290), .A2(n117291), .A3(n117292), .A4(n117293), 
        .ZN(n117289) );
  OAI221_X1 U85216 ( .B1(n99214), .B2(n119966), .C1(n98878), .C2(n119960), .A(
        n117301), .ZN(n117290) );
  OAI221_X1 U85217 ( .B1(n114479), .B2(n120038), .C1(n99280), .C2(n120032), 
        .A(n117294), .ZN(n117293) );
  OAI221_X1 U85218 ( .B1(n114545), .B2(n119990), .C1(n114181), .C2(n119984), 
        .A(n117299), .ZN(n117291) );
  NOR4_X1 U85219 ( .A1(n117267), .A2(n117268), .A3(n117269), .A4(n117270), 
        .ZN(n117266) );
  OAI221_X1 U85220 ( .B1(n99213), .B2(n119966), .C1(n98877), .C2(n119960), .A(
        n117278), .ZN(n117267) );
  OAI221_X1 U85221 ( .B1(n114478), .B2(n120038), .C1(n99279), .C2(n120032), 
        .A(n117271), .ZN(n117270) );
  OAI221_X1 U85222 ( .B1(n114544), .B2(n119990), .C1(n114180), .C2(n119984), 
        .A(n117276), .ZN(n117268) );
  NOR4_X1 U85223 ( .A1(n117244), .A2(n117245), .A3(n117246), .A4(n117247), 
        .ZN(n117243) );
  OAI221_X1 U85224 ( .B1(n99212), .B2(n119966), .C1(n98876), .C2(n119960), .A(
        n117255), .ZN(n117244) );
  OAI221_X1 U85225 ( .B1(n114477), .B2(n120038), .C1(n99278), .C2(n120032), 
        .A(n117248), .ZN(n117247) );
  OAI221_X1 U85226 ( .B1(n114543), .B2(n119990), .C1(n114179), .C2(n119984), 
        .A(n117253), .ZN(n117245) );
  NOR4_X1 U85227 ( .A1(n117221), .A2(n117222), .A3(n117223), .A4(n117224), 
        .ZN(n117220) );
  OAI221_X1 U85228 ( .B1(n99211), .B2(n119966), .C1(n98875), .C2(n119960), .A(
        n117232), .ZN(n117221) );
  OAI221_X1 U85229 ( .B1(n114476), .B2(n120038), .C1(n99277), .C2(n120032), 
        .A(n117225), .ZN(n117224) );
  OAI221_X1 U85230 ( .B1(n114542), .B2(n119990), .C1(n114178), .C2(n119984), 
        .A(n117230), .ZN(n117222) );
  NOR4_X1 U85231 ( .A1(n117198), .A2(n117199), .A3(n117200), .A4(n117201), 
        .ZN(n117197) );
  OAI221_X1 U85232 ( .B1(n99210), .B2(n119966), .C1(n98874), .C2(n119960), .A(
        n117209), .ZN(n117198) );
  OAI221_X1 U85233 ( .B1(n114475), .B2(n120038), .C1(n99276), .C2(n120032), 
        .A(n117202), .ZN(n117201) );
  OAI221_X1 U85234 ( .B1(n114541), .B2(n119990), .C1(n114177), .C2(n119984), 
        .A(n117207), .ZN(n117199) );
  NOR4_X1 U85235 ( .A1(n117175), .A2(n117176), .A3(n117177), .A4(n117178), 
        .ZN(n117174) );
  OAI221_X1 U85236 ( .B1(n99209), .B2(n119966), .C1(n98873), .C2(n119960), .A(
        n117186), .ZN(n117175) );
  OAI221_X1 U85237 ( .B1(n114474), .B2(n120038), .C1(n99275), .C2(n120032), 
        .A(n117179), .ZN(n117178) );
  OAI221_X1 U85238 ( .B1(n114540), .B2(n119990), .C1(n114176), .C2(n119984), 
        .A(n117184), .ZN(n117176) );
  NOR4_X1 U85239 ( .A1(n117152), .A2(n117153), .A3(n117154), .A4(n117155), 
        .ZN(n117151) );
  OAI221_X1 U85240 ( .B1(n99208), .B2(n119966), .C1(n98872), .C2(n119960), .A(
        n117163), .ZN(n117152) );
  OAI221_X1 U85241 ( .B1(n114473), .B2(n120038), .C1(n99274), .C2(n120032), 
        .A(n117156), .ZN(n117155) );
  OAI221_X1 U85242 ( .B1(n114539), .B2(n119990), .C1(n114175), .C2(n119984), 
        .A(n117161), .ZN(n117153) );
  NOR4_X1 U85243 ( .A1(n117129), .A2(n117130), .A3(n117131), .A4(n117132), 
        .ZN(n117128) );
  OAI221_X1 U85244 ( .B1(n99207), .B2(n119967), .C1(n98871), .C2(n119961), .A(
        n117140), .ZN(n117129) );
  OAI221_X1 U85245 ( .B1(n114472), .B2(n120039), .C1(n99273), .C2(n120033), 
        .A(n117133), .ZN(n117132) );
  OAI221_X1 U85246 ( .B1(n114538), .B2(n119991), .C1(n114174), .C2(n119985), 
        .A(n117138), .ZN(n117130) );
  NOR4_X1 U85247 ( .A1(n117106), .A2(n117107), .A3(n117108), .A4(n117109), 
        .ZN(n117105) );
  OAI221_X1 U85248 ( .B1(n99206), .B2(n119967), .C1(n98870), .C2(n119961), .A(
        n117117), .ZN(n117106) );
  OAI221_X1 U85249 ( .B1(n114471), .B2(n120039), .C1(n99272), .C2(n120033), 
        .A(n117110), .ZN(n117109) );
  OAI221_X1 U85250 ( .B1(n114537), .B2(n119991), .C1(n114173), .C2(n119985), 
        .A(n117115), .ZN(n117107) );
  NOR4_X1 U85251 ( .A1(n117083), .A2(n117084), .A3(n117085), .A4(n117086), 
        .ZN(n117082) );
  OAI221_X1 U85252 ( .B1(n99205), .B2(n119967), .C1(n98869), .C2(n119961), .A(
        n117094), .ZN(n117083) );
  OAI221_X1 U85253 ( .B1(n114470), .B2(n120039), .C1(n99271), .C2(n120033), 
        .A(n117087), .ZN(n117086) );
  OAI221_X1 U85254 ( .B1(n114536), .B2(n119991), .C1(n114172), .C2(n119985), 
        .A(n117092), .ZN(n117084) );
  NOR4_X1 U85255 ( .A1(n117060), .A2(n117061), .A3(n117062), .A4(n117063), 
        .ZN(n117059) );
  OAI221_X1 U85256 ( .B1(n99204), .B2(n119967), .C1(n98868), .C2(n119961), .A(
        n117071), .ZN(n117060) );
  OAI221_X1 U85257 ( .B1(n114469), .B2(n120039), .C1(n99270), .C2(n120033), 
        .A(n117064), .ZN(n117063) );
  OAI221_X1 U85258 ( .B1(n114535), .B2(n119991), .C1(n114171), .C2(n119985), 
        .A(n117069), .ZN(n117061) );
  NOR4_X1 U85259 ( .A1(n117037), .A2(n117038), .A3(n117039), .A4(n117040), 
        .ZN(n117036) );
  OAI221_X1 U85260 ( .B1(n99203), .B2(n119967), .C1(n98867), .C2(n119961), .A(
        n117048), .ZN(n117037) );
  OAI221_X1 U85261 ( .B1(n114468), .B2(n120039), .C1(n99269), .C2(n120033), 
        .A(n117041), .ZN(n117040) );
  OAI221_X1 U85262 ( .B1(n114534), .B2(n119991), .C1(n114170), .C2(n119985), 
        .A(n117046), .ZN(n117038) );
  NOR4_X1 U85263 ( .A1(n117014), .A2(n117015), .A3(n117016), .A4(n117017), 
        .ZN(n117013) );
  OAI221_X1 U85264 ( .B1(n99202), .B2(n119967), .C1(n98866), .C2(n119961), .A(
        n117025), .ZN(n117014) );
  OAI221_X1 U85265 ( .B1(n114467), .B2(n120039), .C1(n99268), .C2(n120033), 
        .A(n117018), .ZN(n117017) );
  OAI221_X1 U85266 ( .B1(n114533), .B2(n119991), .C1(n114169), .C2(n119985), 
        .A(n117023), .ZN(n117015) );
  NOR4_X1 U85267 ( .A1(n116991), .A2(n116992), .A3(n116993), .A4(n116994), 
        .ZN(n116990) );
  OAI221_X1 U85268 ( .B1(n99201), .B2(n119967), .C1(n98865), .C2(n119961), .A(
        n117002), .ZN(n116991) );
  OAI221_X1 U85269 ( .B1(n114466), .B2(n120039), .C1(n99267), .C2(n120033), 
        .A(n116995), .ZN(n116994) );
  OAI221_X1 U85270 ( .B1(n114532), .B2(n119991), .C1(n114168), .C2(n119985), 
        .A(n117000), .ZN(n116992) );
  NOR4_X1 U85271 ( .A1(n116968), .A2(n116969), .A3(n116970), .A4(n116971), 
        .ZN(n116967) );
  OAI221_X1 U85272 ( .B1(n99200), .B2(n119967), .C1(n98864), .C2(n119961), .A(
        n116979), .ZN(n116968) );
  OAI221_X1 U85273 ( .B1(n114465), .B2(n120039), .C1(n99266), .C2(n120033), 
        .A(n116972), .ZN(n116971) );
  OAI221_X1 U85274 ( .B1(n114531), .B2(n119991), .C1(n114167), .C2(n119985), 
        .A(n116977), .ZN(n116969) );
  NOR4_X1 U85275 ( .A1(n116945), .A2(n116946), .A3(n116947), .A4(n116948), 
        .ZN(n116944) );
  OAI221_X1 U85276 ( .B1(n99199), .B2(n119967), .C1(n98863), .C2(n119961), .A(
        n116956), .ZN(n116945) );
  OAI221_X1 U85277 ( .B1(n114464), .B2(n120039), .C1(n99265), .C2(n120033), 
        .A(n116949), .ZN(n116948) );
  OAI221_X1 U85278 ( .B1(n114530), .B2(n119991), .C1(n114166), .C2(n119985), 
        .A(n116954), .ZN(n116946) );
  NOR4_X1 U85279 ( .A1(n116922), .A2(n116923), .A3(n116924), .A4(n116925), 
        .ZN(n116921) );
  OAI221_X1 U85280 ( .B1(n99198), .B2(n119967), .C1(n98862), .C2(n119961), .A(
        n116933), .ZN(n116922) );
  OAI221_X1 U85281 ( .B1(n114463), .B2(n120039), .C1(n99264), .C2(n120033), 
        .A(n116926), .ZN(n116925) );
  OAI221_X1 U85282 ( .B1(n114529), .B2(n119991), .C1(n114165), .C2(n119985), 
        .A(n116931), .ZN(n116923) );
  NOR4_X1 U85283 ( .A1(n116899), .A2(n116900), .A3(n116901), .A4(n116902), 
        .ZN(n116898) );
  OAI221_X1 U85284 ( .B1(n99197), .B2(n119967), .C1(n98861), .C2(n119961), .A(
        n116910), .ZN(n116899) );
  OAI221_X1 U85285 ( .B1(n114462), .B2(n120039), .C1(n99263), .C2(n120033), 
        .A(n116903), .ZN(n116902) );
  OAI221_X1 U85286 ( .B1(n114528), .B2(n119991), .C1(n114164), .C2(n119985), 
        .A(n116908), .ZN(n116900) );
  NOR4_X1 U85287 ( .A1(n116876), .A2(n116877), .A3(n116878), .A4(n116879), 
        .ZN(n116875) );
  OAI221_X1 U85288 ( .B1(n99196), .B2(n119967), .C1(n98860), .C2(n119961), .A(
        n116887), .ZN(n116876) );
  OAI221_X1 U85289 ( .B1(n114461), .B2(n120039), .C1(n99262), .C2(n120033), 
        .A(n116880), .ZN(n116879) );
  OAI221_X1 U85290 ( .B1(n114527), .B2(n119991), .C1(n114163), .C2(n119985), 
        .A(n116885), .ZN(n116877) );
  NOR4_X1 U85291 ( .A1(n116853), .A2(n116854), .A3(n116855), .A4(n116856), 
        .ZN(n116852) );
  OAI221_X1 U85292 ( .B1(n99195), .B2(n119968), .C1(n98859), .C2(n119962), .A(
        n116864), .ZN(n116853) );
  OAI221_X1 U85293 ( .B1(n114460), .B2(n120040), .C1(n99261), .C2(n120034), 
        .A(n116857), .ZN(n116856) );
  OAI221_X1 U85294 ( .B1(n114526), .B2(n119992), .C1(n114162), .C2(n119986), 
        .A(n116862), .ZN(n116854) );
  NOR4_X1 U85295 ( .A1(n116830), .A2(n116831), .A3(n116832), .A4(n116833), 
        .ZN(n116829) );
  OAI221_X1 U85296 ( .B1(n99194), .B2(n119968), .C1(n98858), .C2(n119962), .A(
        n116841), .ZN(n116830) );
  OAI221_X1 U85297 ( .B1(n114459), .B2(n120040), .C1(n99260), .C2(n120034), 
        .A(n116834), .ZN(n116833) );
  OAI221_X1 U85298 ( .B1(n114525), .B2(n119992), .C1(n114161), .C2(n119986), 
        .A(n116839), .ZN(n116831) );
  NOR4_X1 U85299 ( .A1(n116807), .A2(n116808), .A3(n116809), .A4(n116810), 
        .ZN(n116806) );
  OAI221_X1 U85300 ( .B1(n99193), .B2(n119968), .C1(n98857), .C2(n119962), .A(
        n116818), .ZN(n116807) );
  OAI221_X1 U85301 ( .B1(n114458), .B2(n120040), .C1(n99259), .C2(n120034), 
        .A(n116811), .ZN(n116810) );
  OAI221_X1 U85302 ( .B1(n114524), .B2(n119992), .C1(n114160), .C2(n119986), 
        .A(n116816), .ZN(n116808) );
  NOR4_X1 U85303 ( .A1(n116784), .A2(n116785), .A3(n116786), .A4(n116787), 
        .ZN(n116783) );
  OAI221_X1 U85304 ( .B1(n99192), .B2(n119968), .C1(n98856), .C2(n119962), .A(
        n116795), .ZN(n116784) );
  OAI221_X1 U85305 ( .B1(n114457), .B2(n120040), .C1(n99258), .C2(n120034), 
        .A(n116788), .ZN(n116787) );
  OAI221_X1 U85306 ( .B1(n114523), .B2(n119992), .C1(n114159), .C2(n119986), 
        .A(n116793), .ZN(n116785) );
  NOR4_X1 U85307 ( .A1(n116761), .A2(n116762), .A3(n116763), .A4(n116764), 
        .ZN(n116760) );
  OAI221_X1 U85308 ( .B1(n99191), .B2(n119968), .C1(n98855), .C2(n119962), .A(
        n116772), .ZN(n116761) );
  OAI221_X1 U85309 ( .B1(n114456), .B2(n120040), .C1(n99257), .C2(n120034), 
        .A(n116765), .ZN(n116764) );
  OAI221_X1 U85310 ( .B1(n114522), .B2(n119992), .C1(n114158), .C2(n119986), 
        .A(n116770), .ZN(n116762) );
  NOR4_X1 U85311 ( .A1(n116738), .A2(n116739), .A3(n116740), .A4(n116741), 
        .ZN(n116737) );
  OAI221_X1 U85312 ( .B1(n99190), .B2(n119968), .C1(n98854), .C2(n119962), .A(
        n116749), .ZN(n116738) );
  OAI221_X1 U85313 ( .B1(n114455), .B2(n120040), .C1(n99256), .C2(n120034), 
        .A(n116742), .ZN(n116741) );
  OAI221_X1 U85314 ( .B1(n114521), .B2(n119992), .C1(n114157), .C2(n119986), 
        .A(n116747), .ZN(n116739) );
  NOR4_X1 U85315 ( .A1(n116715), .A2(n116716), .A3(n116717), .A4(n116718), 
        .ZN(n116714) );
  OAI221_X1 U85316 ( .B1(n99189), .B2(n119968), .C1(n98853), .C2(n119962), .A(
        n116726), .ZN(n116715) );
  OAI221_X1 U85317 ( .B1(n114454), .B2(n120040), .C1(n99255), .C2(n120034), 
        .A(n116719), .ZN(n116718) );
  OAI221_X1 U85318 ( .B1(n114520), .B2(n119992), .C1(n114156), .C2(n119986), 
        .A(n116724), .ZN(n116716) );
  NOR4_X1 U85319 ( .A1(n116692), .A2(n116693), .A3(n116694), .A4(n116695), 
        .ZN(n116691) );
  OAI221_X1 U85320 ( .B1(n99188), .B2(n119968), .C1(n98852), .C2(n119962), .A(
        n116703), .ZN(n116692) );
  OAI221_X1 U85321 ( .B1(n114453), .B2(n120040), .C1(n99254), .C2(n120034), 
        .A(n116696), .ZN(n116695) );
  OAI221_X1 U85322 ( .B1(n114519), .B2(n119992), .C1(n114155), .C2(n119986), 
        .A(n116701), .ZN(n116693) );
  NOR4_X1 U85323 ( .A1(n116669), .A2(n116670), .A3(n116671), .A4(n116672), 
        .ZN(n116668) );
  OAI221_X1 U85324 ( .B1(n99187), .B2(n119968), .C1(n98851), .C2(n119962), .A(
        n116680), .ZN(n116669) );
  OAI221_X1 U85325 ( .B1(n114452), .B2(n120040), .C1(n99253), .C2(n120034), 
        .A(n116673), .ZN(n116672) );
  OAI221_X1 U85326 ( .B1(n114518), .B2(n119992), .C1(n114154), .C2(n119986), 
        .A(n116678), .ZN(n116670) );
  NOR4_X1 U85327 ( .A1(n116646), .A2(n116647), .A3(n116648), .A4(n116649), 
        .ZN(n116645) );
  OAI221_X1 U85328 ( .B1(n99186), .B2(n119968), .C1(n98850), .C2(n119962), .A(
        n116657), .ZN(n116646) );
  OAI221_X1 U85329 ( .B1(n114451), .B2(n120040), .C1(n99252), .C2(n120034), 
        .A(n116650), .ZN(n116649) );
  OAI221_X1 U85330 ( .B1(n114517), .B2(n119992), .C1(n114153), .C2(n119986), 
        .A(n116655), .ZN(n116647) );
  NOR4_X1 U85331 ( .A1(n116623), .A2(n116624), .A3(n116625), .A4(n116626), 
        .ZN(n116622) );
  OAI221_X1 U85332 ( .B1(n99185), .B2(n119968), .C1(n98849), .C2(n119962), .A(
        n116634), .ZN(n116623) );
  OAI221_X1 U85333 ( .B1(n114450), .B2(n120040), .C1(n99251), .C2(n120034), 
        .A(n116627), .ZN(n116626) );
  OAI221_X1 U85334 ( .B1(n114516), .B2(n119992), .C1(n114152), .C2(n119986), 
        .A(n116632), .ZN(n116624) );
  NOR4_X1 U85335 ( .A1(n116600), .A2(n116601), .A3(n116602), .A4(n116603), 
        .ZN(n116599) );
  OAI221_X1 U85336 ( .B1(n99184), .B2(n119968), .C1(n98848), .C2(n119962), .A(
        n116611), .ZN(n116600) );
  OAI221_X1 U85337 ( .B1(n114449), .B2(n120040), .C1(n99250), .C2(n120034), 
        .A(n116604), .ZN(n116603) );
  OAI221_X1 U85338 ( .B1(n114515), .B2(n119992), .C1(n114151), .C2(n119986), 
        .A(n116609), .ZN(n116601) );
  NOR4_X1 U85339 ( .A1(n115151), .A2(n115152), .A3(n115153), .A4(n115154), 
        .ZN(n115150) );
  OAI221_X1 U85340 ( .B1(n114528), .B2(n120165), .C1(n114462), .C2(n120159), 
        .A(n115162), .ZN(n115151) );
  OAI221_X1 U85341 ( .B1(n98999), .B2(n120189), .C1(n114396), .C2(n120183), 
        .A(n115160), .ZN(n115152) );
  OAI221_X1 U85342 ( .B1(n99598), .B2(n120237), .C1(n114005), .C2(n120231), 
        .A(n115155), .ZN(n115154) );
  NOR4_X1 U85343 ( .A1(n115123), .A2(n115124), .A3(n115125), .A4(n115126), 
        .ZN(n115122) );
  OAI221_X1 U85344 ( .B1(n114527), .B2(n120165), .C1(n114461), .C2(n120159), 
        .A(n115134), .ZN(n115123) );
  OAI221_X1 U85345 ( .B1(n98998), .B2(n120189), .C1(n114395), .C2(n120183), 
        .A(n115132), .ZN(n115124) );
  OAI221_X1 U85346 ( .B1(n99597), .B2(n120237), .C1(n114004), .C2(n120231), 
        .A(n115127), .ZN(n115126) );
  NOR4_X1 U85347 ( .A1(n115095), .A2(n115096), .A3(n115097), .A4(n115098), 
        .ZN(n115094) );
  OAI221_X1 U85348 ( .B1(n114526), .B2(n120166), .C1(n114460), .C2(n120160), 
        .A(n115106), .ZN(n115095) );
  OAI221_X1 U85349 ( .B1(n98997), .B2(n120190), .C1(n114394), .C2(n120184), 
        .A(n115104), .ZN(n115096) );
  OAI221_X1 U85350 ( .B1(n99596), .B2(n120238), .C1(n114003), .C2(n120232), 
        .A(n115099), .ZN(n115098) );
  NOR4_X1 U85351 ( .A1(n115067), .A2(n115068), .A3(n115069), .A4(n115070), 
        .ZN(n115066) );
  OAI221_X1 U85352 ( .B1(n114525), .B2(n120166), .C1(n114459), .C2(n120160), 
        .A(n115078), .ZN(n115067) );
  OAI221_X1 U85353 ( .B1(n98996), .B2(n120190), .C1(n114393), .C2(n120184), 
        .A(n115076), .ZN(n115068) );
  OAI221_X1 U85354 ( .B1(n99595), .B2(n120238), .C1(n114002), .C2(n120232), 
        .A(n115071), .ZN(n115070) );
  NOR4_X1 U85355 ( .A1(n115039), .A2(n115040), .A3(n115041), .A4(n115042), 
        .ZN(n115038) );
  OAI221_X1 U85356 ( .B1(n114524), .B2(n120166), .C1(n114458), .C2(n120160), 
        .A(n115050), .ZN(n115039) );
  OAI221_X1 U85357 ( .B1(n98995), .B2(n120190), .C1(n114392), .C2(n120184), 
        .A(n115048), .ZN(n115040) );
  OAI221_X1 U85358 ( .B1(n99594), .B2(n120238), .C1(n114001), .C2(n120232), 
        .A(n115043), .ZN(n115042) );
  NOR4_X1 U85359 ( .A1(n115011), .A2(n115012), .A3(n115013), .A4(n115014), 
        .ZN(n115010) );
  OAI221_X1 U85360 ( .B1(n114523), .B2(n120166), .C1(n114457), .C2(n120160), 
        .A(n115022), .ZN(n115011) );
  OAI221_X1 U85361 ( .B1(n98994), .B2(n120190), .C1(n114391), .C2(n120184), 
        .A(n115020), .ZN(n115012) );
  OAI221_X1 U85362 ( .B1(n99593), .B2(n120238), .C1(n114000), .C2(n120232), 
        .A(n115015), .ZN(n115014) );
  NOR4_X1 U85363 ( .A1(n114983), .A2(n114984), .A3(n114985), .A4(n114986), 
        .ZN(n114982) );
  OAI221_X1 U85364 ( .B1(n114522), .B2(n120166), .C1(n114456), .C2(n120160), 
        .A(n114994), .ZN(n114983) );
  OAI221_X1 U85365 ( .B1(n98993), .B2(n120190), .C1(n114390), .C2(n120184), 
        .A(n114992), .ZN(n114984) );
  OAI221_X1 U85366 ( .B1(n99592), .B2(n120238), .C1(n113999), .C2(n120232), 
        .A(n114987), .ZN(n114986) );
  NOR4_X1 U85367 ( .A1(n114955), .A2(n114956), .A3(n114957), .A4(n114958), 
        .ZN(n114954) );
  OAI221_X1 U85368 ( .B1(n114521), .B2(n120166), .C1(n114455), .C2(n120160), 
        .A(n114966), .ZN(n114955) );
  OAI221_X1 U85369 ( .B1(n98992), .B2(n120190), .C1(n114389), .C2(n120184), 
        .A(n114964), .ZN(n114956) );
  OAI221_X1 U85370 ( .B1(n99591), .B2(n120238), .C1(n113998), .C2(n120232), 
        .A(n114959), .ZN(n114958) );
  NOR4_X1 U85371 ( .A1(n114927), .A2(n114928), .A3(n114929), .A4(n114930), 
        .ZN(n114926) );
  OAI221_X1 U85372 ( .B1(n114520), .B2(n120166), .C1(n114454), .C2(n120160), 
        .A(n114938), .ZN(n114927) );
  OAI221_X1 U85373 ( .B1(n98991), .B2(n120190), .C1(n114388), .C2(n120184), 
        .A(n114936), .ZN(n114928) );
  OAI221_X1 U85374 ( .B1(n99590), .B2(n120238), .C1(n113997), .C2(n120232), 
        .A(n114931), .ZN(n114930) );
  NOR4_X1 U85375 ( .A1(n114899), .A2(n114900), .A3(n114901), .A4(n114902), 
        .ZN(n114898) );
  OAI221_X1 U85376 ( .B1(n114519), .B2(n120166), .C1(n114453), .C2(n120160), 
        .A(n114910), .ZN(n114899) );
  OAI221_X1 U85377 ( .B1(n98990), .B2(n120190), .C1(n114387), .C2(n120184), 
        .A(n114908), .ZN(n114900) );
  OAI221_X1 U85378 ( .B1(n99589), .B2(n120238), .C1(n113996), .C2(n120232), 
        .A(n114903), .ZN(n114902) );
  NOR4_X1 U85379 ( .A1(n114871), .A2(n114872), .A3(n114873), .A4(n114874), 
        .ZN(n114870) );
  OAI221_X1 U85380 ( .B1(n114518), .B2(n120166), .C1(n114452), .C2(n120160), 
        .A(n114882), .ZN(n114871) );
  OAI221_X1 U85381 ( .B1(n98989), .B2(n120190), .C1(n114386), .C2(n120184), 
        .A(n114880), .ZN(n114872) );
  OAI221_X1 U85382 ( .B1(n99588), .B2(n120238), .C1(n113995), .C2(n120232), 
        .A(n114875), .ZN(n114874) );
  NOR4_X1 U85383 ( .A1(n114843), .A2(n114844), .A3(n114845), .A4(n114846), 
        .ZN(n114842) );
  OAI221_X1 U85384 ( .B1(n114517), .B2(n120166), .C1(n114451), .C2(n120160), 
        .A(n114854), .ZN(n114843) );
  OAI221_X1 U85385 ( .B1(n98988), .B2(n120190), .C1(n114385), .C2(n120184), 
        .A(n114852), .ZN(n114844) );
  OAI221_X1 U85386 ( .B1(n99587), .B2(n120238), .C1(n113994), .C2(n120232), 
        .A(n114847), .ZN(n114846) );
  NOR4_X1 U85387 ( .A1(n114815), .A2(n114816), .A3(n114817), .A4(n114818), 
        .ZN(n114814) );
  OAI221_X1 U85388 ( .B1(n114516), .B2(n120166), .C1(n114450), .C2(n120160), 
        .A(n114826), .ZN(n114815) );
  OAI221_X1 U85389 ( .B1(n98987), .B2(n120190), .C1(n114384), .C2(n120184), 
        .A(n114824), .ZN(n114816) );
  OAI221_X1 U85390 ( .B1(n99586), .B2(n120238), .C1(n113993), .C2(n120232), 
        .A(n114819), .ZN(n114818) );
  NOR4_X1 U85391 ( .A1(n114787), .A2(n114788), .A3(n114789), .A4(n114790), 
        .ZN(n114786) );
  OAI221_X1 U85392 ( .B1(n114515), .B2(n120166), .C1(n114449), .C2(n120160), 
        .A(n114798), .ZN(n114787) );
  OAI221_X1 U85393 ( .B1(n98986), .B2(n120190), .C1(n114383), .C2(n120184), 
        .A(n114796), .ZN(n114788) );
  OAI221_X1 U85394 ( .B1(n99585), .B2(n120238), .C1(n113992), .C2(n120232), 
        .A(n114791), .ZN(n114790) );
  NOR4_X1 U85395 ( .A1(n116439), .A2(n116440), .A3(n116441), .A4(n116442), 
        .ZN(n116438) );
  OAI221_X1 U85396 ( .B1(n114574), .B2(n120162), .C1(n114508), .C2(n120156), 
        .A(n116460), .ZN(n116439) );
  OAI221_X1 U85397 ( .B1(n99045), .B2(n120186), .C1(n114442), .C2(n120180), 
        .A(n116455), .ZN(n116440) );
  OAI221_X1 U85398 ( .B1(n99644), .B2(n120234), .C1(n114051), .C2(n120228), 
        .A(n116443), .ZN(n116442) );
  NOR4_X1 U85399 ( .A1(n116411), .A2(n116412), .A3(n116413), .A4(n116414), 
        .ZN(n116410) );
  OAI221_X1 U85400 ( .B1(n114573), .B2(n120162), .C1(n114507), .C2(n120156), 
        .A(n116422), .ZN(n116411) );
  OAI221_X1 U85401 ( .B1(n99044), .B2(n120186), .C1(n114441), .C2(n120180), 
        .A(n116420), .ZN(n116412) );
  OAI221_X1 U85402 ( .B1(n99643), .B2(n120234), .C1(n114050), .C2(n120228), 
        .A(n116415), .ZN(n116414) );
  NOR4_X1 U85403 ( .A1(n116383), .A2(n116384), .A3(n116385), .A4(n116386), 
        .ZN(n116382) );
  OAI221_X1 U85404 ( .B1(n114572), .B2(n120162), .C1(n114506), .C2(n120156), 
        .A(n116394), .ZN(n116383) );
  OAI221_X1 U85405 ( .B1(n99043), .B2(n120186), .C1(n114440), .C2(n120180), 
        .A(n116392), .ZN(n116384) );
  OAI221_X1 U85406 ( .B1(n99642), .B2(n120234), .C1(n114049), .C2(n120228), 
        .A(n116387), .ZN(n116386) );
  NOR4_X1 U85407 ( .A1(n116355), .A2(n116356), .A3(n116357), .A4(n116358), 
        .ZN(n116354) );
  OAI221_X1 U85408 ( .B1(n114571), .B2(n120162), .C1(n114505), .C2(n120156), 
        .A(n116366), .ZN(n116355) );
  OAI221_X1 U85409 ( .B1(n99042), .B2(n120186), .C1(n114439), .C2(n120180), 
        .A(n116364), .ZN(n116356) );
  OAI221_X1 U85410 ( .B1(n99641), .B2(n120234), .C1(n114048), .C2(n120228), 
        .A(n116359), .ZN(n116358) );
  NOR4_X1 U85411 ( .A1(n117785), .A2(n117786), .A3(n117787), .A4(n117788), 
        .ZN(n117784) );
  OAI221_X1 U85412 ( .B1(n99236), .B2(n119964), .C1(n98900), .C2(n119958), .A(
        n117796), .ZN(n117785) );
  OAI221_X1 U85413 ( .B1(n114501), .B2(n120036), .C1(n99302), .C2(n120030), 
        .A(n117789), .ZN(n117788) );
  OAI221_X1 U85414 ( .B1(n114567), .B2(n119988), .C1(n114203), .C2(n119982), 
        .A(n117794), .ZN(n117786) );
  NOR4_X1 U85415 ( .A1(n117763), .A2(n117764), .A3(n117765), .A4(n117766), 
        .ZN(n117762) );
  OAI221_X1 U85416 ( .B1(n99235), .B2(n119964), .C1(n98899), .C2(n119958), .A(
        n117774), .ZN(n117763) );
  OAI221_X1 U85417 ( .B1(n114500), .B2(n120036), .C1(n99301), .C2(n120030), 
        .A(n117767), .ZN(n117766) );
  OAI221_X1 U85418 ( .B1(n114566), .B2(n119988), .C1(n114202), .C2(n119982), 
        .A(n117772), .ZN(n117764) );
  NOR4_X1 U85419 ( .A1(n117741), .A2(n117742), .A3(n117743), .A4(n117744), 
        .ZN(n117740) );
  OAI221_X1 U85420 ( .B1(n99234), .B2(n119964), .C1(n98898), .C2(n119958), .A(
        n117752), .ZN(n117741) );
  OAI221_X1 U85421 ( .B1(n114499), .B2(n120036), .C1(n99300), .C2(n120030), 
        .A(n117745), .ZN(n117744) );
  OAI221_X1 U85422 ( .B1(n114565), .B2(n119988), .C1(n114201), .C2(n119982), 
        .A(n117750), .ZN(n117742) );
  NOR4_X1 U85423 ( .A1(n117719), .A2(n117720), .A3(n117721), .A4(n117722), 
        .ZN(n117718) );
  OAI221_X1 U85424 ( .B1(n99233), .B2(n119964), .C1(n98897), .C2(n119958), .A(
        n117730), .ZN(n117719) );
  OAI221_X1 U85425 ( .B1(n114498), .B2(n120036), .C1(n99299), .C2(n120030), 
        .A(n117723), .ZN(n117722) );
  OAI221_X1 U85426 ( .B1(n114564), .B2(n119988), .C1(n114200), .C2(n119982), 
        .A(n117728), .ZN(n117720) );
  NOR4_X1 U85427 ( .A1(n117939), .A2(n117940), .A3(n117941), .A4(n117942), 
        .ZN(n117938) );
  OAI221_X1 U85428 ( .B1(n99243), .B2(n119964), .C1(n98907), .C2(n119958), .A(
        n117960), .ZN(n117939) );
  OAI221_X1 U85429 ( .B1(n114508), .B2(n120036), .C1(n99309), .C2(n120030), 
        .A(n117943), .ZN(n117942) );
  OAI221_X1 U85430 ( .B1(n114574), .B2(n119988), .C1(n114210), .C2(n119982), 
        .A(n117956), .ZN(n117940) );
  NOR4_X1 U85431 ( .A1(n117917), .A2(n117918), .A3(n117919), .A4(n117920), 
        .ZN(n117916) );
  OAI221_X1 U85432 ( .B1(n99242), .B2(n119964), .C1(n98906), .C2(n119958), .A(
        n117928), .ZN(n117917) );
  OAI221_X1 U85433 ( .B1(n114507), .B2(n120036), .C1(n99308), .C2(n120030), 
        .A(n117921), .ZN(n117920) );
  OAI221_X1 U85434 ( .B1(n114573), .B2(n119988), .C1(n114209), .C2(n119982), 
        .A(n117926), .ZN(n117918) );
  NOR4_X1 U85435 ( .A1(n117895), .A2(n117896), .A3(n117897), .A4(n117898), 
        .ZN(n117894) );
  OAI221_X1 U85436 ( .B1(n99241), .B2(n119964), .C1(n98905), .C2(n119958), .A(
        n117906), .ZN(n117895) );
  OAI221_X1 U85437 ( .B1(n114506), .B2(n120036), .C1(n99307), .C2(n120030), 
        .A(n117899), .ZN(n117898) );
  OAI221_X1 U85438 ( .B1(n114572), .B2(n119988), .C1(n114208), .C2(n119982), 
        .A(n117904), .ZN(n117896) );
  NOR4_X1 U85439 ( .A1(n117873), .A2(n117874), .A3(n117875), .A4(n117876), 
        .ZN(n117872) );
  OAI221_X1 U85440 ( .B1(n99240), .B2(n119964), .C1(n98904), .C2(n119958), .A(
        n117884), .ZN(n117873) );
  OAI221_X1 U85441 ( .B1(n114505), .B2(n120036), .C1(n99306), .C2(n120030), 
        .A(n117877), .ZN(n117876) );
  OAI221_X1 U85442 ( .B1(n114571), .B2(n119988), .C1(n114207), .C2(n119982), 
        .A(n117882), .ZN(n117874) );
  NOR4_X1 U85443 ( .A1(n117851), .A2(n117852), .A3(n117853), .A4(n117854), 
        .ZN(n117850) );
  OAI221_X1 U85444 ( .B1(n99239), .B2(n119964), .C1(n98903), .C2(n119958), .A(
        n117862), .ZN(n117851) );
  OAI221_X1 U85445 ( .B1(n114504), .B2(n120036), .C1(n99305), .C2(n120030), 
        .A(n117855), .ZN(n117854) );
  OAI221_X1 U85446 ( .B1(n114570), .B2(n119988), .C1(n114206), .C2(n119982), 
        .A(n117860), .ZN(n117852) );
  NOR4_X1 U85447 ( .A1(n117829), .A2(n117830), .A3(n117831), .A4(n117832), 
        .ZN(n117828) );
  OAI221_X1 U85448 ( .B1(n99238), .B2(n119964), .C1(n98902), .C2(n119958), .A(
        n117840), .ZN(n117829) );
  OAI221_X1 U85449 ( .B1(n114503), .B2(n120036), .C1(n99304), .C2(n120030), 
        .A(n117833), .ZN(n117832) );
  OAI221_X1 U85450 ( .B1(n114569), .B2(n119988), .C1(n114205), .C2(n119982), 
        .A(n117838), .ZN(n117830) );
  NOR4_X1 U85451 ( .A1(n117807), .A2(n117808), .A3(n117809), .A4(n117810), 
        .ZN(n117806) );
  OAI221_X1 U85452 ( .B1(n99237), .B2(n119964), .C1(n98901), .C2(n119958), .A(
        n117818), .ZN(n117807) );
  OAI221_X1 U85453 ( .B1(n114502), .B2(n120036), .C1(n99303), .C2(n120030), 
        .A(n117811), .ZN(n117810) );
  OAI221_X1 U85454 ( .B1(n114568), .B2(n119988), .C1(n114204), .C2(n119982), 
        .A(n117816), .ZN(n117808) );
  NOR4_X1 U85455 ( .A1(n116327), .A2(n116328), .A3(n116329), .A4(n116330), 
        .ZN(n116326) );
  OAI221_X1 U85456 ( .B1(n114570), .B2(n120162), .C1(n114504), .C2(n120156), 
        .A(n116338), .ZN(n116327) );
  OAI221_X1 U85457 ( .B1(n99041), .B2(n120186), .C1(n114438), .C2(n120180), 
        .A(n116336), .ZN(n116328) );
  OAI221_X1 U85458 ( .B1(n99640), .B2(n120234), .C1(n114047), .C2(n120228), 
        .A(n116331), .ZN(n116330) );
  NOR4_X1 U85459 ( .A1(n116299), .A2(n116300), .A3(n116301), .A4(n116302), 
        .ZN(n116298) );
  OAI221_X1 U85460 ( .B1(n114569), .B2(n120162), .C1(n114503), .C2(n120156), 
        .A(n116310), .ZN(n116299) );
  OAI221_X1 U85461 ( .B1(n99040), .B2(n120186), .C1(n114437), .C2(n120180), 
        .A(n116308), .ZN(n116300) );
  OAI221_X1 U85462 ( .B1(n99639), .B2(n120234), .C1(n114046), .C2(n120228), 
        .A(n116303), .ZN(n116302) );
  NOR4_X1 U85463 ( .A1(n116271), .A2(n116272), .A3(n116273), .A4(n116274), 
        .ZN(n116270) );
  OAI221_X1 U85464 ( .B1(n114568), .B2(n120162), .C1(n114502), .C2(n120156), 
        .A(n116282), .ZN(n116271) );
  OAI221_X1 U85465 ( .B1(n99039), .B2(n120186), .C1(n114436), .C2(n120180), 
        .A(n116280), .ZN(n116272) );
  OAI221_X1 U85466 ( .B1(n99638), .B2(n120234), .C1(n114045), .C2(n120228), 
        .A(n116275), .ZN(n116274) );
  NOR4_X1 U85467 ( .A1(n116243), .A2(n116244), .A3(n116245), .A4(n116246), 
        .ZN(n116242) );
  OAI221_X1 U85468 ( .B1(n114567), .B2(n120162), .C1(n114501), .C2(n120156), 
        .A(n116254), .ZN(n116243) );
  OAI221_X1 U85469 ( .B1(n99038), .B2(n120186), .C1(n114435), .C2(n120180), 
        .A(n116252), .ZN(n116244) );
  OAI221_X1 U85470 ( .B1(n99637), .B2(n120234), .C1(n114044), .C2(n120228), 
        .A(n116247), .ZN(n116246) );
  NOR4_X1 U85471 ( .A1(n116215), .A2(n116216), .A3(n116217), .A4(n116218), 
        .ZN(n116214) );
  OAI221_X1 U85472 ( .B1(n114566), .B2(n120162), .C1(n114500), .C2(n120156), 
        .A(n116226), .ZN(n116215) );
  OAI221_X1 U85473 ( .B1(n99037), .B2(n120186), .C1(n114434), .C2(n120180), 
        .A(n116224), .ZN(n116216) );
  OAI221_X1 U85474 ( .B1(n99636), .B2(n120234), .C1(n114043), .C2(n120228), 
        .A(n116219), .ZN(n116218) );
  NOR4_X1 U85475 ( .A1(n116187), .A2(n116188), .A3(n116189), .A4(n116190), 
        .ZN(n116186) );
  OAI221_X1 U85476 ( .B1(n114565), .B2(n120162), .C1(n114499), .C2(n120156), 
        .A(n116198), .ZN(n116187) );
  OAI221_X1 U85477 ( .B1(n99036), .B2(n120186), .C1(n114433), .C2(n120180), 
        .A(n116196), .ZN(n116188) );
  OAI221_X1 U85478 ( .B1(n99635), .B2(n120234), .C1(n114042), .C2(n120228), 
        .A(n116191), .ZN(n116190) );
  NOR4_X1 U85479 ( .A1(n116159), .A2(n116160), .A3(n116161), .A4(n116162), 
        .ZN(n116158) );
  OAI221_X1 U85480 ( .B1(n114564), .B2(n120162), .C1(n114498), .C2(n120156), 
        .A(n116170), .ZN(n116159) );
  OAI221_X1 U85481 ( .B1(n99035), .B2(n120186), .C1(n114432), .C2(n120180), 
        .A(n116168), .ZN(n116160) );
  OAI221_X1 U85482 ( .B1(n99634), .B2(n120234), .C1(n114041), .C2(n120228), 
        .A(n116163), .ZN(n116162) );
  NOR4_X1 U85483 ( .A1(n116131), .A2(n116132), .A3(n116133), .A4(n116134), 
        .ZN(n116130) );
  OAI221_X1 U85484 ( .B1(n114563), .B2(n120162), .C1(n114497), .C2(n120156), 
        .A(n116142), .ZN(n116131) );
  OAI221_X1 U85485 ( .B1(n99034), .B2(n120186), .C1(n114431), .C2(n120180), 
        .A(n116140), .ZN(n116132) );
  OAI221_X1 U85486 ( .B1(n99633), .B2(n120234), .C1(n114040), .C2(n120228), 
        .A(n116135), .ZN(n116134) );
  NOR4_X1 U85487 ( .A1(n116103), .A2(n116104), .A3(n116105), .A4(n116106), 
        .ZN(n116102) );
  OAI221_X1 U85488 ( .B1(n114562), .B2(n120163), .C1(n114496), .C2(n120157), 
        .A(n116114), .ZN(n116103) );
  OAI221_X1 U85489 ( .B1(n99033), .B2(n120187), .C1(n114430), .C2(n120181), 
        .A(n116112), .ZN(n116104) );
  OAI221_X1 U85490 ( .B1(n99632), .B2(n120235), .C1(n114039), .C2(n120229), 
        .A(n116107), .ZN(n116106) );
  NOR4_X1 U85491 ( .A1(n116075), .A2(n116076), .A3(n116077), .A4(n116078), 
        .ZN(n116074) );
  OAI221_X1 U85492 ( .B1(n114561), .B2(n120163), .C1(n114495), .C2(n120157), 
        .A(n116086), .ZN(n116075) );
  OAI221_X1 U85493 ( .B1(n99032), .B2(n120187), .C1(n114429), .C2(n120181), 
        .A(n116084), .ZN(n116076) );
  OAI221_X1 U85494 ( .B1(n99631), .B2(n120235), .C1(n114038), .C2(n120229), 
        .A(n116079), .ZN(n116078) );
  NOR4_X1 U85495 ( .A1(n116047), .A2(n116048), .A3(n116049), .A4(n116050), 
        .ZN(n116046) );
  OAI221_X1 U85496 ( .B1(n114560), .B2(n120163), .C1(n114494), .C2(n120157), 
        .A(n116058), .ZN(n116047) );
  OAI221_X1 U85497 ( .B1(n99031), .B2(n120187), .C1(n114428), .C2(n120181), 
        .A(n116056), .ZN(n116048) );
  OAI221_X1 U85498 ( .B1(n99630), .B2(n120235), .C1(n114037), .C2(n120229), 
        .A(n116051), .ZN(n116050) );
  NOR4_X1 U85499 ( .A1(n116019), .A2(n116020), .A3(n116021), .A4(n116022), 
        .ZN(n116018) );
  OAI221_X1 U85500 ( .B1(n114559), .B2(n120163), .C1(n114493), .C2(n120157), 
        .A(n116030), .ZN(n116019) );
  OAI221_X1 U85501 ( .B1(n99030), .B2(n120187), .C1(n114427), .C2(n120181), 
        .A(n116028), .ZN(n116020) );
  OAI221_X1 U85502 ( .B1(n99629), .B2(n120235), .C1(n114036), .C2(n120229), 
        .A(n116023), .ZN(n116022) );
  NOR4_X1 U85503 ( .A1(n115991), .A2(n115992), .A3(n115993), .A4(n115994), 
        .ZN(n115990) );
  OAI221_X1 U85504 ( .B1(n114558), .B2(n120163), .C1(n114492), .C2(n120157), 
        .A(n116002), .ZN(n115991) );
  OAI221_X1 U85505 ( .B1(n99029), .B2(n120187), .C1(n114426), .C2(n120181), 
        .A(n116000), .ZN(n115992) );
  OAI221_X1 U85506 ( .B1(n99628), .B2(n120235), .C1(n114035), .C2(n120229), 
        .A(n115995), .ZN(n115994) );
  NOR4_X1 U85507 ( .A1(n115963), .A2(n115964), .A3(n115965), .A4(n115966), 
        .ZN(n115962) );
  OAI221_X1 U85508 ( .B1(n114557), .B2(n120163), .C1(n114491), .C2(n120157), 
        .A(n115974), .ZN(n115963) );
  OAI221_X1 U85509 ( .B1(n99028), .B2(n120187), .C1(n114425), .C2(n120181), 
        .A(n115972), .ZN(n115964) );
  OAI221_X1 U85510 ( .B1(n99627), .B2(n120235), .C1(n114034), .C2(n120229), 
        .A(n115967), .ZN(n115966) );
  NOR4_X1 U85511 ( .A1(n115935), .A2(n115936), .A3(n115937), .A4(n115938), 
        .ZN(n115934) );
  OAI221_X1 U85512 ( .B1(n114556), .B2(n120163), .C1(n114490), .C2(n120157), 
        .A(n115946), .ZN(n115935) );
  OAI221_X1 U85513 ( .B1(n99027), .B2(n120187), .C1(n114424), .C2(n120181), 
        .A(n115944), .ZN(n115936) );
  OAI221_X1 U85514 ( .B1(n99626), .B2(n120235), .C1(n114033), .C2(n120229), 
        .A(n115939), .ZN(n115938) );
  NOR4_X1 U85515 ( .A1(n115907), .A2(n115908), .A3(n115909), .A4(n115910), 
        .ZN(n115906) );
  OAI221_X1 U85516 ( .B1(n114555), .B2(n120163), .C1(n114489), .C2(n120157), 
        .A(n115918), .ZN(n115907) );
  OAI221_X1 U85517 ( .B1(n99026), .B2(n120187), .C1(n114423), .C2(n120181), 
        .A(n115916), .ZN(n115908) );
  OAI221_X1 U85518 ( .B1(n99625), .B2(n120235), .C1(n114032), .C2(n120229), 
        .A(n115911), .ZN(n115910) );
  NOR4_X1 U85519 ( .A1(n115879), .A2(n115880), .A3(n115881), .A4(n115882), 
        .ZN(n115878) );
  OAI221_X1 U85520 ( .B1(n114554), .B2(n120163), .C1(n114488), .C2(n120157), 
        .A(n115890), .ZN(n115879) );
  OAI221_X1 U85521 ( .B1(n99025), .B2(n120187), .C1(n114422), .C2(n120181), 
        .A(n115888), .ZN(n115880) );
  OAI221_X1 U85522 ( .B1(n99624), .B2(n120235), .C1(n114031), .C2(n120229), 
        .A(n115883), .ZN(n115882) );
  NOR4_X1 U85523 ( .A1(n115851), .A2(n115852), .A3(n115853), .A4(n115854), 
        .ZN(n115850) );
  OAI221_X1 U85524 ( .B1(n114553), .B2(n120163), .C1(n114487), .C2(n120157), 
        .A(n115862), .ZN(n115851) );
  OAI221_X1 U85525 ( .B1(n99024), .B2(n120187), .C1(n114421), .C2(n120181), 
        .A(n115860), .ZN(n115852) );
  OAI221_X1 U85526 ( .B1(n99623), .B2(n120235), .C1(n114030), .C2(n120229), 
        .A(n115855), .ZN(n115854) );
  NOR4_X1 U85527 ( .A1(n115823), .A2(n115824), .A3(n115825), .A4(n115826), 
        .ZN(n115822) );
  OAI221_X1 U85528 ( .B1(n114552), .B2(n120163), .C1(n114486), .C2(n120157), 
        .A(n115834), .ZN(n115823) );
  OAI221_X1 U85529 ( .B1(n99023), .B2(n120187), .C1(n114420), .C2(n120181), 
        .A(n115832), .ZN(n115824) );
  OAI221_X1 U85530 ( .B1(n99622), .B2(n120235), .C1(n114029), .C2(n120229), 
        .A(n115827), .ZN(n115826) );
  NOR4_X1 U85531 ( .A1(n115795), .A2(n115796), .A3(n115797), .A4(n115798), 
        .ZN(n115794) );
  OAI221_X1 U85532 ( .B1(n114551), .B2(n120163), .C1(n114485), .C2(n120157), 
        .A(n115806), .ZN(n115795) );
  OAI221_X1 U85533 ( .B1(n99022), .B2(n120187), .C1(n114419), .C2(n120181), 
        .A(n115804), .ZN(n115796) );
  OAI221_X1 U85534 ( .B1(n99621), .B2(n120235), .C1(n114028), .C2(n120229), 
        .A(n115799), .ZN(n115798) );
  NOR4_X1 U85535 ( .A1(n115767), .A2(n115768), .A3(n115769), .A4(n115770), 
        .ZN(n115766) );
  OAI221_X1 U85536 ( .B1(n114550), .B2(n120164), .C1(n114484), .C2(n120158), 
        .A(n115778), .ZN(n115767) );
  OAI221_X1 U85537 ( .B1(n99021), .B2(n120188), .C1(n114418), .C2(n120182), 
        .A(n115776), .ZN(n115768) );
  OAI221_X1 U85538 ( .B1(n99620), .B2(n120236), .C1(n114027), .C2(n120230), 
        .A(n115771), .ZN(n115770) );
  NOR4_X1 U85539 ( .A1(n115739), .A2(n115740), .A3(n115741), .A4(n115742), 
        .ZN(n115738) );
  OAI221_X1 U85540 ( .B1(n114549), .B2(n120164), .C1(n114483), .C2(n120158), 
        .A(n115750), .ZN(n115739) );
  OAI221_X1 U85541 ( .B1(n99020), .B2(n120188), .C1(n114417), .C2(n120182), 
        .A(n115748), .ZN(n115740) );
  OAI221_X1 U85542 ( .B1(n99619), .B2(n120236), .C1(n114026), .C2(n120230), 
        .A(n115743), .ZN(n115742) );
  NOR4_X1 U85543 ( .A1(n115711), .A2(n115712), .A3(n115713), .A4(n115714), 
        .ZN(n115710) );
  OAI221_X1 U85544 ( .B1(n114548), .B2(n120164), .C1(n114482), .C2(n120158), 
        .A(n115722), .ZN(n115711) );
  OAI221_X1 U85545 ( .B1(n99019), .B2(n120188), .C1(n114416), .C2(n120182), 
        .A(n115720), .ZN(n115712) );
  OAI221_X1 U85546 ( .B1(n99618), .B2(n120236), .C1(n114025), .C2(n120230), 
        .A(n115715), .ZN(n115714) );
  NOR4_X1 U85547 ( .A1(n115683), .A2(n115684), .A3(n115685), .A4(n115686), 
        .ZN(n115682) );
  OAI221_X1 U85548 ( .B1(n114547), .B2(n120164), .C1(n114481), .C2(n120158), 
        .A(n115694), .ZN(n115683) );
  OAI221_X1 U85549 ( .B1(n99018), .B2(n120188), .C1(n114415), .C2(n120182), 
        .A(n115692), .ZN(n115684) );
  OAI221_X1 U85550 ( .B1(n99617), .B2(n120236), .C1(n114024), .C2(n120230), 
        .A(n115687), .ZN(n115686) );
  NOR4_X1 U85551 ( .A1(n115655), .A2(n115656), .A3(n115657), .A4(n115658), 
        .ZN(n115654) );
  OAI221_X1 U85552 ( .B1(n114546), .B2(n120164), .C1(n114480), .C2(n120158), 
        .A(n115666), .ZN(n115655) );
  OAI221_X1 U85553 ( .B1(n99017), .B2(n120188), .C1(n114414), .C2(n120182), 
        .A(n115664), .ZN(n115656) );
  OAI221_X1 U85554 ( .B1(n99616), .B2(n120236), .C1(n114023), .C2(n120230), 
        .A(n115659), .ZN(n115658) );
  NOR4_X1 U85555 ( .A1(n115627), .A2(n115628), .A3(n115629), .A4(n115630), 
        .ZN(n115626) );
  OAI221_X1 U85556 ( .B1(n114545), .B2(n120164), .C1(n114479), .C2(n120158), 
        .A(n115638), .ZN(n115627) );
  OAI221_X1 U85557 ( .B1(n99016), .B2(n120188), .C1(n114413), .C2(n120182), 
        .A(n115636), .ZN(n115628) );
  OAI221_X1 U85558 ( .B1(n99615), .B2(n120236), .C1(n114022), .C2(n120230), 
        .A(n115631), .ZN(n115630) );
  NOR4_X1 U85559 ( .A1(n115599), .A2(n115600), .A3(n115601), .A4(n115602), 
        .ZN(n115598) );
  OAI221_X1 U85560 ( .B1(n114544), .B2(n120164), .C1(n114478), .C2(n120158), 
        .A(n115610), .ZN(n115599) );
  OAI221_X1 U85561 ( .B1(n99015), .B2(n120188), .C1(n114412), .C2(n120182), 
        .A(n115608), .ZN(n115600) );
  OAI221_X1 U85562 ( .B1(n99614), .B2(n120236), .C1(n114021), .C2(n120230), 
        .A(n115603), .ZN(n115602) );
  NOR4_X1 U85563 ( .A1(n115571), .A2(n115572), .A3(n115573), .A4(n115574), 
        .ZN(n115570) );
  OAI221_X1 U85564 ( .B1(n114543), .B2(n120164), .C1(n114477), .C2(n120158), 
        .A(n115582), .ZN(n115571) );
  OAI221_X1 U85565 ( .B1(n99014), .B2(n120188), .C1(n114411), .C2(n120182), 
        .A(n115580), .ZN(n115572) );
  OAI221_X1 U85566 ( .B1(n99613), .B2(n120236), .C1(n114020), .C2(n120230), 
        .A(n115575), .ZN(n115574) );
  NOR4_X1 U85567 ( .A1(n115543), .A2(n115544), .A3(n115545), .A4(n115546), 
        .ZN(n115542) );
  OAI221_X1 U85568 ( .B1(n114542), .B2(n120164), .C1(n114476), .C2(n120158), 
        .A(n115554), .ZN(n115543) );
  OAI221_X1 U85569 ( .B1(n99013), .B2(n120188), .C1(n114410), .C2(n120182), 
        .A(n115552), .ZN(n115544) );
  OAI221_X1 U85570 ( .B1(n99612), .B2(n120236), .C1(n114019), .C2(n120230), 
        .A(n115547), .ZN(n115546) );
  NOR4_X1 U85571 ( .A1(n115515), .A2(n115516), .A3(n115517), .A4(n115518), 
        .ZN(n115514) );
  OAI221_X1 U85572 ( .B1(n114541), .B2(n120164), .C1(n114475), .C2(n120158), 
        .A(n115526), .ZN(n115515) );
  OAI221_X1 U85573 ( .B1(n99012), .B2(n120188), .C1(n114409), .C2(n120182), 
        .A(n115524), .ZN(n115516) );
  OAI221_X1 U85574 ( .B1(n99611), .B2(n120236), .C1(n114018), .C2(n120230), 
        .A(n115519), .ZN(n115518) );
  NOR4_X1 U85575 ( .A1(n115487), .A2(n115488), .A3(n115489), .A4(n115490), 
        .ZN(n115486) );
  OAI221_X1 U85576 ( .B1(n114540), .B2(n120164), .C1(n114474), .C2(n120158), 
        .A(n115498), .ZN(n115487) );
  OAI221_X1 U85577 ( .B1(n99011), .B2(n120188), .C1(n114408), .C2(n120182), 
        .A(n115496), .ZN(n115488) );
  OAI221_X1 U85578 ( .B1(n99610), .B2(n120236), .C1(n114017), .C2(n120230), 
        .A(n115491), .ZN(n115490) );
  NOR4_X1 U85579 ( .A1(n115459), .A2(n115460), .A3(n115461), .A4(n115462), 
        .ZN(n115458) );
  OAI221_X1 U85580 ( .B1(n114539), .B2(n120164), .C1(n114473), .C2(n120158), 
        .A(n115470), .ZN(n115459) );
  OAI221_X1 U85581 ( .B1(n99010), .B2(n120188), .C1(n114407), .C2(n120182), 
        .A(n115468), .ZN(n115460) );
  OAI221_X1 U85582 ( .B1(n99609), .B2(n120236), .C1(n114016), .C2(n120230), 
        .A(n115463), .ZN(n115462) );
  NOR4_X1 U85583 ( .A1(n115431), .A2(n115432), .A3(n115433), .A4(n115434), 
        .ZN(n115430) );
  OAI221_X1 U85584 ( .B1(n114538), .B2(n120165), .C1(n114472), .C2(n120159), 
        .A(n115442), .ZN(n115431) );
  OAI221_X1 U85585 ( .B1(n99009), .B2(n120189), .C1(n114406), .C2(n120183), 
        .A(n115440), .ZN(n115432) );
  OAI221_X1 U85586 ( .B1(n99608), .B2(n120237), .C1(n114015), .C2(n120231), 
        .A(n115435), .ZN(n115434) );
  NOR4_X1 U85587 ( .A1(n115403), .A2(n115404), .A3(n115405), .A4(n115406), 
        .ZN(n115402) );
  OAI221_X1 U85588 ( .B1(n114537), .B2(n120165), .C1(n114471), .C2(n120159), 
        .A(n115414), .ZN(n115403) );
  OAI221_X1 U85589 ( .B1(n99008), .B2(n120189), .C1(n114405), .C2(n120183), 
        .A(n115412), .ZN(n115404) );
  OAI221_X1 U85590 ( .B1(n99607), .B2(n120237), .C1(n114014), .C2(n120231), 
        .A(n115407), .ZN(n115406) );
  NOR4_X1 U85591 ( .A1(n115375), .A2(n115376), .A3(n115377), .A4(n115378), 
        .ZN(n115374) );
  OAI221_X1 U85592 ( .B1(n114536), .B2(n120165), .C1(n114470), .C2(n120159), 
        .A(n115386), .ZN(n115375) );
  OAI221_X1 U85593 ( .B1(n99007), .B2(n120189), .C1(n114404), .C2(n120183), 
        .A(n115384), .ZN(n115376) );
  OAI221_X1 U85594 ( .B1(n99606), .B2(n120237), .C1(n114013), .C2(n120231), 
        .A(n115379), .ZN(n115378) );
  NOR4_X1 U85595 ( .A1(n115347), .A2(n115348), .A3(n115349), .A4(n115350), 
        .ZN(n115346) );
  OAI221_X1 U85596 ( .B1(n114535), .B2(n120165), .C1(n114469), .C2(n120159), 
        .A(n115358), .ZN(n115347) );
  OAI221_X1 U85597 ( .B1(n99006), .B2(n120189), .C1(n114403), .C2(n120183), 
        .A(n115356), .ZN(n115348) );
  OAI221_X1 U85598 ( .B1(n99605), .B2(n120237), .C1(n114012), .C2(n120231), 
        .A(n115351), .ZN(n115350) );
  NOR4_X1 U85599 ( .A1(n115319), .A2(n115320), .A3(n115321), .A4(n115322), 
        .ZN(n115318) );
  OAI221_X1 U85600 ( .B1(n114534), .B2(n120165), .C1(n114468), .C2(n120159), 
        .A(n115330), .ZN(n115319) );
  OAI221_X1 U85601 ( .B1(n99005), .B2(n120189), .C1(n114402), .C2(n120183), 
        .A(n115328), .ZN(n115320) );
  OAI221_X1 U85602 ( .B1(n99604), .B2(n120237), .C1(n114011), .C2(n120231), 
        .A(n115323), .ZN(n115322) );
  NOR4_X1 U85603 ( .A1(n115291), .A2(n115292), .A3(n115293), .A4(n115294), 
        .ZN(n115290) );
  OAI221_X1 U85604 ( .B1(n114533), .B2(n120165), .C1(n114467), .C2(n120159), 
        .A(n115302), .ZN(n115291) );
  OAI221_X1 U85605 ( .B1(n99004), .B2(n120189), .C1(n114401), .C2(n120183), 
        .A(n115300), .ZN(n115292) );
  OAI221_X1 U85606 ( .B1(n99603), .B2(n120237), .C1(n114010), .C2(n120231), 
        .A(n115295), .ZN(n115294) );
  NOR4_X1 U85607 ( .A1(n115263), .A2(n115264), .A3(n115265), .A4(n115266), 
        .ZN(n115262) );
  OAI221_X1 U85608 ( .B1(n114532), .B2(n120165), .C1(n114466), .C2(n120159), 
        .A(n115274), .ZN(n115263) );
  OAI221_X1 U85609 ( .B1(n99003), .B2(n120189), .C1(n114400), .C2(n120183), 
        .A(n115272), .ZN(n115264) );
  OAI221_X1 U85610 ( .B1(n99602), .B2(n120237), .C1(n114009), .C2(n120231), 
        .A(n115267), .ZN(n115266) );
  NOR4_X1 U85611 ( .A1(n115235), .A2(n115236), .A3(n115237), .A4(n115238), 
        .ZN(n115234) );
  OAI221_X1 U85612 ( .B1(n114531), .B2(n120165), .C1(n114465), .C2(n120159), 
        .A(n115246), .ZN(n115235) );
  OAI221_X1 U85613 ( .B1(n99002), .B2(n120189), .C1(n114399), .C2(n120183), 
        .A(n115244), .ZN(n115236) );
  OAI221_X1 U85614 ( .B1(n99601), .B2(n120237), .C1(n114008), .C2(n120231), 
        .A(n115239), .ZN(n115238) );
  NOR4_X1 U85615 ( .A1(n115207), .A2(n115208), .A3(n115209), .A4(n115210), 
        .ZN(n115206) );
  OAI221_X1 U85616 ( .B1(n114530), .B2(n120165), .C1(n114464), .C2(n120159), 
        .A(n115218), .ZN(n115207) );
  OAI221_X1 U85617 ( .B1(n99001), .B2(n120189), .C1(n114398), .C2(n120183), 
        .A(n115216), .ZN(n115208) );
  OAI221_X1 U85618 ( .B1(n99600), .B2(n120237), .C1(n114007), .C2(n120231), 
        .A(n115211), .ZN(n115210) );
  NOR4_X1 U85619 ( .A1(n115179), .A2(n115180), .A3(n115181), .A4(n115182), 
        .ZN(n115178) );
  OAI221_X1 U85620 ( .B1(n114529), .B2(n120165), .C1(n114463), .C2(n120159), 
        .A(n115190), .ZN(n115179) );
  OAI221_X1 U85621 ( .B1(n99000), .B2(n120189), .C1(n114397), .C2(n120183), 
        .A(n115188), .ZN(n115180) );
  OAI221_X1 U85622 ( .B1(n99599), .B2(n120237), .C1(n114006), .C2(n120231), 
        .A(n115183), .ZN(n115182) );
  AOI221_X1 U85623 ( .B1(n120089), .B2(n118982), .C1(n120083), .C2(n118546), 
        .A(n114779), .ZN(n114758) );
  OAI22_X1 U85624 ( .A1(n98718), .A2(n120077), .B1(n99918), .B2(n120071), .ZN(
        n114779) );
  AOI221_X1 U85625 ( .B1(n120089), .B2(n118983), .C1(n120083), .C2(n118547), 
        .A(n114753), .ZN(n114732) );
  OAI22_X1 U85626 ( .A1(n98717), .A2(n120077), .B1(n99917), .B2(n120071), .ZN(
        n114753) );
  AOI221_X1 U85627 ( .B1(n120089), .B2(n118984), .C1(n120083), .C2(n118548), 
        .A(n114727), .ZN(n114706) );
  OAI22_X1 U85628 ( .A1(n98716), .A2(n120077), .B1(n99916), .B2(n120071), .ZN(
        n114727) );
  AOI221_X1 U85629 ( .B1(n120089), .B2(n118985), .C1(n120083), .C2(n118549), 
        .A(n114695), .ZN(n114647) );
  OAI22_X1 U85630 ( .A1(n98714), .A2(n120077), .B1(n99914), .B2(n120071), .ZN(
        n114695) );
  AOI221_X1 U85631 ( .B1(n119867), .B2(n95525), .C1(n119861), .C2(n117985), 
        .A(n116595), .ZN(n116575) );
  OAI22_X1 U85632 ( .A1(n98652), .A2(n119855), .B1(n99584), .B2(n119849), .ZN(
        n116595) );
  AOI221_X1 U85633 ( .B1(n119867), .B2(n95526), .C1(n119861), .C2(n117986), 
        .A(n116574), .ZN(n116554) );
  OAI22_X1 U85634 ( .A1(n98651), .A2(n119855), .B1(n99583), .B2(n119849), .ZN(
        n116574) );
  AOI221_X1 U85635 ( .B1(n119867), .B2(n95527), .C1(n119861), .C2(n117987), 
        .A(n116553), .ZN(n116533) );
  OAI22_X1 U85636 ( .A1(n98650), .A2(n119855), .B1(n99582), .B2(n119849), .ZN(
        n116553) );
  AOI221_X1 U85637 ( .B1(n119867), .B2(n95528), .C1(n119861), .C2(n117988), 
        .A(n116530), .ZN(n116479) );
  OAI22_X1 U85638 ( .A1(n98648), .A2(n119855), .B1(n99580), .B2(n119849), .ZN(
        n116530) );
  NAND2_X1 U85639 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .ZN(n113986) );
  NAND2_X1 U85640 ( .A1(ADD_WR[1]), .A2(n114375), .ZN(n113908) );
  NAND2_X1 U85641 ( .A1(ADD_WR[2]), .A2(n114376), .ZN(n113913) );
  OAI221_X1 U85642 ( .B1(n99584), .B2(n120239), .C1(n89969), .C2(n120233), .A(
        n114765), .ZN(n114764) );
  AOI22_X1 U85643 ( .A1(n120227), .A2(n109895), .B1(n120216), .B2(OUT1[60]), 
        .ZN(n114765) );
  OAI221_X1 U85644 ( .B1(n99583), .B2(n120239), .C1(n89968), .C2(n120233), .A(
        n114739), .ZN(n114738) );
  AOI22_X1 U85645 ( .A1(n120227), .A2(n109896), .B1(n120216), .B2(OUT1[61]), 
        .ZN(n114739) );
  OAI221_X1 U85646 ( .B1(n99582), .B2(n120239), .C1(n89967), .C2(n120233), .A(
        n114713), .ZN(n114712) );
  AOI22_X1 U85647 ( .A1(n120227), .A2(n109897), .B1(n120216), .B2(OUT1[62]), 
        .ZN(n114713) );
  OAI221_X1 U85648 ( .B1(n99580), .B2(n120239), .C1(n89965), .C2(n120233), .A(
        n114656), .ZN(n114653) );
  AOI22_X1 U85649 ( .A1(n120227), .A2(n109898), .B1(n120218), .B2(OUT1[63]), 
        .ZN(n114656) );
  OAI221_X1 U85650 ( .B1(n114448), .B2(n120041), .C1(n99249), .C2(n120035), 
        .A(n116583), .ZN(n116582) );
  AOI22_X1 U85651 ( .A1(n120029), .A2(n109903), .B1(n120018), .B2(OUT2[60]), 
        .ZN(n116583) );
  OAI221_X1 U85652 ( .B1(n114447), .B2(n120041), .C1(n99248), .C2(n120035), 
        .A(n116562), .ZN(n116561) );
  AOI22_X1 U85653 ( .A1(n120029), .A2(n109904), .B1(n120018), .B2(OUT2[61]), 
        .ZN(n116562) );
  OAI221_X1 U85654 ( .B1(n114446), .B2(n120041), .C1(n99247), .C2(n120035), 
        .A(n116541), .ZN(n116540) );
  AOI22_X1 U85655 ( .A1(n120029), .A2(n109905), .B1(n120018), .B2(OUT2[62]), 
        .ZN(n116541) );
  OAI221_X1 U85656 ( .B1(n114444), .B2(n120041), .C1(n99245), .C2(n120035), 
        .A(n116489), .ZN(n116486) );
  AOI22_X1 U85657 ( .A1(n120029), .A2(n109906), .B1(n120020), .B2(OUT2[63]), 
        .ZN(n116489) );
  OAI221_X1 U85658 ( .B1(n114164), .B2(n120213), .C1(n98666), .C2(n120207), 
        .A(n115157), .ZN(n115153) );
  AOI22_X1 U85659 ( .A1(n120201), .A2(n118610), .B1(n120195), .B2(n119238), 
        .ZN(n115157) );
  OAI221_X1 U85660 ( .B1(n114163), .B2(n120213), .C1(n98665), .C2(n120207), 
        .A(n115129), .ZN(n115125) );
  AOI22_X1 U85661 ( .A1(n120201), .A2(n118611), .B1(n120195), .B2(n119239), 
        .ZN(n115129) );
  OAI221_X1 U85662 ( .B1(n114162), .B2(n120214), .C1(n98664), .C2(n120208), 
        .A(n115101), .ZN(n115097) );
  AOI22_X1 U85663 ( .A1(n120202), .A2(n118612), .B1(n120196), .B2(n119240), 
        .ZN(n115101) );
  OAI221_X1 U85664 ( .B1(n114161), .B2(n120214), .C1(n98663), .C2(n120208), 
        .A(n115073), .ZN(n115069) );
  AOI22_X1 U85665 ( .A1(n120202), .A2(n118613), .B1(n120196), .B2(n119241), 
        .ZN(n115073) );
  OAI221_X1 U85666 ( .B1(n114160), .B2(n120214), .C1(n98662), .C2(n120208), 
        .A(n115045), .ZN(n115041) );
  AOI22_X1 U85667 ( .A1(n120202), .A2(n118614), .B1(n120196), .B2(n119242), 
        .ZN(n115045) );
  OAI221_X1 U85668 ( .B1(n114159), .B2(n120214), .C1(n98661), .C2(n120208), 
        .A(n115017), .ZN(n115013) );
  AOI22_X1 U85669 ( .A1(n120202), .A2(n118615), .B1(n120196), .B2(n119243), 
        .ZN(n115017) );
  OAI221_X1 U85670 ( .B1(n114158), .B2(n120214), .C1(n98660), .C2(n120208), 
        .A(n114989), .ZN(n114985) );
  AOI22_X1 U85671 ( .A1(n120202), .A2(n118616), .B1(n120196), .B2(n119244), 
        .ZN(n114989) );
  OAI221_X1 U85672 ( .B1(n114157), .B2(n120214), .C1(n98659), .C2(n120208), 
        .A(n114961), .ZN(n114957) );
  AOI22_X1 U85673 ( .A1(n120202), .A2(n118617), .B1(n120196), .B2(n119245), 
        .ZN(n114961) );
  OAI221_X1 U85674 ( .B1(n114156), .B2(n120214), .C1(n98658), .C2(n120208), 
        .A(n114933), .ZN(n114929) );
  AOI22_X1 U85675 ( .A1(n120202), .A2(n118618), .B1(n120196), .B2(n119246), 
        .ZN(n114933) );
  OAI221_X1 U85676 ( .B1(n114155), .B2(n120214), .C1(n98657), .C2(n120208), 
        .A(n114905), .ZN(n114901) );
  AOI22_X1 U85677 ( .A1(n120202), .A2(n118619), .B1(n120196), .B2(n119247), 
        .ZN(n114905) );
  OAI221_X1 U85678 ( .B1(n114154), .B2(n120214), .C1(n98656), .C2(n120208), 
        .A(n114877), .ZN(n114873) );
  AOI22_X1 U85679 ( .A1(n120202), .A2(n118620), .B1(n120196), .B2(n119248), 
        .ZN(n114877) );
  OAI221_X1 U85680 ( .B1(n114153), .B2(n120214), .C1(n98655), .C2(n120208), 
        .A(n114849), .ZN(n114845) );
  AOI22_X1 U85681 ( .A1(n120202), .A2(n118621), .B1(n120196), .B2(n119249), 
        .ZN(n114849) );
  OAI221_X1 U85682 ( .B1(n114152), .B2(n120214), .C1(n98654), .C2(n120208), 
        .A(n114821), .ZN(n114817) );
  AOI22_X1 U85683 ( .A1(n120202), .A2(n118622), .B1(n120196), .B2(n119250), 
        .ZN(n114821) );
  OAI221_X1 U85684 ( .B1(n114151), .B2(n120214), .C1(n98653), .C2(n120208), 
        .A(n114793), .ZN(n114789) );
  AOI22_X1 U85685 ( .A1(n120202), .A2(n118623), .B1(n120196), .B2(n119251), 
        .ZN(n114793) );
  OAI221_X1 U85686 ( .B1(n114198), .B2(n120211), .C1(n98700), .C2(n120205), 
        .A(n116109), .ZN(n116105) );
  AOI22_X1 U85687 ( .A1(n120199), .A2(n118624), .B1(n120193), .B2(n119252), 
        .ZN(n116109) );
  OAI221_X1 U85688 ( .B1(n114197), .B2(n120211), .C1(n98699), .C2(n120205), 
        .A(n116081), .ZN(n116077) );
  AOI22_X1 U85689 ( .A1(n120199), .A2(n118625), .B1(n120193), .B2(n119253), 
        .ZN(n116081) );
  OAI221_X1 U85690 ( .B1(n114196), .B2(n120211), .C1(n98698), .C2(n120205), 
        .A(n116053), .ZN(n116049) );
  AOI22_X1 U85691 ( .A1(n120199), .A2(n118626), .B1(n120193), .B2(n119254), 
        .ZN(n116053) );
  OAI221_X1 U85692 ( .B1(n114195), .B2(n120211), .C1(n98697), .C2(n120205), 
        .A(n116025), .ZN(n116021) );
  AOI22_X1 U85693 ( .A1(n120199), .A2(n118627), .B1(n120193), .B2(n119255), 
        .ZN(n116025) );
  OAI221_X1 U85694 ( .B1(n114194), .B2(n120211), .C1(n98696), .C2(n120205), 
        .A(n115997), .ZN(n115993) );
  AOI22_X1 U85695 ( .A1(n120199), .A2(n118628), .B1(n120193), .B2(n119256), 
        .ZN(n115997) );
  OAI221_X1 U85696 ( .B1(n114193), .B2(n120211), .C1(n98695), .C2(n120205), 
        .A(n115969), .ZN(n115965) );
  AOI22_X1 U85697 ( .A1(n120199), .A2(n118629), .B1(n120193), .B2(n119257), 
        .ZN(n115969) );
  OAI221_X1 U85698 ( .B1(n114192), .B2(n120211), .C1(n98694), .C2(n120205), 
        .A(n115941), .ZN(n115937) );
  AOI22_X1 U85699 ( .A1(n120199), .A2(n118630), .B1(n120193), .B2(n119258), 
        .ZN(n115941) );
  OAI221_X1 U85700 ( .B1(n114191), .B2(n120211), .C1(n98693), .C2(n120205), 
        .A(n115913), .ZN(n115909) );
  AOI22_X1 U85701 ( .A1(n120199), .A2(n118631), .B1(n120193), .B2(n119259), 
        .ZN(n115913) );
  OAI221_X1 U85702 ( .B1(n114190), .B2(n120211), .C1(n98692), .C2(n120205), 
        .A(n115885), .ZN(n115881) );
  AOI22_X1 U85703 ( .A1(n120199), .A2(n118632), .B1(n120193), .B2(n119260), 
        .ZN(n115885) );
  OAI221_X1 U85704 ( .B1(n114189), .B2(n120211), .C1(n98691), .C2(n120205), 
        .A(n115857), .ZN(n115853) );
  AOI22_X1 U85705 ( .A1(n120199), .A2(n118633), .B1(n120193), .B2(n119261), 
        .ZN(n115857) );
  OAI221_X1 U85706 ( .B1(n114188), .B2(n120211), .C1(n98690), .C2(n120205), 
        .A(n115829), .ZN(n115825) );
  AOI22_X1 U85707 ( .A1(n120199), .A2(n118634), .B1(n120193), .B2(n119262), 
        .ZN(n115829) );
  OAI221_X1 U85708 ( .B1(n114187), .B2(n120211), .C1(n98689), .C2(n120205), 
        .A(n115801), .ZN(n115797) );
  AOI22_X1 U85709 ( .A1(n120199), .A2(n118635), .B1(n120193), .B2(n119263), 
        .ZN(n115801) );
  OAI221_X1 U85710 ( .B1(n114186), .B2(n120212), .C1(n98688), .C2(n120206), 
        .A(n115773), .ZN(n115769) );
  AOI22_X1 U85711 ( .A1(n120200), .A2(n118636), .B1(n120194), .B2(n119264), 
        .ZN(n115773) );
  OAI221_X1 U85712 ( .B1(n114185), .B2(n120212), .C1(n98687), .C2(n120206), 
        .A(n115745), .ZN(n115741) );
  AOI22_X1 U85713 ( .A1(n120200), .A2(n118637), .B1(n120194), .B2(n119265), 
        .ZN(n115745) );
  OAI221_X1 U85714 ( .B1(n114184), .B2(n120212), .C1(n98686), .C2(n120206), 
        .A(n115717), .ZN(n115713) );
  AOI22_X1 U85715 ( .A1(n120200), .A2(n118638), .B1(n120194), .B2(n119266), 
        .ZN(n115717) );
  OAI221_X1 U85716 ( .B1(n114183), .B2(n120212), .C1(n98685), .C2(n120206), 
        .A(n115689), .ZN(n115685) );
  AOI22_X1 U85717 ( .A1(n120200), .A2(n118639), .B1(n120194), .B2(n119267), 
        .ZN(n115689) );
  OAI221_X1 U85718 ( .B1(n114182), .B2(n120212), .C1(n98684), .C2(n120206), 
        .A(n115661), .ZN(n115657) );
  AOI22_X1 U85719 ( .A1(n120200), .A2(n118640), .B1(n120194), .B2(n119268), 
        .ZN(n115661) );
  OAI221_X1 U85720 ( .B1(n114181), .B2(n120212), .C1(n98683), .C2(n120206), 
        .A(n115633), .ZN(n115629) );
  AOI22_X1 U85721 ( .A1(n120200), .A2(n118641), .B1(n120194), .B2(n119269), 
        .ZN(n115633) );
  OAI221_X1 U85722 ( .B1(n114180), .B2(n120212), .C1(n98682), .C2(n120206), 
        .A(n115605), .ZN(n115601) );
  AOI22_X1 U85723 ( .A1(n120200), .A2(n118642), .B1(n120194), .B2(n119270), 
        .ZN(n115605) );
  OAI221_X1 U85724 ( .B1(n114179), .B2(n120212), .C1(n98681), .C2(n120206), 
        .A(n115577), .ZN(n115573) );
  AOI22_X1 U85725 ( .A1(n120200), .A2(n118643), .B1(n120194), .B2(n119271), 
        .ZN(n115577) );
  OAI221_X1 U85726 ( .B1(n114178), .B2(n120212), .C1(n98680), .C2(n120206), 
        .A(n115549), .ZN(n115545) );
  AOI22_X1 U85727 ( .A1(n120200), .A2(n118644), .B1(n120194), .B2(n119272), 
        .ZN(n115549) );
  OAI221_X1 U85728 ( .B1(n114177), .B2(n120212), .C1(n98679), .C2(n120206), 
        .A(n115521), .ZN(n115517) );
  AOI22_X1 U85729 ( .A1(n120200), .A2(n118645), .B1(n120194), .B2(n119273), 
        .ZN(n115521) );
  OAI221_X1 U85730 ( .B1(n114176), .B2(n120212), .C1(n98678), .C2(n120206), 
        .A(n115493), .ZN(n115489) );
  AOI22_X1 U85731 ( .A1(n120200), .A2(n118646), .B1(n120194), .B2(n119274), 
        .ZN(n115493) );
  OAI221_X1 U85732 ( .B1(n114175), .B2(n120212), .C1(n98677), .C2(n120206), 
        .A(n115465), .ZN(n115461) );
  AOI22_X1 U85733 ( .A1(n120200), .A2(n118647), .B1(n120194), .B2(n119275), 
        .ZN(n115465) );
  OAI221_X1 U85734 ( .B1(n114174), .B2(n120213), .C1(n98676), .C2(n120207), 
        .A(n115437), .ZN(n115433) );
  AOI22_X1 U85735 ( .A1(n120201), .A2(n118648), .B1(n120195), .B2(n119276), 
        .ZN(n115437) );
  OAI221_X1 U85736 ( .B1(n114173), .B2(n120213), .C1(n98675), .C2(n120207), 
        .A(n115409), .ZN(n115405) );
  AOI22_X1 U85737 ( .A1(n120201), .A2(n118649), .B1(n120195), .B2(n119277), 
        .ZN(n115409) );
  OAI221_X1 U85738 ( .B1(n114172), .B2(n120213), .C1(n98674), .C2(n120207), 
        .A(n115381), .ZN(n115377) );
  AOI22_X1 U85739 ( .A1(n120201), .A2(n118650), .B1(n120195), .B2(n119278), 
        .ZN(n115381) );
  OAI221_X1 U85740 ( .B1(n114171), .B2(n120213), .C1(n98673), .C2(n120207), 
        .A(n115353), .ZN(n115349) );
  AOI22_X1 U85741 ( .A1(n120201), .A2(n118651), .B1(n120195), .B2(n119279), 
        .ZN(n115353) );
  OAI221_X1 U85742 ( .B1(n114170), .B2(n120213), .C1(n98672), .C2(n120207), 
        .A(n115325), .ZN(n115321) );
  AOI22_X1 U85743 ( .A1(n120201), .A2(n118652), .B1(n120195), .B2(n119280), 
        .ZN(n115325) );
  OAI221_X1 U85744 ( .B1(n114169), .B2(n120213), .C1(n98671), .C2(n120207), 
        .A(n115297), .ZN(n115293) );
  AOI22_X1 U85745 ( .A1(n120201), .A2(n118653), .B1(n120195), .B2(n119281), 
        .ZN(n115297) );
  OAI221_X1 U85746 ( .B1(n114168), .B2(n120213), .C1(n98670), .C2(n120207), 
        .A(n115269), .ZN(n115265) );
  AOI22_X1 U85747 ( .A1(n120201), .A2(n118654), .B1(n120195), .B2(n119282), 
        .ZN(n115269) );
  OAI221_X1 U85748 ( .B1(n114167), .B2(n120213), .C1(n98669), .C2(n120207), 
        .A(n115241), .ZN(n115237) );
  AOI22_X1 U85749 ( .A1(n120201), .A2(n118655), .B1(n120195), .B2(n119283), 
        .ZN(n115241) );
  OAI221_X1 U85750 ( .B1(n114166), .B2(n120213), .C1(n98668), .C2(n120207), 
        .A(n115213), .ZN(n115209) );
  AOI22_X1 U85751 ( .A1(n120201), .A2(n118656), .B1(n120195), .B2(n119284), 
        .ZN(n115213) );
  OAI221_X1 U85752 ( .B1(n114165), .B2(n120213), .C1(n98667), .C2(n120207), 
        .A(n115185), .ZN(n115181) );
  AOI22_X1 U85753 ( .A1(n120201), .A2(n118657), .B1(n120195), .B2(n119285), 
        .ZN(n115185) );
  OAI221_X1 U85754 ( .B1(n114210), .B2(n120210), .C1(n98712), .C2(n120204), 
        .A(n116449), .ZN(n116441) );
  AOI22_X1 U85755 ( .A1(n120198), .A2(n118658), .B1(n120192), .B2(n119286), 
        .ZN(n116449) );
  OAI221_X1 U85756 ( .B1(n114209), .B2(n120210), .C1(n98711), .C2(n120204), 
        .A(n116417), .ZN(n116413) );
  AOI22_X1 U85757 ( .A1(n120198), .A2(n118659), .B1(n120192), .B2(n119287), 
        .ZN(n116417) );
  OAI221_X1 U85758 ( .B1(n114208), .B2(n120210), .C1(n98710), .C2(n120204), 
        .A(n116389), .ZN(n116385) );
  AOI22_X1 U85759 ( .A1(n120198), .A2(n118660), .B1(n120192), .B2(n119288), 
        .ZN(n116389) );
  OAI221_X1 U85760 ( .B1(n114207), .B2(n120210), .C1(n98709), .C2(n120204), 
        .A(n116361), .ZN(n116357) );
  AOI22_X1 U85761 ( .A1(n120198), .A2(n118661), .B1(n120192), .B2(n119289), 
        .ZN(n116361) );
  OAI221_X1 U85762 ( .B1(n114206), .B2(n120210), .C1(n98708), .C2(n120204), 
        .A(n116333), .ZN(n116329) );
  AOI22_X1 U85763 ( .A1(n120198), .A2(n118662), .B1(n120192), .B2(n119290), 
        .ZN(n116333) );
  OAI221_X1 U85764 ( .B1(n114205), .B2(n120210), .C1(n98707), .C2(n120204), 
        .A(n116305), .ZN(n116301) );
  AOI22_X1 U85765 ( .A1(n120198), .A2(n118663), .B1(n120192), .B2(n119291), 
        .ZN(n116305) );
  OAI221_X1 U85766 ( .B1(n114204), .B2(n120210), .C1(n98706), .C2(n120204), 
        .A(n116277), .ZN(n116273) );
  AOI22_X1 U85767 ( .A1(n120198), .A2(n118664), .B1(n120192), .B2(n119292), 
        .ZN(n116277) );
  OAI221_X1 U85768 ( .B1(n114203), .B2(n120210), .C1(n98705), .C2(n120204), 
        .A(n116249), .ZN(n116245) );
  AOI22_X1 U85769 ( .A1(n120198), .A2(n118665), .B1(n120192), .B2(n119293), 
        .ZN(n116249) );
  OAI221_X1 U85770 ( .B1(n114202), .B2(n120210), .C1(n98704), .C2(n120204), 
        .A(n116221), .ZN(n116217) );
  AOI22_X1 U85771 ( .A1(n120198), .A2(n118666), .B1(n120192), .B2(n119294), 
        .ZN(n116221) );
  OAI221_X1 U85772 ( .B1(n114201), .B2(n120210), .C1(n98703), .C2(n120204), 
        .A(n116193), .ZN(n116189) );
  AOI22_X1 U85773 ( .A1(n120198), .A2(n118667), .B1(n120192), .B2(n119295), 
        .ZN(n116193) );
  OAI221_X1 U85774 ( .B1(n114200), .B2(n120210), .C1(n98702), .C2(n120204), 
        .A(n116165), .ZN(n116161) );
  AOI22_X1 U85775 ( .A1(n120198), .A2(n118668), .B1(n120192), .B2(n119296), 
        .ZN(n116165) );
  OAI221_X1 U85776 ( .B1(n114199), .B2(n120210), .C1(n98701), .C2(n120204), 
        .A(n116137), .ZN(n116133) );
  AOI22_X1 U85777 ( .A1(n120198), .A2(n118669), .B1(n120192), .B2(n119297), 
        .ZN(n116137) );
  OAI221_X1 U85778 ( .B1(n114127), .B2(n120191), .C1(n114382), .C2(n120185), 
        .A(n114769), .ZN(n114762) );
  AOI22_X1 U85779 ( .A1(n120179), .A2(n117974), .B1(n120173), .B2(n119110), 
        .ZN(n114769) );
  OAI221_X1 U85780 ( .B1(n114126), .B2(n120191), .C1(n114381), .C2(n120185), 
        .A(n114743), .ZN(n114736) );
  AOI22_X1 U85781 ( .A1(n120179), .A2(n117975), .B1(n120173), .B2(n119111), 
        .ZN(n114743) );
  OAI221_X1 U85782 ( .B1(n114125), .B2(n120191), .C1(n114380), .C2(n120185), 
        .A(n114717), .ZN(n114710) );
  AOI22_X1 U85783 ( .A1(n120179), .A2(n117976), .B1(n120173), .B2(n119112), 
        .ZN(n114717) );
  OAI221_X1 U85784 ( .B1(n114123), .B2(n120191), .C1(n114378), .C2(n120185), 
        .A(n114668), .ZN(n114651) );
  AOI22_X1 U85785 ( .A1(n120179), .A2(n117977), .B1(n120173), .B2(n119113), 
        .ZN(n114668) );
  OAI221_X1 U85786 ( .B1(n114514), .B2(n119993), .C1(n114150), .C2(n119987), 
        .A(n116587), .ZN(n116580) );
  AOI22_X1 U85787 ( .A1(n119981), .A2(n111041), .B1(n119975), .B2(n117993), 
        .ZN(n116587) );
  OAI221_X1 U85788 ( .B1(n114513), .B2(n119993), .C1(n114149), .C2(n119987), 
        .A(n116566), .ZN(n116559) );
  AOI22_X1 U85789 ( .A1(n119981), .A2(n111042), .B1(n119975), .B2(n117994), 
        .ZN(n116566) );
  OAI221_X1 U85790 ( .B1(n114512), .B2(n119993), .C1(n114148), .C2(n119987), 
        .A(n116545), .ZN(n116538) );
  AOI22_X1 U85791 ( .A1(n119981), .A2(n111043), .B1(n119975), .B2(n117995), 
        .ZN(n116545) );
  OAI221_X1 U85792 ( .B1(n114510), .B2(n119993), .C1(n114146), .C2(n119987), 
        .A(n116501), .ZN(n116484) );
  AOI22_X1 U85793 ( .A1(n119981), .A2(n111044), .B1(n119975), .B2(n117996), 
        .ZN(n116501) );
  OAI221_X1 U85794 ( .B1(n114514), .B2(n120167), .C1(n114448), .C2(n120161), 
        .A(n114771), .ZN(n114761) );
  AOI22_X1 U85795 ( .A1(n120155), .A2(n111045), .B1(n120149), .B2(n119046), 
        .ZN(n114771) );
  OAI221_X1 U85796 ( .B1(n114513), .B2(n120167), .C1(n114447), .C2(n120161), 
        .A(n114745), .ZN(n114735) );
  AOI22_X1 U85797 ( .A1(n120155), .A2(n111046), .B1(n120149), .B2(n119047), 
        .ZN(n114745) );
  OAI221_X1 U85798 ( .B1(n114512), .B2(n120167), .C1(n114446), .C2(n120161), 
        .A(n114719), .ZN(n114709) );
  AOI22_X1 U85799 ( .A1(n120155), .A2(n111047), .B1(n120149), .B2(n119048), 
        .ZN(n114719) );
  OAI221_X1 U85800 ( .B1(n114510), .B2(n120167), .C1(n114444), .C2(n120161), 
        .A(n114674), .ZN(n114650) );
  AOI22_X1 U85801 ( .A1(n120155), .A2(n111048), .B1(n120149), .B2(n119049), 
        .ZN(n114674) );
  OAI221_X1 U85802 ( .B1(n99183), .B2(n119969), .C1(n113985), .C2(n119963), 
        .A(n116588), .ZN(n116579) );
  AOI22_X1 U85803 ( .A1(n119957), .A2(n117981), .B1(n119951), .B2(n117974), 
        .ZN(n116588) );
  OAI221_X1 U85804 ( .B1(n99182), .B2(n119969), .C1(n113984), .C2(n119963), 
        .A(n116567), .ZN(n116558) );
  AOI22_X1 U85805 ( .A1(n119957), .A2(n117982), .B1(n119951), .B2(n117975), 
        .ZN(n116567) );
  OAI221_X1 U85806 ( .B1(n99181), .B2(n119969), .C1(n113983), .C2(n119963), 
        .A(n116546), .ZN(n116537) );
  AOI22_X1 U85807 ( .A1(n119957), .A2(n117983), .B1(n119951), .B2(n117976), 
        .ZN(n116546) );
  OAI221_X1 U85808 ( .B1(n99179), .B2(n119969), .C1(n113981), .C2(n119963), 
        .A(n116506), .ZN(n116483) );
  AOI22_X1 U85809 ( .A1(n119957), .A2(n117984), .B1(n119951), .B2(n117977), 
        .ZN(n116506) );
  OAI22_X1 U85810 ( .A1(n99051), .A2(n120143), .B1(n89500), .B2(n120137), .ZN(
        n114776) );
  OAI22_X1 U85811 ( .A1(n99050), .A2(n120143), .B1(n89498), .B2(n120137), .ZN(
        n114750) );
  OAI22_X1 U85812 ( .A1(n99049), .A2(n120143), .B1(n89496), .B2(n120137), .ZN(
        n114724) );
  OAI22_X1 U85813 ( .A1(n99047), .A2(n120143), .B1(n89493), .B2(n120137), .ZN(
        n114681) );
  OAI22_X1 U85814 ( .A1(n99720), .A2(n119945), .B1(n89500), .B2(n119939), .ZN(
        n116592) );
  OAI22_X1 U85815 ( .A1(n99719), .A2(n119945), .B1(n89498), .B2(n119939), .ZN(
        n116571) );
  OAI22_X1 U85816 ( .A1(n99718), .A2(n119945), .B1(n89496), .B2(n119939), .ZN(
        n116550) );
  OAI22_X1 U85817 ( .A1(n99716), .A2(n119945), .B1(n89493), .B2(n119939), .ZN(
        n116512) );
  OAI22_X1 U85818 ( .A1(n90310), .A2(n120131), .B1(n114239), .B2(n120125), 
        .ZN(n114775) );
  OAI22_X1 U85819 ( .A1(n90309), .A2(n120131), .B1(n114238), .B2(n120125), 
        .ZN(n114749) );
  OAI22_X1 U85820 ( .A1(n90308), .A2(n120131), .B1(n114237), .B2(n120125), 
        .ZN(n114723) );
  OAI22_X1 U85821 ( .A1(n90306), .A2(n120131), .B1(n114235), .B2(n120125), 
        .ZN(n114680) );
  OAI22_X1 U85822 ( .A1(n90715), .A2(n119933), .B1(n99051), .B2(n119927), .ZN(
        n116591) );
  OAI22_X1 U85823 ( .A1(n90714), .A2(n119933), .B1(n99050), .B2(n119927), .ZN(
        n116570) );
  OAI22_X1 U85824 ( .A1(n90713), .A2(n119933), .B1(n99049), .B2(n119927), .ZN(
        n116549) );
  OAI22_X1 U85825 ( .A1(n90711), .A2(n119933), .B1(n99047), .B2(n119927), .ZN(
        n116511) );
  OAI22_X1 U85826 ( .A1(n89969), .A2(n119879), .B1(n99450), .B2(n119873), .ZN(
        n116594) );
  OAI22_X1 U85827 ( .A1(n89968), .A2(n119879), .B1(n99449), .B2(n119873), .ZN(
        n116573) );
  OAI22_X1 U85828 ( .A1(n89967), .A2(n119879), .B1(n99448), .B2(n119873), .ZN(
        n116552) );
  OAI22_X1 U85829 ( .A1(n89965), .A2(n119879), .B1(n99446), .B2(n119873), .ZN(
        n116525) );
  OAI22_X1 U85830 ( .A1(n90516), .A2(n120119), .B1(n90035), .B2(n120113), .ZN(
        n114774) );
  OAI22_X1 U85831 ( .A1(n90515), .A2(n120119), .B1(n90034), .B2(n120113), .ZN(
        n114748) );
  OAI22_X1 U85832 ( .A1(n90514), .A2(n120119), .B1(n90033), .B2(n120113), .ZN(
        n114722) );
  OAI22_X1 U85833 ( .A1(n90512), .A2(n120119), .B1(n90031), .B2(n120113), .ZN(
        n114679) );
  OAI22_X1 U85834 ( .A1(n98718), .A2(n119921), .B1(n90377), .B2(n119915), .ZN(
        n116590) );
  OAI22_X1 U85835 ( .A1(n98717), .A2(n119921), .B1(n90376), .B2(n119915), .ZN(
        n116569) );
  OAI22_X1 U85836 ( .A1(n98716), .A2(n119921), .B1(n90375), .B2(n119915), .ZN(
        n116548) );
  OAI22_X1 U85837 ( .A1(n98714), .A2(n119921), .B1(n90373), .B2(n119915), .ZN(
        n116510) );
  OAI22_X1 U85838 ( .A1(n90764), .A2(n119928), .B1(n99100), .B2(n119922), .ZN(
        n117711) );
  OAI22_X1 U85839 ( .A1(n90763), .A2(n119929), .B1(n99099), .B2(n119923), .ZN(
        n117689) );
  OAI22_X1 U85840 ( .A1(n90762), .A2(n119929), .B1(n99098), .B2(n119923), .ZN(
        n117667) );
  OAI22_X1 U85841 ( .A1(n90761), .A2(n119929), .B1(n99097), .B2(n119923), .ZN(
        n117645) );
  OAI22_X1 U85842 ( .A1(n90760), .A2(n119929), .B1(n99096), .B2(n119923), .ZN(
        n117623) );
  OAI22_X1 U85843 ( .A1(n90759), .A2(n119929), .B1(n99095), .B2(n119923), .ZN(
        n117601) );
  OAI22_X1 U85844 ( .A1(n90758), .A2(n119929), .B1(n99094), .B2(n119923), .ZN(
        n117579) );
  OAI22_X1 U85845 ( .A1(n90757), .A2(n119929), .B1(n99093), .B2(n119923), .ZN(
        n117557) );
  OAI22_X1 U85846 ( .A1(n90756), .A2(n119929), .B1(n99092), .B2(n119923), .ZN(
        n117534) );
  OAI22_X1 U85847 ( .A1(n90755), .A2(n119929), .B1(n99091), .B2(n119923), .ZN(
        n117511) );
  OAI22_X1 U85848 ( .A1(n90754), .A2(n119929), .B1(n99090), .B2(n119923), .ZN(
        n117488) );
  OAI22_X1 U85849 ( .A1(n90753), .A2(n119929), .B1(n99089), .B2(n119923), .ZN(
        n117465) );
  OAI22_X1 U85850 ( .A1(n90752), .A2(n119929), .B1(n99088), .B2(n119923), .ZN(
        n117442) );
  OAI22_X1 U85851 ( .A1(n90751), .A2(n119930), .B1(n99087), .B2(n119924), .ZN(
        n117419) );
  OAI22_X1 U85852 ( .A1(n90750), .A2(n119930), .B1(n99086), .B2(n119924), .ZN(
        n117396) );
  OAI22_X1 U85853 ( .A1(n90749), .A2(n119930), .B1(n99085), .B2(n119924), .ZN(
        n117373) );
  OAI22_X1 U85854 ( .A1(n90748), .A2(n119930), .B1(n99084), .B2(n119924), .ZN(
        n117350) );
  OAI22_X1 U85855 ( .A1(n90747), .A2(n119930), .B1(n99083), .B2(n119924), .ZN(
        n117327) );
  OAI22_X1 U85856 ( .A1(n90746), .A2(n119930), .B1(n99082), .B2(n119924), .ZN(
        n117304) );
  OAI22_X1 U85857 ( .A1(n90745), .A2(n119930), .B1(n99081), .B2(n119924), .ZN(
        n117281) );
  OAI22_X1 U85858 ( .A1(n90744), .A2(n119930), .B1(n99080), .B2(n119924), .ZN(
        n117258) );
  OAI22_X1 U85859 ( .A1(n90743), .A2(n119930), .B1(n99079), .B2(n119924), .ZN(
        n117235) );
  OAI22_X1 U85860 ( .A1(n90742), .A2(n119930), .B1(n99078), .B2(n119924), .ZN(
        n117212) );
  OAI22_X1 U85861 ( .A1(n90741), .A2(n119930), .B1(n99077), .B2(n119924), .ZN(
        n117189) );
  OAI22_X1 U85862 ( .A1(n90740), .A2(n119930), .B1(n99076), .B2(n119924), .ZN(
        n117166) );
  OAI22_X1 U85863 ( .A1(n90739), .A2(n119931), .B1(n99075), .B2(n119925), .ZN(
        n117143) );
  OAI22_X1 U85864 ( .A1(n90738), .A2(n119931), .B1(n99074), .B2(n119925), .ZN(
        n117120) );
  OAI22_X1 U85865 ( .A1(n90737), .A2(n119931), .B1(n99073), .B2(n119925), .ZN(
        n117097) );
  OAI22_X1 U85866 ( .A1(n90736), .A2(n119931), .B1(n99072), .B2(n119925), .ZN(
        n117074) );
  OAI22_X1 U85867 ( .A1(n90735), .A2(n119931), .B1(n99071), .B2(n119925), .ZN(
        n117051) );
  OAI22_X1 U85868 ( .A1(n90734), .A2(n119931), .B1(n99070), .B2(n119925), .ZN(
        n117028) );
  OAI22_X1 U85869 ( .A1(n90733), .A2(n119931), .B1(n99069), .B2(n119925), .ZN(
        n117005) );
  OAI22_X1 U85870 ( .A1(n90732), .A2(n119931), .B1(n99068), .B2(n119925), .ZN(
        n116982) );
  OAI22_X1 U85871 ( .A1(n90731), .A2(n119931), .B1(n99067), .B2(n119925), .ZN(
        n116959) );
  OAI22_X1 U85872 ( .A1(n90730), .A2(n119931), .B1(n99066), .B2(n119925), .ZN(
        n116936) );
  OAI22_X1 U85873 ( .A1(n90729), .A2(n119931), .B1(n99065), .B2(n119925), .ZN(
        n116913) );
  OAI22_X1 U85874 ( .A1(n90728), .A2(n119931), .B1(n99064), .B2(n119925), .ZN(
        n116890) );
  OAI22_X1 U85875 ( .A1(n90727), .A2(n119932), .B1(n99063), .B2(n119926), .ZN(
        n116867) );
  OAI22_X1 U85876 ( .A1(n90726), .A2(n119932), .B1(n99062), .B2(n119926), .ZN(
        n116844) );
  OAI22_X1 U85877 ( .A1(n90725), .A2(n119932), .B1(n99061), .B2(n119926), .ZN(
        n116821) );
  OAI22_X1 U85878 ( .A1(n90724), .A2(n119932), .B1(n99060), .B2(n119926), .ZN(
        n116798) );
  OAI22_X1 U85879 ( .A1(n90723), .A2(n119932), .B1(n99059), .B2(n119926), .ZN(
        n116775) );
  OAI22_X1 U85880 ( .A1(n90722), .A2(n119932), .B1(n99058), .B2(n119926), .ZN(
        n116752) );
  OAI22_X1 U85881 ( .A1(n90721), .A2(n119932), .B1(n99057), .B2(n119926), .ZN(
        n116729) );
  OAI22_X1 U85882 ( .A1(n90720), .A2(n119932), .B1(n99056), .B2(n119926), .ZN(
        n116706) );
  OAI22_X1 U85883 ( .A1(n90719), .A2(n119932), .B1(n99055), .B2(n119926), .ZN(
        n116683) );
  OAI22_X1 U85884 ( .A1(n90718), .A2(n119932), .B1(n99054), .B2(n119926), .ZN(
        n116660) );
  OAI22_X1 U85885 ( .A1(n90717), .A2(n119932), .B1(n99053), .B2(n119926), .ZN(
        n116637) );
  OAI22_X1 U85886 ( .A1(n90716), .A2(n119932), .B1(n99052), .B2(n119926), .ZN(
        n116614) );
  OAI22_X1 U85887 ( .A1(n90768), .A2(n119928), .B1(n99104), .B2(n119922), .ZN(
        n117799) );
  OAI22_X1 U85888 ( .A1(n90767), .A2(n119928), .B1(n99103), .B2(n119922), .ZN(
        n117777) );
  OAI22_X1 U85889 ( .A1(n90766), .A2(n119928), .B1(n99102), .B2(n119922), .ZN(
        n117755) );
  OAI22_X1 U85890 ( .A1(n90765), .A2(n119928), .B1(n99101), .B2(n119922), .ZN(
        n117733) );
  OAI22_X1 U85891 ( .A1(n90775), .A2(n119928), .B1(n99111), .B2(n119922), .ZN(
        n117965) );
  OAI22_X1 U85892 ( .A1(n90774), .A2(n119928), .B1(n99110), .B2(n119922), .ZN(
        n117931) );
  OAI22_X1 U85893 ( .A1(n90773), .A2(n119928), .B1(n99109), .B2(n119922), .ZN(
        n117909) );
  OAI22_X1 U85894 ( .A1(n90772), .A2(n119928), .B1(n99108), .B2(n119922), .ZN(
        n117887) );
  OAI22_X1 U85895 ( .A1(n90771), .A2(n119928), .B1(n99107), .B2(n119922), .ZN(
        n117865) );
  OAI22_X1 U85896 ( .A1(n90770), .A2(n119928), .B1(n99106), .B2(n119922), .ZN(
        n117843) );
  OAI22_X1 U85897 ( .A1(n90769), .A2(n119928), .B1(n99105), .B2(n119922), .ZN(
        n117821) );
  OAI22_X1 U85898 ( .A1(n98701), .A2(n119850), .B1(n99633), .B2(n119844), .ZN(
        n117714) );
  OAI22_X1 U85899 ( .A1(n98700), .A2(n119851), .B1(n99632), .B2(n119845), .ZN(
        n117692) );
  OAI22_X1 U85900 ( .A1(n98699), .A2(n119851), .B1(n99631), .B2(n119845), .ZN(
        n117670) );
  OAI22_X1 U85901 ( .A1(n98698), .A2(n119851), .B1(n99630), .B2(n119845), .ZN(
        n117648) );
  OAI22_X1 U85902 ( .A1(n98697), .A2(n119851), .B1(n99629), .B2(n119845), .ZN(
        n117626) );
  OAI22_X1 U85903 ( .A1(n98696), .A2(n119851), .B1(n99628), .B2(n119845), .ZN(
        n117604) );
  OAI22_X1 U85904 ( .A1(n98695), .A2(n119851), .B1(n99627), .B2(n119845), .ZN(
        n117582) );
  OAI22_X1 U85905 ( .A1(n98694), .A2(n119851), .B1(n99626), .B2(n119845), .ZN(
        n117560) );
  OAI22_X1 U85906 ( .A1(n98693), .A2(n119851), .B1(n99625), .B2(n119845), .ZN(
        n117538) );
  OAI22_X1 U85907 ( .A1(n98692), .A2(n119851), .B1(n99624), .B2(n119845), .ZN(
        n117515) );
  OAI22_X1 U85908 ( .A1(n98691), .A2(n119851), .B1(n99623), .B2(n119845), .ZN(
        n117492) );
  OAI22_X1 U85909 ( .A1(n98690), .A2(n119851), .B1(n99622), .B2(n119845), .ZN(
        n117469) );
  OAI22_X1 U85910 ( .A1(n98689), .A2(n119851), .B1(n99621), .B2(n119845), .ZN(
        n117446) );
  OAI22_X1 U85911 ( .A1(n98688), .A2(n119852), .B1(n99620), .B2(n119846), .ZN(
        n117423) );
  OAI22_X1 U85912 ( .A1(n98687), .A2(n119852), .B1(n99619), .B2(n119846), .ZN(
        n117400) );
  OAI22_X1 U85913 ( .A1(n98686), .A2(n119852), .B1(n99618), .B2(n119846), .ZN(
        n117377) );
  OAI22_X1 U85914 ( .A1(n98685), .A2(n119852), .B1(n99617), .B2(n119846), .ZN(
        n117354) );
  OAI22_X1 U85915 ( .A1(n98684), .A2(n119852), .B1(n99616), .B2(n119846), .ZN(
        n117331) );
  OAI22_X1 U85916 ( .A1(n98683), .A2(n119852), .B1(n99615), .B2(n119846), .ZN(
        n117308) );
  OAI22_X1 U85917 ( .A1(n98682), .A2(n119852), .B1(n99614), .B2(n119846), .ZN(
        n117285) );
  OAI22_X1 U85918 ( .A1(n98681), .A2(n119852), .B1(n99613), .B2(n119846), .ZN(
        n117262) );
  OAI22_X1 U85919 ( .A1(n98680), .A2(n119852), .B1(n99612), .B2(n119846), .ZN(
        n117239) );
  OAI22_X1 U85920 ( .A1(n98679), .A2(n119852), .B1(n99611), .B2(n119846), .ZN(
        n117216) );
  OAI22_X1 U85921 ( .A1(n98678), .A2(n119852), .B1(n99610), .B2(n119846), .ZN(
        n117193) );
  OAI22_X1 U85922 ( .A1(n98677), .A2(n119852), .B1(n99609), .B2(n119846), .ZN(
        n117170) );
  OAI22_X1 U85923 ( .A1(n98676), .A2(n119853), .B1(n99608), .B2(n119847), .ZN(
        n117147) );
  OAI22_X1 U85924 ( .A1(n98675), .A2(n119853), .B1(n99607), .B2(n119847), .ZN(
        n117124) );
  OAI22_X1 U85925 ( .A1(n98674), .A2(n119853), .B1(n99606), .B2(n119847), .ZN(
        n117101) );
  OAI22_X1 U85926 ( .A1(n98673), .A2(n119853), .B1(n99605), .B2(n119847), .ZN(
        n117078) );
  OAI22_X1 U85927 ( .A1(n98672), .A2(n119853), .B1(n99604), .B2(n119847), .ZN(
        n117055) );
  OAI22_X1 U85928 ( .A1(n98671), .A2(n119853), .B1(n99603), .B2(n119847), .ZN(
        n117032) );
  OAI22_X1 U85929 ( .A1(n98670), .A2(n119853), .B1(n99602), .B2(n119847), .ZN(
        n117009) );
  OAI22_X1 U85930 ( .A1(n98669), .A2(n119853), .B1(n99601), .B2(n119847), .ZN(
        n116986) );
  OAI22_X1 U85931 ( .A1(n98668), .A2(n119853), .B1(n99600), .B2(n119847), .ZN(
        n116963) );
  OAI22_X1 U85932 ( .A1(n98667), .A2(n119853), .B1(n99599), .B2(n119847), .ZN(
        n116940) );
  OAI22_X1 U85933 ( .A1(n98666), .A2(n119853), .B1(n99598), .B2(n119847), .ZN(
        n116917) );
  OAI22_X1 U85934 ( .A1(n98665), .A2(n119853), .B1(n99597), .B2(n119847), .ZN(
        n116894) );
  OAI22_X1 U85935 ( .A1(n98664), .A2(n119854), .B1(n99596), .B2(n119848), .ZN(
        n116871) );
  OAI22_X1 U85936 ( .A1(n98663), .A2(n119854), .B1(n99595), .B2(n119848), .ZN(
        n116848) );
  OAI22_X1 U85937 ( .A1(n98662), .A2(n119854), .B1(n99594), .B2(n119848), .ZN(
        n116825) );
  OAI22_X1 U85938 ( .A1(n98661), .A2(n119854), .B1(n99593), .B2(n119848), .ZN(
        n116802) );
  OAI22_X1 U85939 ( .A1(n98660), .A2(n119854), .B1(n99592), .B2(n119848), .ZN(
        n116779) );
  OAI22_X1 U85940 ( .A1(n98659), .A2(n119854), .B1(n99591), .B2(n119848), .ZN(
        n116756) );
  OAI22_X1 U85941 ( .A1(n98658), .A2(n119854), .B1(n99590), .B2(n119848), .ZN(
        n116733) );
  OAI22_X1 U85942 ( .A1(n98657), .A2(n119854), .B1(n99589), .B2(n119848), .ZN(
        n116710) );
  OAI22_X1 U85943 ( .A1(n98656), .A2(n119854), .B1(n99588), .B2(n119848), .ZN(
        n116687) );
  OAI22_X1 U85944 ( .A1(n98655), .A2(n119854), .B1(n99587), .B2(n119848), .ZN(
        n116664) );
  OAI22_X1 U85945 ( .A1(n98654), .A2(n119854), .B1(n99586), .B2(n119848), .ZN(
        n116641) );
  OAI22_X1 U85946 ( .A1(n98653), .A2(n119854), .B1(n99585), .B2(n119848), .ZN(
        n116618) );
  OAI22_X1 U85947 ( .A1(n98732), .A2(n120075), .B1(n99932), .B2(n120069), .ZN(
        n115171) );
  OAI22_X1 U85948 ( .A1(n98731), .A2(n120075), .B1(n99931), .B2(n120069), .ZN(
        n115143) );
  OAI22_X1 U85949 ( .A1(n98730), .A2(n120076), .B1(n99930), .B2(n120070), .ZN(
        n115115) );
  OAI22_X1 U85950 ( .A1(n98729), .A2(n120076), .B1(n99929), .B2(n120070), .ZN(
        n115087) );
  OAI22_X1 U85951 ( .A1(n98728), .A2(n120076), .B1(n99928), .B2(n120070), .ZN(
        n115059) );
  OAI22_X1 U85952 ( .A1(n98727), .A2(n120076), .B1(n99927), .B2(n120070), .ZN(
        n115031) );
  OAI22_X1 U85953 ( .A1(n98726), .A2(n120076), .B1(n99926), .B2(n120070), .ZN(
        n115003) );
  OAI22_X1 U85954 ( .A1(n98725), .A2(n120076), .B1(n99925), .B2(n120070), .ZN(
        n114975) );
  OAI22_X1 U85955 ( .A1(n98724), .A2(n120076), .B1(n99924), .B2(n120070), .ZN(
        n114947) );
  OAI22_X1 U85956 ( .A1(n98723), .A2(n120076), .B1(n99923), .B2(n120070), .ZN(
        n114919) );
  OAI22_X1 U85957 ( .A1(n98722), .A2(n120076), .B1(n99922), .B2(n120070), .ZN(
        n114891) );
  OAI22_X1 U85958 ( .A1(n98721), .A2(n120076), .B1(n99921), .B2(n120070), .ZN(
        n114863) );
  OAI22_X1 U85959 ( .A1(n98720), .A2(n120076), .B1(n99920), .B2(n120070), .ZN(
        n114835) );
  OAI22_X1 U85960 ( .A1(n98719), .A2(n120076), .B1(n99919), .B2(n120070), .ZN(
        n114807) );
  OAI22_X1 U85961 ( .A1(n98778), .A2(n120072), .B1(n99978), .B2(n120066), .ZN(
        n116474) );
  OAI22_X1 U85962 ( .A1(n98777), .A2(n120072), .B1(n99977), .B2(n120066), .ZN(
        n116431) );
  OAI22_X1 U85963 ( .A1(n98776), .A2(n120072), .B1(n99976), .B2(n120066), .ZN(
        n116403) );
  OAI22_X1 U85964 ( .A1(n98775), .A2(n120072), .B1(n99975), .B2(n120066), .ZN(
        n116375) );
  OAI22_X1 U85965 ( .A1(n98705), .A2(n119850), .B1(n99637), .B2(n119844), .ZN(
        n117802) );
  OAI22_X1 U85966 ( .A1(n98704), .A2(n119850), .B1(n99636), .B2(n119844), .ZN(
        n117780) );
  OAI22_X1 U85967 ( .A1(n98703), .A2(n119850), .B1(n99635), .B2(n119844), .ZN(
        n117758) );
  OAI22_X1 U85968 ( .A1(n98702), .A2(n119850), .B1(n99634), .B2(n119844), .ZN(
        n117736) );
  OAI22_X1 U85969 ( .A1(n98712), .A2(n119850), .B1(n99644), .B2(n119844), .ZN(
        n117972) );
  OAI22_X1 U85970 ( .A1(n98711), .A2(n119850), .B1(n99643), .B2(n119844), .ZN(
        n117934) );
  OAI22_X1 U85971 ( .A1(n98710), .A2(n119850), .B1(n99642), .B2(n119844), .ZN(
        n117912) );
  OAI22_X1 U85972 ( .A1(n98709), .A2(n119850), .B1(n99641), .B2(n119844), .ZN(
        n117890) );
  OAI22_X1 U85973 ( .A1(n98708), .A2(n119850), .B1(n99640), .B2(n119844), .ZN(
        n117868) );
  OAI22_X1 U85974 ( .A1(n98707), .A2(n119850), .B1(n99639), .B2(n119844), .ZN(
        n117846) );
  OAI22_X1 U85975 ( .A1(n98706), .A2(n119850), .B1(n99638), .B2(n119844), .ZN(
        n117824) );
  OAI22_X1 U85976 ( .A1(n98774), .A2(n120072), .B1(n99974), .B2(n120066), .ZN(
        n116347) );
  OAI22_X1 U85977 ( .A1(n98773), .A2(n120072), .B1(n99973), .B2(n120066), .ZN(
        n116319) );
  OAI22_X1 U85978 ( .A1(n98772), .A2(n120072), .B1(n99972), .B2(n120066), .ZN(
        n116291) );
  OAI22_X1 U85979 ( .A1(n98771), .A2(n120072), .B1(n99971), .B2(n120066), .ZN(
        n116263) );
  OAI22_X1 U85980 ( .A1(n98770), .A2(n120072), .B1(n99970), .B2(n120066), .ZN(
        n116235) );
  OAI22_X1 U85981 ( .A1(n98769), .A2(n120072), .B1(n99969), .B2(n120066), .ZN(
        n116207) );
  OAI22_X1 U85982 ( .A1(n98768), .A2(n120072), .B1(n99968), .B2(n120066), .ZN(
        n116179) );
  OAI22_X1 U85983 ( .A1(n98767), .A2(n120072), .B1(n99967), .B2(n120066), .ZN(
        n116151) );
  OAI22_X1 U85984 ( .A1(n98766), .A2(n120073), .B1(n99966), .B2(n120067), .ZN(
        n116123) );
  OAI22_X1 U85985 ( .A1(n98765), .A2(n120073), .B1(n99965), .B2(n120067), .ZN(
        n116095) );
  OAI22_X1 U85986 ( .A1(n98764), .A2(n120073), .B1(n99964), .B2(n120067), .ZN(
        n116067) );
  OAI22_X1 U85987 ( .A1(n98763), .A2(n120073), .B1(n99963), .B2(n120067), .ZN(
        n116039) );
  OAI22_X1 U85988 ( .A1(n98762), .A2(n120073), .B1(n99962), .B2(n120067), .ZN(
        n116011) );
  OAI22_X1 U85989 ( .A1(n98761), .A2(n120073), .B1(n99961), .B2(n120067), .ZN(
        n115983) );
  OAI22_X1 U85990 ( .A1(n98760), .A2(n120073), .B1(n99960), .B2(n120067), .ZN(
        n115955) );
  OAI22_X1 U85991 ( .A1(n98759), .A2(n120073), .B1(n99959), .B2(n120067), .ZN(
        n115927) );
  OAI22_X1 U85992 ( .A1(n98758), .A2(n120073), .B1(n99958), .B2(n120067), .ZN(
        n115899) );
  OAI22_X1 U85993 ( .A1(n98757), .A2(n120073), .B1(n99957), .B2(n120067), .ZN(
        n115871) );
  OAI22_X1 U85994 ( .A1(n98756), .A2(n120073), .B1(n99956), .B2(n120067), .ZN(
        n115843) );
  OAI22_X1 U85995 ( .A1(n98755), .A2(n120073), .B1(n99955), .B2(n120067), .ZN(
        n115815) );
  OAI22_X1 U85996 ( .A1(n98754), .A2(n120074), .B1(n99954), .B2(n120068), .ZN(
        n115787) );
  OAI22_X1 U85997 ( .A1(n98753), .A2(n120074), .B1(n99953), .B2(n120068), .ZN(
        n115759) );
  OAI22_X1 U85998 ( .A1(n98752), .A2(n120074), .B1(n99952), .B2(n120068), .ZN(
        n115731) );
  OAI22_X1 U85999 ( .A1(n98751), .A2(n120074), .B1(n99951), .B2(n120068), .ZN(
        n115703) );
  OAI22_X1 U86000 ( .A1(n98750), .A2(n120074), .B1(n99950), .B2(n120068), .ZN(
        n115675) );
  OAI22_X1 U86001 ( .A1(n98749), .A2(n120074), .B1(n99949), .B2(n120068), .ZN(
        n115647) );
  OAI22_X1 U86002 ( .A1(n98748), .A2(n120074), .B1(n99948), .B2(n120068), .ZN(
        n115619) );
  OAI22_X1 U86003 ( .A1(n98747), .A2(n120074), .B1(n99947), .B2(n120068), .ZN(
        n115591) );
  OAI22_X1 U86004 ( .A1(n98746), .A2(n120074), .B1(n99946), .B2(n120068), .ZN(
        n115563) );
  OAI22_X1 U86005 ( .A1(n98745), .A2(n120074), .B1(n99945), .B2(n120068), .ZN(
        n115535) );
  OAI22_X1 U86006 ( .A1(n98744), .A2(n120074), .B1(n99944), .B2(n120068), .ZN(
        n115507) );
  OAI22_X1 U86007 ( .A1(n98743), .A2(n120074), .B1(n99943), .B2(n120068), .ZN(
        n115479) );
  OAI22_X1 U86008 ( .A1(n98742), .A2(n120075), .B1(n99942), .B2(n120069), .ZN(
        n115451) );
  OAI22_X1 U86009 ( .A1(n98741), .A2(n120075), .B1(n99941), .B2(n120069), .ZN(
        n115423) );
  OAI22_X1 U86010 ( .A1(n98740), .A2(n120075), .B1(n99940), .B2(n120069), .ZN(
        n115395) );
  OAI22_X1 U86011 ( .A1(n98739), .A2(n120075), .B1(n99939), .B2(n120069), .ZN(
        n115367) );
  OAI22_X1 U86012 ( .A1(n98738), .A2(n120075), .B1(n99938), .B2(n120069), .ZN(
        n115339) );
  OAI22_X1 U86013 ( .A1(n98737), .A2(n120075), .B1(n99937), .B2(n120069), .ZN(
        n115311) );
  OAI22_X1 U86014 ( .A1(n98736), .A2(n120075), .B1(n99936), .B2(n120069), .ZN(
        n115283) );
  OAI22_X1 U86015 ( .A1(n98735), .A2(n120075), .B1(n99935), .B2(n120069), .ZN(
        n115255) );
  OAI22_X1 U86016 ( .A1(n98734), .A2(n120075), .B1(n99934), .B2(n120069), .ZN(
        n115227) );
  OAI22_X1 U86017 ( .A1(n98733), .A2(n120075), .B1(n99933), .B2(n120069), .ZN(
        n115199) );
  OAI22_X1 U86018 ( .A1(n114040), .A2(n119874), .B1(n99499), .B2(n119868), 
        .ZN(n117713) );
  OAI22_X1 U86019 ( .A1(n114039), .A2(n119875), .B1(n99498), .B2(n119869), 
        .ZN(n117691) );
  OAI22_X1 U86020 ( .A1(n114038), .A2(n119875), .B1(n99497), .B2(n119869), 
        .ZN(n117669) );
  OAI22_X1 U86021 ( .A1(n114037), .A2(n119875), .B1(n99496), .B2(n119869), 
        .ZN(n117647) );
  OAI22_X1 U86022 ( .A1(n114036), .A2(n119875), .B1(n99495), .B2(n119869), 
        .ZN(n117625) );
  OAI22_X1 U86023 ( .A1(n114035), .A2(n119875), .B1(n99494), .B2(n119869), 
        .ZN(n117603) );
  OAI22_X1 U86024 ( .A1(n114034), .A2(n119875), .B1(n99493), .B2(n119869), 
        .ZN(n117581) );
  OAI22_X1 U86025 ( .A1(n114033), .A2(n119875), .B1(n99492), .B2(n119869), 
        .ZN(n117559) );
  OAI22_X1 U86026 ( .A1(n114032), .A2(n119875), .B1(n99491), .B2(n119869), 
        .ZN(n117537) );
  OAI22_X1 U86027 ( .A1(n114031), .A2(n119875), .B1(n99490), .B2(n119869), 
        .ZN(n117514) );
  OAI22_X1 U86028 ( .A1(n114030), .A2(n119875), .B1(n99489), .B2(n119869), 
        .ZN(n117491) );
  OAI22_X1 U86029 ( .A1(n114029), .A2(n119875), .B1(n99488), .B2(n119869), 
        .ZN(n117468) );
  OAI22_X1 U86030 ( .A1(n114028), .A2(n119875), .B1(n99487), .B2(n119869), 
        .ZN(n117445) );
  OAI22_X1 U86031 ( .A1(n114027), .A2(n119876), .B1(n99486), .B2(n119870), 
        .ZN(n117422) );
  OAI22_X1 U86032 ( .A1(n114026), .A2(n119876), .B1(n99485), .B2(n119870), 
        .ZN(n117399) );
  OAI22_X1 U86033 ( .A1(n114025), .A2(n119876), .B1(n99484), .B2(n119870), 
        .ZN(n117376) );
  OAI22_X1 U86034 ( .A1(n114024), .A2(n119876), .B1(n99483), .B2(n119870), 
        .ZN(n117353) );
  OAI22_X1 U86035 ( .A1(n114023), .A2(n119876), .B1(n99482), .B2(n119870), 
        .ZN(n117330) );
  OAI22_X1 U86036 ( .A1(n114022), .A2(n119876), .B1(n99481), .B2(n119870), 
        .ZN(n117307) );
  OAI22_X1 U86037 ( .A1(n114021), .A2(n119876), .B1(n99480), .B2(n119870), 
        .ZN(n117284) );
  OAI22_X1 U86038 ( .A1(n114020), .A2(n119876), .B1(n99479), .B2(n119870), 
        .ZN(n117261) );
  OAI22_X1 U86039 ( .A1(n114019), .A2(n119876), .B1(n99478), .B2(n119870), 
        .ZN(n117238) );
  OAI22_X1 U86040 ( .A1(n114018), .A2(n119876), .B1(n99477), .B2(n119870), 
        .ZN(n117215) );
  OAI22_X1 U86041 ( .A1(n114017), .A2(n119876), .B1(n99476), .B2(n119870), 
        .ZN(n117192) );
  OAI22_X1 U86042 ( .A1(n114016), .A2(n119876), .B1(n99475), .B2(n119870), 
        .ZN(n117169) );
  OAI22_X1 U86043 ( .A1(n114015), .A2(n119877), .B1(n99474), .B2(n119871), 
        .ZN(n117146) );
  OAI22_X1 U86044 ( .A1(n114014), .A2(n119877), .B1(n99473), .B2(n119871), 
        .ZN(n117123) );
  OAI22_X1 U86045 ( .A1(n114013), .A2(n119877), .B1(n99472), .B2(n119871), 
        .ZN(n117100) );
  OAI22_X1 U86046 ( .A1(n114012), .A2(n119877), .B1(n99471), .B2(n119871), 
        .ZN(n117077) );
  OAI22_X1 U86047 ( .A1(n114011), .A2(n119877), .B1(n99470), .B2(n119871), 
        .ZN(n117054) );
  OAI22_X1 U86048 ( .A1(n114010), .A2(n119877), .B1(n99469), .B2(n119871), 
        .ZN(n117031) );
  OAI22_X1 U86049 ( .A1(n114009), .A2(n119877), .B1(n99468), .B2(n119871), 
        .ZN(n117008) );
  OAI22_X1 U86050 ( .A1(n114008), .A2(n119877), .B1(n99467), .B2(n119871), 
        .ZN(n116985) );
  OAI22_X1 U86051 ( .A1(n114007), .A2(n119877), .B1(n99466), .B2(n119871), 
        .ZN(n116962) );
  OAI22_X1 U86052 ( .A1(n114006), .A2(n119877), .B1(n99465), .B2(n119871), 
        .ZN(n116939) );
  OAI22_X1 U86053 ( .A1(n114005), .A2(n119877), .B1(n99464), .B2(n119871), 
        .ZN(n116916) );
  OAI22_X1 U86054 ( .A1(n114004), .A2(n119877), .B1(n99463), .B2(n119871), 
        .ZN(n116893) );
  OAI22_X1 U86055 ( .A1(n114003), .A2(n119878), .B1(n99462), .B2(n119872), 
        .ZN(n116870) );
  OAI22_X1 U86056 ( .A1(n114002), .A2(n119878), .B1(n99461), .B2(n119872), 
        .ZN(n116847) );
  OAI22_X1 U86057 ( .A1(n114001), .A2(n119878), .B1(n99460), .B2(n119872), 
        .ZN(n116824) );
  OAI22_X1 U86058 ( .A1(n114000), .A2(n119878), .B1(n99459), .B2(n119872), 
        .ZN(n116801) );
  OAI22_X1 U86059 ( .A1(n113999), .A2(n119878), .B1(n99458), .B2(n119872), 
        .ZN(n116778) );
  OAI22_X1 U86060 ( .A1(n113998), .A2(n119878), .B1(n99457), .B2(n119872), 
        .ZN(n116755) );
  OAI22_X1 U86061 ( .A1(n113997), .A2(n119878), .B1(n99456), .B2(n119872), 
        .ZN(n116732) );
  OAI22_X1 U86062 ( .A1(n113996), .A2(n119878), .B1(n99455), .B2(n119872), 
        .ZN(n116709) );
  OAI22_X1 U86063 ( .A1(n113995), .A2(n119878), .B1(n99454), .B2(n119872), 
        .ZN(n116686) );
  OAI22_X1 U86064 ( .A1(n113994), .A2(n119878), .B1(n99453), .B2(n119872), 
        .ZN(n116663) );
  OAI22_X1 U86065 ( .A1(n113993), .A2(n119878), .B1(n99452), .B2(n119872), 
        .ZN(n116640) );
  OAI22_X1 U86066 ( .A1(n113992), .A2(n119878), .B1(n99451), .B2(n119872), 
        .ZN(n116617) );
  OAI22_X1 U86067 ( .A1(n114044), .A2(n119874), .B1(n99503), .B2(n119868), 
        .ZN(n117801) );
  OAI22_X1 U86068 ( .A1(n114043), .A2(n119874), .B1(n99502), .B2(n119868), 
        .ZN(n117779) );
  OAI22_X1 U86069 ( .A1(n114042), .A2(n119874), .B1(n99501), .B2(n119868), 
        .ZN(n117757) );
  OAI22_X1 U86070 ( .A1(n114041), .A2(n119874), .B1(n99500), .B2(n119868), 
        .ZN(n117735) );
  OAI22_X1 U86071 ( .A1(n114051), .A2(n119874), .B1(n99510), .B2(n119868), 
        .ZN(n117969) );
  OAI22_X1 U86072 ( .A1(n114050), .A2(n119874), .B1(n99509), .B2(n119868), 
        .ZN(n117933) );
  OAI22_X1 U86073 ( .A1(n114049), .A2(n119874), .B1(n99508), .B2(n119868), 
        .ZN(n117911) );
  OAI22_X1 U86074 ( .A1(n114048), .A2(n119874), .B1(n99507), .B2(n119868), 
        .ZN(n117889) );
  OAI22_X1 U86075 ( .A1(n114047), .A2(n119874), .B1(n99506), .B2(n119868), 
        .ZN(n117867) );
  OAI22_X1 U86076 ( .A1(n114046), .A2(n119874), .B1(n99505), .B2(n119868), 
        .ZN(n117845) );
  OAI22_X1 U86077 ( .A1(n114045), .A2(n119874), .B1(n99504), .B2(n119868), 
        .ZN(n117823) );
  OAI22_X1 U86078 ( .A1(n99769), .A2(n119940), .B1(n113868), .B2(n119934), 
        .ZN(n117712) );
  OAI22_X1 U86079 ( .A1(n99768), .A2(n119941), .B1(n113866), .B2(n119935), 
        .ZN(n117690) );
  OAI22_X1 U86080 ( .A1(n99767), .A2(n119941), .B1(n113864), .B2(n119935), 
        .ZN(n117668) );
  OAI22_X1 U86081 ( .A1(n99766), .A2(n119941), .B1(n113862), .B2(n119935), 
        .ZN(n117646) );
  OAI22_X1 U86082 ( .A1(n99765), .A2(n119941), .B1(n113860), .B2(n119935), 
        .ZN(n117624) );
  OAI22_X1 U86083 ( .A1(n99764), .A2(n119941), .B1(n113858), .B2(n119935), 
        .ZN(n117602) );
  OAI22_X1 U86084 ( .A1(n99763), .A2(n119941), .B1(n113856), .B2(n119935), 
        .ZN(n117580) );
  OAI22_X1 U86085 ( .A1(n99762), .A2(n119941), .B1(n113854), .B2(n119935), 
        .ZN(n117558) );
  OAI22_X1 U86086 ( .A1(n99761), .A2(n119941), .B1(n113852), .B2(n119935), 
        .ZN(n117535) );
  OAI22_X1 U86087 ( .A1(n99760), .A2(n119941), .B1(n113850), .B2(n119935), 
        .ZN(n117512) );
  OAI22_X1 U86088 ( .A1(n99759), .A2(n119941), .B1(n113848), .B2(n119935), 
        .ZN(n117489) );
  OAI22_X1 U86089 ( .A1(n99758), .A2(n119941), .B1(n113846), .B2(n119935), 
        .ZN(n117466) );
  OAI22_X1 U86090 ( .A1(n99757), .A2(n119941), .B1(n113844), .B2(n119935), 
        .ZN(n117443) );
  OAI22_X1 U86091 ( .A1(n99756), .A2(n119942), .B1(n113842), .B2(n119936), 
        .ZN(n117420) );
  OAI22_X1 U86092 ( .A1(n99755), .A2(n119942), .B1(n113840), .B2(n119936), 
        .ZN(n117397) );
  OAI22_X1 U86093 ( .A1(n99754), .A2(n119942), .B1(n113838), .B2(n119936), 
        .ZN(n117374) );
  OAI22_X1 U86094 ( .A1(n99753), .A2(n119942), .B1(n113836), .B2(n119936), 
        .ZN(n117351) );
  OAI22_X1 U86095 ( .A1(n99752), .A2(n119942), .B1(n113834), .B2(n119936), 
        .ZN(n117328) );
  OAI22_X1 U86096 ( .A1(n99751), .A2(n119942), .B1(n113832), .B2(n119936), 
        .ZN(n117305) );
  OAI22_X1 U86097 ( .A1(n99750), .A2(n119942), .B1(n113830), .B2(n119936), 
        .ZN(n117282) );
  OAI22_X1 U86098 ( .A1(n99749), .A2(n119942), .B1(n113828), .B2(n119936), 
        .ZN(n117259) );
  OAI22_X1 U86099 ( .A1(n99748), .A2(n119942), .B1(n113826), .B2(n119936), 
        .ZN(n117236) );
  OAI22_X1 U86100 ( .A1(n99747), .A2(n119942), .B1(n113824), .B2(n119936), 
        .ZN(n117213) );
  OAI22_X1 U86101 ( .A1(n99746), .A2(n119942), .B1(n113822), .B2(n119936), 
        .ZN(n117190) );
  OAI22_X1 U86102 ( .A1(n99745), .A2(n119942), .B1(n113820), .B2(n119936), 
        .ZN(n117167) );
  OAI22_X1 U86103 ( .A1(n99744), .A2(n119943), .B1(n113818), .B2(n119937), 
        .ZN(n117144) );
  OAI22_X1 U86104 ( .A1(n99743), .A2(n119943), .B1(n113816), .B2(n119937), 
        .ZN(n117121) );
  OAI22_X1 U86105 ( .A1(n99742), .A2(n119943), .B1(n113814), .B2(n119937), 
        .ZN(n117098) );
  OAI22_X1 U86106 ( .A1(n99741), .A2(n119943), .B1(n113812), .B2(n119937), 
        .ZN(n117075) );
  OAI22_X1 U86107 ( .A1(n99740), .A2(n119943), .B1(n113810), .B2(n119937), 
        .ZN(n117052) );
  OAI22_X1 U86108 ( .A1(n99739), .A2(n119943), .B1(n113808), .B2(n119937), 
        .ZN(n117029) );
  OAI22_X1 U86109 ( .A1(n99738), .A2(n119943), .B1(n113806), .B2(n119937), 
        .ZN(n117006) );
  OAI22_X1 U86110 ( .A1(n99737), .A2(n119943), .B1(n113804), .B2(n119937), 
        .ZN(n116983) );
  OAI22_X1 U86111 ( .A1(n99736), .A2(n119943), .B1(n113802), .B2(n119937), 
        .ZN(n116960) );
  OAI22_X1 U86112 ( .A1(n99735), .A2(n119943), .B1(n113800), .B2(n119937), 
        .ZN(n116937) );
  OAI22_X1 U86113 ( .A1(n99734), .A2(n119943), .B1(n113798), .B2(n119937), 
        .ZN(n116914) );
  OAI22_X1 U86114 ( .A1(n99733), .A2(n119943), .B1(n113796), .B2(n119937), 
        .ZN(n116891) );
  OAI22_X1 U86115 ( .A1(n99732), .A2(n119944), .B1(n113794), .B2(n119938), 
        .ZN(n116868) );
  OAI22_X1 U86116 ( .A1(n99731), .A2(n119944), .B1(n113792), .B2(n119938), 
        .ZN(n116845) );
  OAI22_X1 U86117 ( .A1(n99730), .A2(n119944), .B1(n113790), .B2(n119938), 
        .ZN(n116822) );
  OAI22_X1 U86118 ( .A1(n99729), .A2(n119944), .B1(n113788), .B2(n119938), 
        .ZN(n116799) );
  OAI22_X1 U86119 ( .A1(n99728), .A2(n119944), .B1(n113786), .B2(n119938), 
        .ZN(n116776) );
  OAI22_X1 U86120 ( .A1(n99727), .A2(n119944), .B1(n113784), .B2(n119938), 
        .ZN(n116753) );
  OAI22_X1 U86121 ( .A1(n99726), .A2(n119944), .B1(n113782), .B2(n119938), 
        .ZN(n116730) );
  OAI22_X1 U86122 ( .A1(n99725), .A2(n119944), .B1(n113780), .B2(n119938), 
        .ZN(n116707) );
  OAI22_X1 U86123 ( .A1(n99724), .A2(n119944), .B1(n113778), .B2(n119938), 
        .ZN(n116684) );
  OAI22_X1 U86124 ( .A1(n99723), .A2(n119944), .B1(n113776), .B2(n119938), 
        .ZN(n116661) );
  OAI22_X1 U86125 ( .A1(n99722), .A2(n119944), .B1(n113774), .B2(n119938), 
        .ZN(n116638) );
  OAI22_X1 U86126 ( .A1(n99721), .A2(n119944), .B1(n113772), .B2(n119938), 
        .ZN(n116615) );
  OAI22_X1 U86127 ( .A1(n99065), .A2(n120141), .B1(n113798), .B2(n120135), 
        .ZN(n115168) );
  OAI22_X1 U86128 ( .A1(n99064), .A2(n120141), .B1(n113796), .B2(n120135), 
        .ZN(n115140) );
  OAI22_X1 U86129 ( .A1(n99063), .A2(n120142), .B1(n113794), .B2(n120136), 
        .ZN(n115112) );
  OAI22_X1 U86130 ( .A1(n99062), .A2(n120142), .B1(n113792), .B2(n120136), 
        .ZN(n115084) );
  OAI22_X1 U86131 ( .A1(n99061), .A2(n120142), .B1(n113790), .B2(n120136), 
        .ZN(n115056) );
  OAI22_X1 U86132 ( .A1(n99060), .A2(n120142), .B1(n113788), .B2(n120136), 
        .ZN(n115028) );
  OAI22_X1 U86133 ( .A1(n99059), .A2(n120142), .B1(n113786), .B2(n120136), 
        .ZN(n115000) );
  OAI22_X1 U86134 ( .A1(n99058), .A2(n120142), .B1(n113784), .B2(n120136), 
        .ZN(n114972) );
  OAI22_X1 U86135 ( .A1(n99057), .A2(n120142), .B1(n113782), .B2(n120136), 
        .ZN(n114944) );
  OAI22_X1 U86136 ( .A1(n99056), .A2(n120142), .B1(n113780), .B2(n120136), 
        .ZN(n114916) );
  OAI22_X1 U86137 ( .A1(n99055), .A2(n120142), .B1(n113778), .B2(n120136), 
        .ZN(n114888) );
  OAI22_X1 U86138 ( .A1(n99054), .A2(n120142), .B1(n113776), .B2(n120136), 
        .ZN(n114860) );
  OAI22_X1 U86139 ( .A1(n99053), .A2(n120142), .B1(n113774), .B2(n120136), 
        .ZN(n114832) );
  OAI22_X1 U86140 ( .A1(n99052), .A2(n120142), .B1(n113772), .B2(n120136), 
        .ZN(n114804) );
  OAI22_X1 U86141 ( .A1(n99111), .A2(n120138), .B1(n113890), .B2(n120132), 
        .ZN(n116468) );
  OAI22_X1 U86142 ( .A1(n99110), .A2(n120138), .B1(n113888), .B2(n120132), 
        .ZN(n116428) );
  OAI22_X1 U86143 ( .A1(n99109), .A2(n120138), .B1(n113886), .B2(n120132), 
        .ZN(n116400) );
  OAI22_X1 U86144 ( .A1(n99108), .A2(n120138), .B1(n113884), .B2(n120132), 
        .ZN(n116372) );
  OAI22_X1 U86145 ( .A1(n99773), .A2(n119940), .B1(n113876), .B2(n119934), 
        .ZN(n117800) );
  OAI22_X1 U86146 ( .A1(n99772), .A2(n119940), .B1(n113874), .B2(n119934), 
        .ZN(n117778) );
  OAI22_X1 U86147 ( .A1(n99771), .A2(n119940), .B1(n113872), .B2(n119934), 
        .ZN(n117756) );
  OAI22_X1 U86148 ( .A1(n99770), .A2(n119940), .B1(n113870), .B2(n119934), 
        .ZN(n117734) );
  OAI22_X1 U86149 ( .A1(n99780), .A2(n119940), .B1(n113890), .B2(n119934), 
        .ZN(n117966) );
  OAI22_X1 U86150 ( .A1(n99779), .A2(n119940), .B1(n113888), .B2(n119934), 
        .ZN(n117932) );
  OAI22_X1 U86151 ( .A1(n99778), .A2(n119940), .B1(n113886), .B2(n119934), 
        .ZN(n117910) );
  OAI22_X1 U86152 ( .A1(n99777), .A2(n119940), .B1(n113884), .B2(n119934), 
        .ZN(n117888) );
  OAI22_X1 U86153 ( .A1(n99776), .A2(n119940), .B1(n113882), .B2(n119934), 
        .ZN(n117866) );
  OAI22_X1 U86154 ( .A1(n99775), .A2(n119940), .B1(n113880), .B2(n119934), 
        .ZN(n117844) );
  OAI22_X1 U86155 ( .A1(n99774), .A2(n119940), .B1(n113878), .B2(n119934), 
        .ZN(n117822) );
  OAI22_X1 U86156 ( .A1(n99107), .A2(n120138), .B1(n113882), .B2(n120132), 
        .ZN(n116344) );
  OAI22_X1 U86157 ( .A1(n99106), .A2(n120138), .B1(n113880), .B2(n120132), 
        .ZN(n116316) );
  OAI22_X1 U86158 ( .A1(n99105), .A2(n120138), .B1(n113878), .B2(n120132), 
        .ZN(n116288) );
  OAI22_X1 U86159 ( .A1(n99104), .A2(n120138), .B1(n113876), .B2(n120132), 
        .ZN(n116260) );
  OAI22_X1 U86160 ( .A1(n99103), .A2(n120138), .B1(n113874), .B2(n120132), 
        .ZN(n116232) );
  OAI22_X1 U86161 ( .A1(n99102), .A2(n120138), .B1(n113872), .B2(n120132), 
        .ZN(n116204) );
  OAI22_X1 U86162 ( .A1(n99101), .A2(n120138), .B1(n113870), .B2(n120132), 
        .ZN(n116176) );
  OAI22_X1 U86163 ( .A1(n99100), .A2(n120138), .B1(n113868), .B2(n120132), 
        .ZN(n116148) );
  OAI22_X1 U86164 ( .A1(n99099), .A2(n120139), .B1(n113866), .B2(n120133), 
        .ZN(n116120) );
  OAI22_X1 U86165 ( .A1(n99098), .A2(n120139), .B1(n113864), .B2(n120133), 
        .ZN(n116092) );
  OAI22_X1 U86166 ( .A1(n99097), .A2(n120139), .B1(n113862), .B2(n120133), 
        .ZN(n116064) );
  OAI22_X1 U86167 ( .A1(n99096), .A2(n120139), .B1(n113860), .B2(n120133), 
        .ZN(n116036) );
  OAI22_X1 U86168 ( .A1(n99095), .A2(n120139), .B1(n113858), .B2(n120133), 
        .ZN(n116008) );
  OAI22_X1 U86169 ( .A1(n99094), .A2(n120139), .B1(n113856), .B2(n120133), 
        .ZN(n115980) );
  OAI22_X1 U86170 ( .A1(n99093), .A2(n120139), .B1(n113854), .B2(n120133), 
        .ZN(n115952) );
  OAI22_X1 U86171 ( .A1(n99092), .A2(n120139), .B1(n113852), .B2(n120133), 
        .ZN(n115924) );
  OAI22_X1 U86172 ( .A1(n99091), .A2(n120139), .B1(n113850), .B2(n120133), 
        .ZN(n115896) );
  OAI22_X1 U86173 ( .A1(n99090), .A2(n120139), .B1(n113848), .B2(n120133), 
        .ZN(n115868) );
  OAI22_X1 U86174 ( .A1(n99089), .A2(n120139), .B1(n113846), .B2(n120133), 
        .ZN(n115840) );
  OAI22_X1 U86175 ( .A1(n99088), .A2(n120139), .B1(n113844), .B2(n120133), 
        .ZN(n115812) );
  OAI22_X1 U86176 ( .A1(n99087), .A2(n120140), .B1(n113842), .B2(n120134), 
        .ZN(n115784) );
  OAI22_X1 U86177 ( .A1(n99086), .A2(n120140), .B1(n113840), .B2(n120134), 
        .ZN(n115756) );
  OAI22_X1 U86178 ( .A1(n99085), .A2(n120140), .B1(n113838), .B2(n120134), 
        .ZN(n115728) );
  OAI22_X1 U86179 ( .A1(n99084), .A2(n120140), .B1(n113836), .B2(n120134), 
        .ZN(n115700) );
  OAI22_X1 U86180 ( .A1(n99083), .A2(n120140), .B1(n113834), .B2(n120134), 
        .ZN(n115672) );
  OAI22_X1 U86181 ( .A1(n99082), .A2(n120140), .B1(n113832), .B2(n120134), 
        .ZN(n115644) );
  OAI22_X1 U86182 ( .A1(n99081), .A2(n120140), .B1(n113830), .B2(n120134), 
        .ZN(n115616) );
  OAI22_X1 U86183 ( .A1(n99080), .A2(n120140), .B1(n113828), .B2(n120134), 
        .ZN(n115588) );
  OAI22_X1 U86184 ( .A1(n99079), .A2(n120140), .B1(n113826), .B2(n120134), 
        .ZN(n115560) );
  OAI22_X1 U86185 ( .A1(n99078), .A2(n120140), .B1(n113824), .B2(n120134), 
        .ZN(n115532) );
  OAI22_X1 U86186 ( .A1(n99077), .A2(n120140), .B1(n113822), .B2(n120134), 
        .ZN(n115504) );
  OAI22_X1 U86187 ( .A1(n99076), .A2(n120140), .B1(n113820), .B2(n120134), 
        .ZN(n115476) );
  OAI22_X1 U86188 ( .A1(n99075), .A2(n120141), .B1(n113818), .B2(n120135), 
        .ZN(n115448) );
  OAI22_X1 U86189 ( .A1(n99074), .A2(n120141), .B1(n113816), .B2(n120135), 
        .ZN(n115420) );
  OAI22_X1 U86190 ( .A1(n99073), .A2(n120141), .B1(n113814), .B2(n120135), 
        .ZN(n115392) );
  OAI22_X1 U86191 ( .A1(n99072), .A2(n120141), .B1(n113812), .B2(n120135), 
        .ZN(n115364) );
  OAI22_X1 U86192 ( .A1(n99071), .A2(n120141), .B1(n113810), .B2(n120135), 
        .ZN(n115336) );
  OAI22_X1 U86193 ( .A1(n99070), .A2(n120141), .B1(n113808), .B2(n120135), 
        .ZN(n115308) );
  OAI22_X1 U86194 ( .A1(n99069), .A2(n120141), .B1(n113806), .B2(n120135), 
        .ZN(n115280) );
  OAI22_X1 U86195 ( .A1(n99068), .A2(n120141), .B1(n113804), .B2(n120135), 
        .ZN(n115252) );
  OAI22_X1 U86196 ( .A1(n99067), .A2(n120141), .B1(n113802), .B2(n120135), 
        .ZN(n115224) );
  OAI22_X1 U86197 ( .A1(n99066), .A2(n120141), .B1(n113800), .B2(n120135), 
        .ZN(n115196) );
  OAI22_X1 U86198 ( .A1(n98767), .A2(n119916), .B1(n90426), .B2(n119910), .ZN(
        n117710) );
  OAI22_X1 U86199 ( .A1(n98766), .A2(n119917), .B1(n90425), .B2(n119911), .ZN(
        n117688) );
  OAI22_X1 U86200 ( .A1(n98765), .A2(n119917), .B1(n90424), .B2(n119911), .ZN(
        n117666) );
  OAI22_X1 U86201 ( .A1(n98764), .A2(n119917), .B1(n90423), .B2(n119911), .ZN(
        n117644) );
  OAI22_X1 U86202 ( .A1(n98763), .A2(n119917), .B1(n90422), .B2(n119911), .ZN(
        n117622) );
  OAI22_X1 U86203 ( .A1(n98762), .A2(n119917), .B1(n90421), .B2(n119911), .ZN(
        n117600) );
  OAI22_X1 U86204 ( .A1(n98761), .A2(n119917), .B1(n90420), .B2(n119911), .ZN(
        n117578) );
  OAI22_X1 U86205 ( .A1(n98760), .A2(n119917), .B1(n90419), .B2(n119911), .ZN(
        n117556) );
  OAI22_X1 U86206 ( .A1(n98759), .A2(n119917), .B1(n90418), .B2(n119911), .ZN(
        n117533) );
  OAI22_X1 U86207 ( .A1(n98758), .A2(n119917), .B1(n90417), .B2(n119911), .ZN(
        n117510) );
  OAI22_X1 U86208 ( .A1(n98757), .A2(n119917), .B1(n90416), .B2(n119911), .ZN(
        n117487) );
  OAI22_X1 U86209 ( .A1(n98756), .A2(n119917), .B1(n90415), .B2(n119911), .ZN(
        n117464) );
  OAI22_X1 U86210 ( .A1(n98755), .A2(n119917), .B1(n90414), .B2(n119911), .ZN(
        n117441) );
  OAI22_X1 U86211 ( .A1(n98754), .A2(n119918), .B1(n90413), .B2(n119912), .ZN(
        n117418) );
  OAI22_X1 U86212 ( .A1(n98753), .A2(n119918), .B1(n90412), .B2(n119912), .ZN(
        n117395) );
  OAI22_X1 U86213 ( .A1(n98752), .A2(n119918), .B1(n90411), .B2(n119912), .ZN(
        n117372) );
  OAI22_X1 U86214 ( .A1(n98751), .A2(n119918), .B1(n90410), .B2(n119912), .ZN(
        n117349) );
  OAI22_X1 U86215 ( .A1(n98750), .A2(n119918), .B1(n90409), .B2(n119912), .ZN(
        n117326) );
  OAI22_X1 U86216 ( .A1(n98749), .A2(n119918), .B1(n90408), .B2(n119912), .ZN(
        n117303) );
  OAI22_X1 U86217 ( .A1(n98748), .A2(n119918), .B1(n90407), .B2(n119912), .ZN(
        n117280) );
  OAI22_X1 U86218 ( .A1(n98747), .A2(n119918), .B1(n90406), .B2(n119912), .ZN(
        n117257) );
  OAI22_X1 U86219 ( .A1(n98746), .A2(n119918), .B1(n90405), .B2(n119912), .ZN(
        n117234) );
  OAI22_X1 U86220 ( .A1(n98745), .A2(n119918), .B1(n90404), .B2(n119912), .ZN(
        n117211) );
  OAI22_X1 U86221 ( .A1(n98744), .A2(n119918), .B1(n90403), .B2(n119912), .ZN(
        n117188) );
  OAI22_X1 U86222 ( .A1(n98743), .A2(n119918), .B1(n90402), .B2(n119912), .ZN(
        n117165) );
  OAI22_X1 U86223 ( .A1(n98742), .A2(n119919), .B1(n90401), .B2(n119913), .ZN(
        n117142) );
  OAI22_X1 U86224 ( .A1(n98741), .A2(n119919), .B1(n90400), .B2(n119913), .ZN(
        n117119) );
  OAI22_X1 U86225 ( .A1(n98740), .A2(n119919), .B1(n90399), .B2(n119913), .ZN(
        n117096) );
  OAI22_X1 U86226 ( .A1(n98739), .A2(n119919), .B1(n90398), .B2(n119913), .ZN(
        n117073) );
  OAI22_X1 U86227 ( .A1(n98738), .A2(n119919), .B1(n90397), .B2(n119913), .ZN(
        n117050) );
  OAI22_X1 U86228 ( .A1(n98737), .A2(n119919), .B1(n90396), .B2(n119913), .ZN(
        n117027) );
  OAI22_X1 U86229 ( .A1(n98736), .A2(n119919), .B1(n90395), .B2(n119913), .ZN(
        n117004) );
  OAI22_X1 U86230 ( .A1(n98735), .A2(n119919), .B1(n90394), .B2(n119913), .ZN(
        n116981) );
  OAI22_X1 U86231 ( .A1(n98734), .A2(n119919), .B1(n90393), .B2(n119913), .ZN(
        n116958) );
  OAI22_X1 U86232 ( .A1(n98733), .A2(n119919), .B1(n90392), .B2(n119913), .ZN(
        n116935) );
  OAI22_X1 U86233 ( .A1(n98732), .A2(n119919), .B1(n90391), .B2(n119913), .ZN(
        n116912) );
  OAI22_X1 U86234 ( .A1(n98731), .A2(n119919), .B1(n90390), .B2(n119913), .ZN(
        n116889) );
  OAI22_X1 U86235 ( .A1(n98730), .A2(n119920), .B1(n90389), .B2(n119914), .ZN(
        n116866) );
  OAI22_X1 U86236 ( .A1(n98729), .A2(n119920), .B1(n90388), .B2(n119914), .ZN(
        n116843) );
  OAI22_X1 U86237 ( .A1(n98728), .A2(n119920), .B1(n90387), .B2(n119914), .ZN(
        n116820) );
  OAI22_X1 U86238 ( .A1(n98727), .A2(n119920), .B1(n90386), .B2(n119914), .ZN(
        n116797) );
  OAI22_X1 U86239 ( .A1(n98726), .A2(n119920), .B1(n90385), .B2(n119914), .ZN(
        n116774) );
  OAI22_X1 U86240 ( .A1(n98725), .A2(n119920), .B1(n90384), .B2(n119914), .ZN(
        n116751) );
  OAI22_X1 U86241 ( .A1(n98724), .A2(n119920), .B1(n90383), .B2(n119914), .ZN(
        n116728) );
  OAI22_X1 U86242 ( .A1(n98723), .A2(n119920), .B1(n90382), .B2(n119914), .ZN(
        n116705) );
  OAI22_X1 U86243 ( .A1(n98722), .A2(n119920), .B1(n90381), .B2(n119914), .ZN(
        n116682) );
  OAI22_X1 U86244 ( .A1(n98721), .A2(n119920), .B1(n90380), .B2(n119914), .ZN(
        n116659) );
  OAI22_X1 U86245 ( .A1(n98720), .A2(n119920), .B1(n90379), .B2(n119914), .ZN(
        n116636) );
  OAI22_X1 U86246 ( .A1(n98719), .A2(n119920), .B1(n90378), .B2(n119914), .ZN(
        n116613) );
  OAI22_X1 U86247 ( .A1(n90530), .A2(n120117), .B1(n90049), .B2(n120111), .ZN(
        n115166) );
  OAI22_X1 U86248 ( .A1(n90529), .A2(n120117), .B1(n90048), .B2(n120111), .ZN(
        n115138) );
  OAI22_X1 U86249 ( .A1(n90528), .A2(n120118), .B1(n90047), .B2(n120112), .ZN(
        n115110) );
  OAI22_X1 U86250 ( .A1(n90527), .A2(n120118), .B1(n90046), .B2(n120112), .ZN(
        n115082) );
  OAI22_X1 U86251 ( .A1(n90526), .A2(n120118), .B1(n90045), .B2(n120112), .ZN(
        n115054) );
  OAI22_X1 U86252 ( .A1(n90525), .A2(n120118), .B1(n90044), .B2(n120112), .ZN(
        n115026) );
  OAI22_X1 U86253 ( .A1(n90524), .A2(n120118), .B1(n90043), .B2(n120112), .ZN(
        n114998) );
  OAI22_X1 U86254 ( .A1(n90523), .A2(n120118), .B1(n90042), .B2(n120112), .ZN(
        n114970) );
  OAI22_X1 U86255 ( .A1(n90522), .A2(n120118), .B1(n90041), .B2(n120112), .ZN(
        n114942) );
  OAI22_X1 U86256 ( .A1(n90521), .A2(n120118), .B1(n90040), .B2(n120112), .ZN(
        n114914) );
  OAI22_X1 U86257 ( .A1(n90520), .A2(n120118), .B1(n90039), .B2(n120112), .ZN(
        n114886) );
  OAI22_X1 U86258 ( .A1(n90519), .A2(n120118), .B1(n90038), .B2(n120112), .ZN(
        n114858) );
  OAI22_X1 U86259 ( .A1(n90518), .A2(n120118), .B1(n90037), .B2(n120112), .ZN(
        n114830) );
  OAI22_X1 U86260 ( .A1(n90517), .A2(n120118), .B1(n90036), .B2(n120112), .ZN(
        n114802) );
  OAI22_X1 U86261 ( .A1(n114233), .A2(n120114), .B1(n90095), .B2(n120108), 
        .ZN(n116466) );
  OAI22_X1 U86262 ( .A1(n114232), .A2(n120114), .B1(n90094), .B2(n120108), 
        .ZN(n116426) );
  OAI22_X1 U86263 ( .A1(n114231), .A2(n120114), .B1(n90093), .B2(n120108), 
        .ZN(n116398) );
  OAI22_X1 U86264 ( .A1(n114230), .A2(n120114), .B1(n90092), .B2(n120108), 
        .ZN(n116370) );
  OAI22_X1 U86265 ( .A1(n98771), .A2(n119916), .B1(n90430), .B2(n119910), .ZN(
        n117798) );
  OAI22_X1 U86266 ( .A1(n98770), .A2(n119916), .B1(n90429), .B2(n119910), .ZN(
        n117776) );
  OAI22_X1 U86267 ( .A1(n98769), .A2(n119916), .B1(n90428), .B2(n119910), .ZN(
        n117754) );
  OAI22_X1 U86268 ( .A1(n98768), .A2(n119916), .B1(n90427), .B2(n119910), .ZN(
        n117732) );
  OAI22_X1 U86269 ( .A1(n98778), .A2(n119916), .B1(n90437), .B2(n119910), .ZN(
        n117964) );
  OAI22_X1 U86270 ( .A1(n98777), .A2(n119916), .B1(n90436), .B2(n119910), .ZN(
        n117930) );
  OAI22_X1 U86271 ( .A1(n98776), .A2(n119916), .B1(n90435), .B2(n119910), .ZN(
        n117908) );
  OAI22_X1 U86272 ( .A1(n98775), .A2(n119916), .B1(n90434), .B2(n119910), .ZN(
        n117886) );
  OAI22_X1 U86273 ( .A1(n98774), .A2(n119916), .B1(n90433), .B2(n119910), .ZN(
        n117864) );
  OAI22_X1 U86274 ( .A1(n98773), .A2(n119916), .B1(n90432), .B2(n119910), .ZN(
        n117842) );
  OAI22_X1 U86275 ( .A1(n98772), .A2(n119916), .B1(n90431), .B2(n119910), .ZN(
        n117820) );
  OAI22_X1 U86276 ( .A1(n114229), .A2(n120114), .B1(n90091), .B2(n120108), 
        .ZN(n116342) );
  OAI22_X1 U86277 ( .A1(n114228), .A2(n120114), .B1(n90090), .B2(n120108), 
        .ZN(n116314) );
  OAI22_X1 U86278 ( .A1(n114227), .A2(n120114), .B1(n90089), .B2(n120108), 
        .ZN(n116286) );
  OAI22_X1 U86279 ( .A1(n114226), .A2(n120114), .B1(n90088), .B2(n120108), 
        .ZN(n116258) );
  OAI22_X1 U86280 ( .A1(n114225), .A2(n120114), .B1(n90087), .B2(n120108), 
        .ZN(n116230) );
  OAI22_X1 U86281 ( .A1(n114224), .A2(n120114), .B1(n90086), .B2(n120108), 
        .ZN(n116202) );
  OAI22_X1 U86282 ( .A1(n114223), .A2(n120114), .B1(n90085), .B2(n120108), 
        .ZN(n116174) );
  OAI22_X1 U86283 ( .A1(n114222), .A2(n120114), .B1(n90084), .B2(n120108), 
        .ZN(n116146) );
  OAI22_X1 U86284 ( .A1(n114221), .A2(n120115), .B1(n90083), .B2(n120109), 
        .ZN(n116118) );
  OAI22_X1 U86285 ( .A1(n114220), .A2(n120115), .B1(n90082), .B2(n120109), 
        .ZN(n116090) );
  OAI22_X1 U86286 ( .A1(n114219), .A2(n120115), .B1(n90081), .B2(n120109), 
        .ZN(n116062) );
  OAI22_X1 U86287 ( .A1(n114218), .A2(n120115), .B1(n90080), .B2(n120109), 
        .ZN(n116034) );
  OAI22_X1 U86288 ( .A1(n114217), .A2(n120115), .B1(n90079), .B2(n120109), 
        .ZN(n116006) );
  OAI22_X1 U86289 ( .A1(n114216), .A2(n120115), .B1(n90078), .B2(n120109), 
        .ZN(n115978) );
  OAI22_X1 U86290 ( .A1(n114215), .A2(n120115), .B1(n90077), .B2(n120109), 
        .ZN(n115950) );
  OAI22_X1 U86291 ( .A1(n90557), .A2(n120115), .B1(n90076), .B2(n120109), .ZN(
        n115922) );
  OAI22_X1 U86292 ( .A1(n90556), .A2(n120115), .B1(n90075), .B2(n120109), .ZN(
        n115894) );
  OAI22_X1 U86293 ( .A1(n90555), .A2(n120115), .B1(n90074), .B2(n120109), .ZN(
        n115866) );
  OAI22_X1 U86294 ( .A1(n90554), .A2(n120115), .B1(n90073), .B2(n120109), .ZN(
        n115838) );
  OAI22_X1 U86295 ( .A1(n90553), .A2(n120115), .B1(n90072), .B2(n120109), .ZN(
        n115810) );
  OAI22_X1 U86296 ( .A1(n90552), .A2(n120116), .B1(n90071), .B2(n120110), .ZN(
        n115782) );
  OAI22_X1 U86297 ( .A1(n90551), .A2(n120116), .B1(n90070), .B2(n120110), .ZN(
        n115754) );
  OAI22_X1 U86298 ( .A1(n90550), .A2(n120116), .B1(n90069), .B2(n120110), .ZN(
        n115726) );
  OAI22_X1 U86299 ( .A1(n90549), .A2(n120116), .B1(n90068), .B2(n120110), .ZN(
        n115698) );
  OAI22_X1 U86300 ( .A1(n90548), .A2(n120116), .B1(n90067), .B2(n120110), .ZN(
        n115670) );
  OAI22_X1 U86301 ( .A1(n90547), .A2(n120116), .B1(n90066), .B2(n120110), .ZN(
        n115642) );
  OAI22_X1 U86302 ( .A1(n90546), .A2(n120116), .B1(n90065), .B2(n120110), .ZN(
        n115614) );
  OAI22_X1 U86303 ( .A1(n90545), .A2(n120116), .B1(n90064), .B2(n120110), .ZN(
        n115586) );
  OAI22_X1 U86304 ( .A1(n90544), .A2(n120116), .B1(n90063), .B2(n120110), .ZN(
        n115558) );
  OAI22_X1 U86305 ( .A1(n90543), .A2(n120116), .B1(n90062), .B2(n120110), .ZN(
        n115530) );
  OAI22_X1 U86306 ( .A1(n90542), .A2(n120116), .B1(n90061), .B2(n120110), .ZN(
        n115502) );
  OAI22_X1 U86307 ( .A1(n90541), .A2(n120116), .B1(n90060), .B2(n120110), .ZN(
        n115474) );
  OAI22_X1 U86308 ( .A1(n90540), .A2(n120117), .B1(n90059), .B2(n120111), .ZN(
        n115446) );
  OAI22_X1 U86309 ( .A1(n90539), .A2(n120117), .B1(n90058), .B2(n120111), .ZN(
        n115418) );
  OAI22_X1 U86310 ( .A1(n90538), .A2(n120117), .B1(n90057), .B2(n120111), .ZN(
        n115390) );
  OAI22_X1 U86311 ( .A1(n90537), .A2(n120117), .B1(n90056), .B2(n120111), .ZN(
        n115362) );
  OAI22_X1 U86312 ( .A1(n90536), .A2(n120117), .B1(n90055), .B2(n120111), .ZN(
        n115334) );
  OAI22_X1 U86313 ( .A1(n90535), .A2(n120117), .B1(n90054), .B2(n120111), .ZN(
        n115306) );
  OAI22_X1 U86314 ( .A1(n90534), .A2(n120117), .B1(n90053), .B2(n120111), .ZN(
        n115278) );
  OAI22_X1 U86315 ( .A1(n90533), .A2(n120117), .B1(n90052), .B2(n120111), .ZN(
        n115250) );
  OAI22_X1 U86316 ( .A1(n90532), .A2(n120117), .B1(n90051), .B2(n120111), .ZN(
        n115222) );
  OAI22_X1 U86317 ( .A1(n90531), .A2(n120117), .B1(n90050), .B2(n120111), .ZN(
        n115194) );
  OAI22_X1 U86318 ( .A1(n90324), .A2(n120129), .B1(n114253), .B2(n120123), 
        .ZN(n115167) );
  OAI22_X1 U86319 ( .A1(n90323), .A2(n120129), .B1(n114252), .B2(n120123), 
        .ZN(n115139) );
  OAI22_X1 U86320 ( .A1(n90322), .A2(n120130), .B1(n114251), .B2(n120124), 
        .ZN(n115111) );
  OAI22_X1 U86321 ( .A1(n90321), .A2(n120130), .B1(n114250), .B2(n120124), 
        .ZN(n115083) );
  OAI22_X1 U86322 ( .A1(n90320), .A2(n120130), .B1(n114249), .B2(n120124), 
        .ZN(n115055) );
  OAI22_X1 U86323 ( .A1(n90319), .A2(n120130), .B1(n114248), .B2(n120124), 
        .ZN(n115027) );
  OAI22_X1 U86324 ( .A1(n90318), .A2(n120130), .B1(n114247), .B2(n120124), 
        .ZN(n114999) );
  OAI22_X1 U86325 ( .A1(n90317), .A2(n120130), .B1(n114246), .B2(n120124), 
        .ZN(n114971) );
  OAI22_X1 U86326 ( .A1(n90316), .A2(n120130), .B1(n114245), .B2(n120124), 
        .ZN(n114943) );
  OAI22_X1 U86327 ( .A1(n90315), .A2(n120130), .B1(n114244), .B2(n120124), 
        .ZN(n114915) );
  OAI22_X1 U86328 ( .A1(n90314), .A2(n120130), .B1(n114243), .B2(n120124), 
        .ZN(n114887) );
  OAI22_X1 U86329 ( .A1(n90313), .A2(n120130), .B1(n114242), .B2(n120124), 
        .ZN(n114859) );
  OAI22_X1 U86330 ( .A1(n90312), .A2(n120130), .B1(n114241), .B2(n120124), 
        .ZN(n114831) );
  OAI22_X1 U86331 ( .A1(n90311), .A2(n120130), .B1(n114240), .B2(n120124), 
        .ZN(n114803) );
  OAI22_X1 U86332 ( .A1(n90370), .A2(n120126), .B1(n114299), .B2(n120120), 
        .ZN(n116467) );
  OAI22_X1 U86333 ( .A1(n90369), .A2(n120126), .B1(n114298), .B2(n120120), 
        .ZN(n116427) );
  OAI22_X1 U86334 ( .A1(n90368), .A2(n120126), .B1(n114297), .B2(n120120), 
        .ZN(n116399) );
  OAI22_X1 U86335 ( .A1(n90367), .A2(n120126), .B1(n114296), .B2(n120120), 
        .ZN(n116371) );
  OAI22_X1 U86336 ( .A1(n90366), .A2(n120126), .B1(n114295), .B2(n120120), 
        .ZN(n116343) );
  OAI22_X1 U86337 ( .A1(n90365), .A2(n120126), .B1(n114294), .B2(n120120), 
        .ZN(n116315) );
  OAI22_X1 U86338 ( .A1(n90364), .A2(n120126), .B1(n114293), .B2(n120120), 
        .ZN(n116287) );
  OAI22_X1 U86339 ( .A1(n90363), .A2(n120126), .B1(n114292), .B2(n120120), 
        .ZN(n116259) );
  OAI22_X1 U86340 ( .A1(n90362), .A2(n120126), .B1(n114291), .B2(n120120), 
        .ZN(n116231) );
  OAI22_X1 U86341 ( .A1(n90361), .A2(n120126), .B1(n114290), .B2(n120120), 
        .ZN(n116203) );
  OAI22_X1 U86342 ( .A1(n90360), .A2(n120126), .B1(n114289), .B2(n120120), 
        .ZN(n116175) );
  OAI22_X1 U86343 ( .A1(n90359), .A2(n120126), .B1(n114288), .B2(n120120), 
        .ZN(n116147) );
  OAI22_X1 U86344 ( .A1(n90358), .A2(n120127), .B1(n114287), .B2(n120121), 
        .ZN(n116119) );
  OAI22_X1 U86345 ( .A1(n90357), .A2(n120127), .B1(n114286), .B2(n120121), 
        .ZN(n116091) );
  OAI22_X1 U86346 ( .A1(n90356), .A2(n120127), .B1(n114285), .B2(n120121), 
        .ZN(n116063) );
  OAI22_X1 U86347 ( .A1(n90355), .A2(n120127), .B1(n114284), .B2(n120121), 
        .ZN(n116035) );
  OAI22_X1 U86348 ( .A1(n90354), .A2(n120127), .B1(n114283), .B2(n120121), 
        .ZN(n116007) );
  OAI22_X1 U86349 ( .A1(n90353), .A2(n120127), .B1(n114282), .B2(n120121), 
        .ZN(n115979) );
  OAI22_X1 U86350 ( .A1(n90352), .A2(n120127), .B1(n114281), .B2(n120121), 
        .ZN(n115951) );
  OAI22_X1 U86351 ( .A1(n90351), .A2(n120127), .B1(n114280), .B2(n120121), 
        .ZN(n115923) );
  OAI22_X1 U86352 ( .A1(n90350), .A2(n120127), .B1(n114279), .B2(n120121), 
        .ZN(n115895) );
  OAI22_X1 U86353 ( .A1(n90349), .A2(n120127), .B1(n114278), .B2(n120121), 
        .ZN(n115867) );
  OAI22_X1 U86354 ( .A1(n90348), .A2(n120127), .B1(n114277), .B2(n120121), 
        .ZN(n115839) );
  OAI22_X1 U86355 ( .A1(n90347), .A2(n120127), .B1(n114276), .B2(n120121), 
        .ZN(n115811) );
  OAI22_X1 U86356 ( .A1(n90346), .A2(n120128), .B1(n114275), .B2(n120122), 
        .ZN(n115783) );
  OAI22_X1 U86357 ( .A1(n90345), .A2(n120128), .B1(n114274), .B2(n120122), 
        .ZN(n115755) );
  OAI22_X1 U86358 ( .A1(n90344), .A2(n120128), .B1(n114273), .B2(n120122), 
        .ZN(n115727) );
  OAI22_X1 U86359 ( .A1(n90343), .A2(n120128), .B1(n114272), .B2(n120122), 
        .ZN(n115699) );
  OAI22_X1 U86360 ( .A1(n90342), .A2(n120128), .B1(n114271), .B2(n120122), 
        .ZN(n115671) );
  OAI22_X1 U86361 ( .A1(n90341), .A2(n120128), .B1(n114270), .B2(n120122), 
        .ZN(n115643) );
  OAI22_X1 U86362 ( .A1(n90340), .A2(n120128), .B1(n114269), .B2(n120122), 
        .ZN(n115615) );
  OAI22_X1 U86363 ( .A1(n90339), .A2(n120128), .B1(n114268), .B2(n120122), 
        .ZN(n115587) );
  OAI22_X1 U86364 ( .A1(n90338), .A2(n120128), .B1(n114267), .B2(n120122), 
        .ZN(n115559) );
  OAI22_X1 U86365 ( .A1(n90337), .A2(n120128), .B1(n114266), .B2(n120122), 
        .ZN(n115531) );
  OAI22_X1 U86366 ( .A1(n90336), .A2(n120128), .B1(n114265), .B2(n120122), 
        .ZN(n115503) );
  OAI22_X1 U86367 ( .A1(n90335), .A2(n120128), .B1(n114264), .B2(n120122), 
        .ZN(n115475) );
  OAI22_X1 U86368 ( .A1(n90334), .A2(n120129), .B1(n114263), .B2(n120123), 
        .ZN(n115447) );
  OAI22_X1 U86369 ( .A1(n90333), .A2(n120129), .B1(n114262), .B2(n120123), 
        .ZN(n115419) );
  OAI22_X1 U86370 ( .A1(n90332), .A2(n120129), .B1(n114261), .B2(n120123), 
        .ZN(n115391) );
  OAI22_X1 U86371 ( .A1(n90331), .A2(n120129), .B1(n114260), .B2(n120123), 
        .ZN(n115363) );
  OAI22_X1 U86372 ( .A1(n90330), .A2(n120129), .B1(n114259), .B2(n120123), 
        .ZN(n115335) );
  OAI22_X1 U86373 ( .A1(n90329), .A2(n120129), .B1(n114258), .B2(n120123), 
        .ZN(n115307) );
  OAI22_X1 U86374 ( .A1(n90328), .A2(n120129), .B1(n114257), .B2(n120123), 
        .ZN(n115279) );
  OAI22_X1 U86375 ( .A1(n90327), .A2(n120129), .B1(n114256), .B2(n120123), 
        .ZN(n115251) );
  OAI22_X1 U86376 ( .A1(n90326), .A2(n120129), .B1(n114255), .B2(n120123), 
        .ZN(n115223) );
  OAI22_X1 U86377 ( .A1(n90325), .A2(n120129), .B1(n114254), .B2(n120123), 
        .ZN(n115195) );
  OAI22_X1 U86378 ( .A1(n98599), .A2(n120051), .B1(n114596), .B2(n120045), 
        .ZN(n115173) );
  OAI22_X1 U86379 ( .A1(n98598), .A2(n120051), .B1(n114595), .B2(n120045), 
        .ZN(n115145) );
  OAI22_X1 U86380 ( .A1(n98597), .A2(n120052), .B1(n114594), .B2(n120046), 
        .ZN(n115117) );
  OAI22_X1 U86381 ( .A1(n98596), .A2(n120052), .B1(n114593), .B2(n120046), 
        .ZN(n115089) );
  OAI22_X1 U86382 ( .A1(n98595), .A2(n120052), .B1(n114592), .B2(n120046), 
        .ZN(n115061) );
  OAI22_X1 U86383 ( .A1(n98594), .A2(n120052), .B1(n114591), .B2(n120046), 
        .ZN(n115033) );
  OAI22_X1 U86384 ( .A1(n98593), .A2(n120052), .B1(n114590), .B2(n120046), 
        .ZN(n115005) );
  OAI22_X1 U86385 ( .A1(n98592), .A2(n120052), .B1(n114589), .B2(n120046), 
        .ZN(n114977) );
  OAI22_X1 U86386 ( .A1(n98591), .A2(n120052), .B1(n114588), .B2(n120046), 
        .ZN(n114949) );
  OAI22_X1 U86387 ( .A1(n98590), .A2(n120052), .B1(n114587), .B2(n120046), 
        .ZN(n114921) );
  OAI22_X1 U86388 ( .A1(n98589), .A2(n120052), .B1(n114586), .B2(n120046), 
        .ZN(n114893) );
  OAI22_X1 U86389 ( .A1(n98588), .A2(n120052), .B1(n114585), .B2(n120046), 
        .ZN(n114865) );
  OAI22_X1 U86390 ( .A1(n98587), .A2(n120052), .B1(n114584), .B2(n120046), 
        .ZN(n114837) );
  OAI22_X1 U86391 ( .A1(n98586), .A2(n120052), .B1(n114583), .B2(n120046), 
        .ZN(n114809) );
  OAI22_X1 U86392 ( .A1(n98645), .A2(n120048), .B1(n114642), .B2(n120042), 
        .ZN(n116477) );
  OAI22_X1 U86393 ( .A1(n98644), .A2(n120048), .B1(n114641), .B2(n120042), 
        .ZN(n116433) );
  OAI22_X1 U86394 ( .A1(n98643), .A2(n120048), .B1(n114640), .B2(n120042), 
        .ZN(n116405) );
  OAI22_X1 U86395 ( .A1(n98642), .A2(n120048), .B1(n114639), .B2(n120042), 
        .ZN(n116377) );
  OAI22_X1 U86396 ( .A1(n98641), .A2(n120048), .B1(n114638), .B2(n120042), 
        .ZN(n116349) );
  OAI22_X1 U86397 ( .A1(n98640), .A2(n120048), .B1(n114637), .B2(n120042), 
        .ZN(n116321) );
  OAI22_X1 U86398 ( .A1(n98639), .A2(n120048), .B1(n114636), .B2(n120042), 
        .ZN(n116293) );
  OAI22_X1 U86399 ( .A1(n98638), .A2(n120048), .B1(n114635), .B2(n120042), 
        .ZN(n116265) );
  OAI22_X1 U86400 ( .A1(n98637), .A2(n120048), .B1(n114634), .B2(n120042), 
        .ZN(n116237) );
  OAI22_X1 U86401 ( .A1(n98636), .A2(n120048), .B1(n114633), .B2(n120042), 
        .ZN(n116209) );
  OAI22_X1 U86402 ( .A1(n98635), .A2(n120048), .B1(n114632), .B2(n120042), 
        .ZN(n116181) );
  OAI22_X1 U86403 ( .A1(n98634), .A2(n120048), .B1(n114631), .B2(n120042), 
        .ZN(n116153) );
  OAI22_X1 U86404 ( .A1(n98633), .A2(n120049), .B1(n114630), .B2(n120043), 
        .ZN(n116125) );
  OAI22_X1 U86405 ( .A1(n98632), .A2(n120049), .B1(n114629), .B2(n120043), 
        .ZN(n116097) );
  OAI22_X1 U86406 ( .A1(n98631), .A2(n120049), .B1(n114628), .B2(n120043), 
        .ZN(n116069) );
  OAI22_X1 U86407 ( .A1(n98630), .A2(n120049), .B1(n114627), .B2(n120043), 
        .ZN(n116041) );
  OAI22_X1 U86408 ( .A1(n98629), .A2(n120049), .B1(n114626), .B2(n120043), 
        .ZN(n116013) );
  OAI22_X1 U86409 ( .A1(n98628), .A2(n120049), .B1(n114625), .B2(n120043), 
        .ZN(n115985) );
  OAI22_X1 U86410 ( .A1(n98627), .A2(n120049), .B1(n114624), .B2(n120043), 
        .ZN(n115957) );
  OAI22_X1 U86411 ( .A1(n98626), .A2(n120049), .B1(n114623), .B2(n120043), 
        .ZN(n115929) );
  OAI22_X1 U86412 ( .A1(n98625), .A2(n120049), .B1(n114622), .B2(n120043), 
        .ZN(n115901) );
  OAI22_X1 U86413 ( .A1(n98624), .A2(n120049), .B1(n114621), .B2(n120043), 
        .ZN(n115873) );
  OAI22_X1 U86414 ( .A1(n98623), .A2(n120049), .B1(n114620), .B2(n120043), 
        .ZN(n115845) );
  OAI22_X1 U86415 ( .A1(n98622), .A2(n120049), .B1(n114619), .B2(n120043), 
        .ZN(n115817) );
  OAI22_X1 U86416 ( .A1(n98621), .A2(n120050), .B1(n114618), .B2(n120044), 
        .ZN(n115789) );
  OAI22_X1 U86417 ( .A1(n98620), .A2(n120050), .B1(n114617), .B2(n120044), 
        .ZN(n115761) );
  OAI22_X1 U86418 ( .A1(n98619), .A2(n120050), .B1(n114616), .B2(n120044), 
        .ZN(n115733) );
  OAI22_X1 U86419 ( .A1(n98618), .A2(n120050), .B1(n114615), .B2(n120044), 
        .ZN(n115705) );
  OAI22_X1 U86420 ( .A1(n98617), .A2(n120050), .B1(n114614), .B2(n120044), 
        .ZN(n115677) );
  OAI22_X1 U86421 ( .A1(n98616), .A2(n120050), .B1(n114613), .B2(n120044), 
        .ZN(n115649) );
  OAI22_X1 U86422 ( .A1(n98615), .A2(n120050), .B1(n114612), .B2(n120044), 
        .ZN(n115621) );
  OAI22_X1 U86423 ( .A1(n98614), .A2(n120050), .B1(n114611), .B2(n120044), 
        .ZN(n115593) );
  OAI22_X1 U86424 ( .A1(n98613), .A2(n120050), .B1(n114610), .B2(n120044), 
        .ZN(n115565) );
  OAI22_X1 U86425 ( .A1(n98612), .A2(n120050), .B1(n114609), .B2(n120044), 
        .ZN(n115537) );
  OAI22_X1 U86426 ( .A1(n98611), .A2(n120050), .B1(n114608), .B2(n120044), 
        .ZN(n115509) );
  OAI22_X1 U86427 ( .A1(n98610), .A2(n120050), .B1(n114607), .B2(n120044), 
        .ZN(n115481) );
  OAI22_X1 U86428 ( .A1(n98609), .A2(n120051), .B1(n114606), .B2(n120045), 
        .ZN(n115453) );
  OAI22_X1 U86429 ( .A1(n98608), .A2(n120051), .B1(n114605), .B2(n120045), 
        .ZN(n115425) );
  OAI22_X1 U86430 ( .A1(n98607), .A2(n120051), .B1(n114604), .B2(n120045), 
        .ZN(n115397) );
  OAI22_X1 U86431 ( .A1(n98606), .A2(n120051), .B1(n114603), .B2(n120045), 
        .ZN(n115369) );
  OAI22_X1 U86432 ( .A1(n98605), .A2(n120051), .B1(n114602), .B2(n120045), 
        .ZN(n115341) );
  OAI22_X1 U86433 ( .A1(n98604), .A2(n120051), .B1(n114601), .B2(n120045), 
        .ZN(n115313) );
  OAI22_X1 U86434 ( .A1(n98603), .A2(n120051), .B1(n114600), .B2(n120045), 
        .ZN(n115285) );
  OAI22_X1 U86435 ( .A1(n98602), .A2(n120051), .B1(n114599), .B2(n120045), 
        .ZN(n115257) );
  OAI22_X1 U86436 ( .A1(n98601), .A2(n120051), .B1(n114598), .B2(n120045), 
        .ZN(n115229) );
  OAI22_X1 U86437 ( .A1(n98600), .A2(n120051), .B1(n114597), .B2(n120045), 
        .ZN(n115201) );
  OAI22_X1 U86438 ( .A1(n89500), .A2(n120829), .B1(n120826), .B2(n120809), 
        .ZN(n7483) );
  OAI22_X1 U86439 ( .A1(n89498), .A2(n120829), .B1(n120826), .B2(n120812), 
        .ZN(n7484) );
  OAI22_X1 U86440 ( .A1(n89496), .A2(n120829), .B1(n120826), .B2(n120815), 
        .ZN(n7485) );
  OAI22_X1 U86441 ( .A1(n89493), .A2(n120829), .B1(n120826), .B2(n120818), 
        .ZN(n7486) );
  OAI22_X1 U86442 ( .A1(n120622), .A2(n113900), .B1(n120809), .B2(n120616), 
        .ZN(n7419) );
  OAI22_X1 U86443 ( .A1(n120622), .A2(n113899), .B1(n120812), .B2(n120616), 
        .ZN(n7420) );
  OAI22_X1 U86444 ( .A1(n120622), .A2(n113898), .B1(n120815), .B2(n120616), 
        .ZN(n7421) );
  OAI22_X1 U86445 ( .A1(n120622), .A2(n113896), .B1(n120818), .B2(n120616), 
        .ZN(n7422) );
  OAI22_X1 U86446 ( .A1(n99183), .A2(n120475), .B1(n120810), .B2(n120469), 
        .ZN(n6651) );
  OAI22_X1 U86447 ( .A1(n99182), .A2(n120475), .B1(n120813), .B2(n120469), 
        .ZN(n6652) );
  OAI22_X1 U86448 ( .A1(n99181), .A2(n120475), .B1(n120816), .B2(n120469), 
        .ZN(n6653) );
  OAI22_X1 U86449 ( .A1(n99179), .A2(n120475), .B1(n120819), .B2(n120469), 
        .ZN(n6654) );
  OAI22_X1 U86450 ( .A1(n99315), .A2(n120451), .B1(n120810), .B2(n120445), 
        .ZN(n6523) );
  OAI22_X1 U86451 ( .A1(n99314), .A2(n120451), .B1(n120813), .B2(n120445), 
        .ZN(n6524) );
  OAI22_X1 U86452 ( .A1(n99313), .A2(n120451), .B1(n120816), .B2(n120445), 
        .ZN(n6525) );
  OAI22_X1 U86453 ( .A1(n99311), .A2(n120451), .B1(n120819), .B2(n120445), 
        .ZN(n6526) );
  OAI22_X1 U86454 ( .A1(n120524), .A2(n114060), .B1(n120809), .B2(n120517), 
        .ZN(n6907) );
  OAI22_X1 U86455 ( .A1(n120524), .A2(n114059), .B1(n120812), .B2(n120517), 
        .ZN(n6908) );
  OAI22_X1 U86456 ( .A1(n120524), .A2(n114058), .B1(n120815), .B2(n120517), 
        .ZN(n6909) );
  OAI22_X1 U86457 ( .A1(n120524), .A2(n114056), .B1(n120818), .B2(n120517), 
        .ZN(n6910) );
  OAI22_X1 U86458 ( .A1(n99051), .A2(n120499), .B1(n120809), .B2(n120493), 
        .ZN(n6779) );
  OAI22_X1 U86459 ( .A1(n99050), .A2(n120499), .B1(n120812), .B2(n120493), 
        .ZN(n6780) );
  OAI22_X1 U86460 ( .A1(n99049), .A2(n120499), .B1(n120815), .B2(n120493), 
        .ZN(n6781) );
  OAI22_X1 U86461 ( .A1(n99047), .A2(n120499), .B1(n120818), .B2(n120493), 
        .ZN(n6782) );
  OAI22_X1 U86462 ( .A1(n99117), .A2(n120487), .B1(n120810), .B2(n120481), 
        .ZN(n6715) );
  OAI22_X1 U86463 ( .A1(n99116), .A2(n120487), .B1(n120813), .B2(n120481), 
        .ZN(n6716) );
  OAI22_X1 U86464 ( .A1(n99115), .A2(n120487), .B1(n120816), .B2(n120481), 
        .ZN(n6717) );
  OAI22_X1 U86465 ( .A1(n99113), .A2(n120487), .B1(n120819), .B2(n120481), 
        .ZN(n6718) );
  OAI22_X1 U86466 ( .A1(n99249), .A2(n120463), .B1(n120810), .B2(n120457), 
        .ZN(n6587) );
  OAI22_X1 U86467 ( .A1(n99248), .A2(n120463), .B1(n120813), .B2(n120457), 
        .ZN(n6588) );
  OAI22_X1 U86468 ( .A1(n99247), .A2(n120463), .B1(n120816), .B2(n120457), 
        .ZN(n6589) );
  OAI22_X1 U86469 ( .A1(n99245), .A2(n120463), .B1(n120819), .B2(n120457), 
        .ZN(n6590) );
  OAI22_X1 U86470 ( .A1(n98718), .A2(n120586), .B1(n120809), .B2(n120580), 
        .ZN(n7227) );
  OAI22_X1 U86471 ( .A1(n98717), .A2(n120586), .B1(n120812), .B2(n120580), 
        .ZN(n7228) );
  OAI22_X1 U86472 ( .A1(n98716), .A2(n120586), .B1(n120815), .B2(n120580), 
        .ZN(n7229) );
  OAI22_X1 U86473 ( .A1(n98714), .A2(n120586), .B1(n120818), .B2(n120580), 
        .ZN(n7230) );
  OAI22_X1 U86474 ( .A1(n98652), .A2(n120598), .B1(n120809), .B2(n120592), 
        .ZN(n7291) );
  OAI22_X1 U86475 ( .A1(n98651), .A2(n120598), .B1(n120812), .B2(n120592), 
        .ZN(n7292) );
  OAI22_X1 U86476 ( .A1(n98650), .A2(n120598), .B1(n120815), .B2(n120592), 
        .ZN(n7293) );
  OAI22_X1 U86477 ( .A1(n98648), .A2(n120598), .B1(n120818), .B2(n120592), 
        .ZN(n7294) );
  OAI22_X1 U86478 ( .A1(n99584), .A2(n120365), .B1(n120810), .B2(n120359), 
        .ZN(n6075) );
  OAI22_X1 U86479 ( .A1(n99583), .A2(n120365), .B1(n120813), .B2(n120359), 
        .ZN(n6076) );
  OAI22_X1 U86480 ( .A1(n99582), .A2(n120365), .B1(n120816), .B2(n120359), 
        .ZN(n6077) );
  OAI22_X1 U86481 ( .A1(n99580), .A2(n120365), .B1(n120819), .B2(n120359), 
        .ZN(n6078) );
  OAI22_X1 U86482 ( .A1(n120341), .A2(n114310), .B1(n120810), .B2(n120334), 
        .ZN(n5947) );
  OAI22_X1 U86483 ( .A1(n120341), .A2(n114309), .B1(n120813), .B2(n120334), 
        .ZN(n5948) );
  OAI22_X1 U86484 ( .A1(n120341), .A2(n114308), .B1(n120816), .B2(n120334), 
        .ZN(n5949) );
  OAI22_X1 U86485 ( .A1(n120341), .A2(n114306), .B1(n120819), .B2(n120334), 
        .ZN(n5950) );
  OAI22_X1 U86486 ( .A1(n99450), .A2(n120402), .B1(n120810), .B2(n120396), 
        .ZN(n6267) );
  OAI22_X1 U86487 ( .A1(n99449), .A2(n120402), .B1(n120813), .B2(n120396), 
        .ZN(n6268) );
  OAI22_X1 U86488 ( .A1(n99448), .A2(n120402), .B1(n120816), .B2(n120396), 
        .ZN(n6269) );
  OAI22_X1 U86489 ( .A1(n99446), .A2(n120402), .B1(n120819), .B2(n120396), 
        .ZN(n6270) );
  OAI22_X1 U86490 ( .A1(n99720), .A2(n120328), .B1(n120811), .B2(n120322), 
        .ZN(n5883) );
  OAI22_X1 U86491 ( .A1(n99719), .A2(n120328), .B1(n120814), .B2(n120322), 
        .ZN(n5884) );
  OAI22_X1 U86492 ( .A1(n99718), .A2(n120328), .B1(n120817), .B2(n120322), 
        .ZN(n5885) );
  OAI22_X1 U86493 ( .A1(n99716), .A2(n120328), .B1(n120820), .B2(n120322), 
        .ZN(n5886) );
  OAI22_X1 U86494 ( .A1(n99918), .A2(n120277), .B1(n120811), .B2(n120271), 
        .ZN(n5627) );
  OAI22_X1 U86495 ( .A1(n99917), .A2(n120277), .B1(n120814), .B2(n120271), 
        .ZN(n5628) );
  OAI22_X1 U86496 ( .A1(n99916), .A2(n120277), .B1(n120817), .B2(n120271), 
        .ZN(n5629) );
  OAI22_X1 U86497 ( .A1(n99914), .A2(n120277), .B1(n120820), .B2(n120271), 
        .ZN(n5630) );
  OAI22_X1 U86498 ( .A1(n90035), .A2(n120536), .B1(n120809), .B2(n120530), 
        .ZN(n6971) );
  OAI22_X1 U86499 ( .A1(n90034), .A2(n120536), .B1(n120812), .B2(n120530), 
        .ZN(n6972) );
  OAI22_X1 U86500 ( .A1(n90033), .A2(n120536), .B1(n120815), .B2(n120530), 
        .ZN(n6973) );
  OAI22_X1 U86501 ( .A1(n90031), .A2(n120536), .B1(n120818), .B2(n120530), 
        .ZN(n6974) );
  OAI22_X1 U86502 ( .A1(n89969), .A2(n120545), .B1(n120809), .B2(n120542), 
        .ZN(n7035) );
  OAI22_X1 U86503 ( .A1(n89968), .A2(n120545), .B1(n120812), .B2(n120542), 
        .ZN(n7036) );
  OAI22_X1 U86504 ( .A1(n89967), .A2(n120545), .B1(n120815), .B2(n120542), 
        .ZN(n7037) );
  OAI22_X1 U86505 ( .A1(n89965), .A2(n120545), .B1(n120818), .B2(n120542), 
        .ZN(n7038) );
  OAI22_X1 U86506 ( .A1(n90516), .A2(n120385), .B1(n120810), .B2(n120384), 
        .ZN(n6203) );
  OAI22_X1 U86507 ( .A1(n90515), .A2(n120385), .B1(n120813), .B2(n120384), 
        .ZN(n6204) );
  OAI22_X1 U86508 ( .A1(n90514), .A2(n120385), .B1(n120816), .B2(n120384), 
        .ZN(n6205) );
  OAI22_X1 U86509 ( .A1(n90512), .A2(n120387), .B1(n120819), .B2(n120384), 
        .ZN(n6206) );
  OAI22_X1 U86510 ( .A1(n90310), .A2(n120439), .B1(n120810), .B2(n120433), 
        .ZN(n6459) );
  OAI22_X1 U86511 ( .A1(n90309), .A2(n120439), .B1(n120813), .B2(n120433), 
        .ZN(n6460) );
  OAI22_X1 U86512 ( .A1(n90308), .A2(n120439), .B1(n120816), .B2(n120433), 
        .ZN(n6461) );
  OAI22_X1 U86513 ( .A1(n90306), .A2(n120439), .B1(n120819), .B2(n120433), 
        .ZN(n6462) );
  OAI22_X1 U86514 ( .A1(n90377), .A2(n120427), .B1(n120810), .B2(n120421), 
        .ZN(n6395) );
  OAI22_X1 U86515 ( .A1(n90376), .A2(n120427), .B1(n120813), .B2(n120421), 
        .ZN(n6396) );
  OAI22_X1 U86516 ( .A1(n90375), .A2(n120427), .B1(n120816), .B2(n120421), 
        .ZN(n6397) );
  OAI22_X1 U86517 ( .A1(n90373), .A2(n120427), .B1(n120819), .B2(n120421), 
        .ZN(n6398) );
  OAI22_X1 U86518 ( .A1(n90715), .A2(n120353), .B1(n120810), .B2(n120347), 
        .ZN(n6011) );
  OAI22_X1 U86519 ( .A1(n90714), .A2(n120353), .B1(n120813), .B2(n120347), 
        .ZN(n6012) );
  OAI22_X1 U86520 ( .A1(n90713), .A2(n120353), .B1(n120816), .B2(n120347), 
        .ZN(n6013) );
  OAI22_X1 U86521 ( .A1(n90711), .A2(n120353), .B1(n120819), .B2(n120347), 
        .ZN(n6014) );
  AOI22_X1 U86522 ( .A1(n119976), .A2(n118922), .B1(n119970), .B2(n111007), 
        .ZN(n117706) );
  AOI22_X1 U86523 ( .A1(n120024), .A2(n118862), .B1(n120022), .B2(OUT2[11]), 
        .ZN(n117701) );
  AOI22_X1 U86524 ( .A1(n119952), .A2(n118336), .B1(n119946), .B2(n118216), 
        .ZN(n117708) );
  AOI22_X1 U86525 ( .A1(n119977), .A2(n118923), .B1(n119971), .B2(n111008), 
        .ZN(n117684) );
  AOI22_X1 U86526 ( .A1(n120025), .A2(n118863), .B1(n120022), .B2(OUT2[12]), 
        .ZN(n117679) );
  AOI22_X1 U86527 ( .A1(n119953), .A2(n118337), .B1(n119947), .B2(n118217), 
        .ZN(n117686) );
  AOI22_X1 U86528 ( .A1(n119977), .A2(n118924), .B1(n119971), .B2(n111009), 
        .ZN(n117662) );
  AOI22_X1 U86529 ( .A1(n120025), .A2(n118864), .B1(n120022), .B2(OUT2[13]), 
        .ZN(n117657) );
  AOI22_X1 U86530 ( .A1(n119953), .A2(n118338), .B1(n119947), .B2(n118218), 
        .ZN(n117664) );
  AOI22_X1 U86531 ( .A1(n119977), .A2(n118925), .B1(n119971), .B2(n111010), 
        .ZN(n117640) );
  AOI22_X1 U86532 ( .A1(n120025), .A2(n118865), .B1(n120022), .B2(OUT2[14]), 
        .ZN(n117635) );
  AOI22_X1 U86533 ( .A1(n119953), .A2(n118339), .B1(n119947), .B2(n118219), 
        .ZN(n117642) );
  AOI22_X1 U86534 ( .A1(n119977), .A2(n118926), .B1(n119971), .B2(n111011), 
        .ZN(n117618) );
  AOI22_X1 U86535 ( .A1(n120025), .A2(n118866), .B1(n120022), .B2(OUT2[15]), 
        .ZN(n117613) );
  AOI22_X1 U86536 ( .A1(n119953), .A2(n118340), .B1(n119947), .B2(n118220), 
        .ZN(n117620) );
  AOI22_X1 U86537 ( .A1(n119977), .A2(n118927), .B1(n119971), .B2(n111012), 
        .ZN(n117596) );
  AOI22_X1 U86538 ( .A1(n120025), .A2(n118867), .B1(n120022), .B2(OUT2[16]), 
        .ZN(n117591) );
  AOI22_X1 U86539 ( .A1(n119953), .A2(n118341), .B1(n119947), .B2(n118221), 
        .ZN(n117598) );
  AOI22_X1 U86540 ( .A1(n119977), .A2(n118928), .B1(n119971), .B2(n111013), 
        .ZN(n117574) );
  AOI22_X1 U86541 ( .A1(n120025), .A2(n118868), .B1(n120021), .B2(OUT2[17]), 
        .ZN(n117569) );
  AOI22_X1 U86542 ( .A1(n119953), .A2(n118342), .B1(n119947), .B2(n118222), 
        .ZN(n117576) );
  AOI22_X1 U86543 ( .A1(n119977), .A2(n118929), .B1(n119971), .B2(n111014), 
        .ZN(n117552) );
  AOI22_X1 U86544 ( .A1(n120025), .A2(n118869), .B1(n120021), .B2(OUT2[18]), 
        .ZN(n117547) );
  AOI22_X1 U86545 ( .A1(n119953), .A2(n118343), .B1(n119947), .B2(n118223), 
        .ZN(n117554) );
  AOI22_X1 U86546 ( .A1(n119977), .A2(n118930), .B1(n119971), .B2(n111015), 
        .ZN(n117529) );
  AOI22_X1 U86547 ( .A1(n120025), .A2(n118870), .B1(n120021), .B2(OUT2[19]), 
        .ZN(n117524) );
  AOI22_X1 U86548 ( .A1(n119953), .A2(n118344), .B1(n119947), .B2(n118224), 
        .ZN(n117531) );
  AOI22_X1 U86549 ( .A1(n119977), .A2(n118931), .B1(n119971), .B2(n111016), 
        .ZN(n117506) );
  AOI22_X1 U86550 ( .A1(n120025), .A2(n118871), .B1(n120021), .B2(OUT2[20]), 
        .ZN(n117501) );
  AOI22_X1 U86551 ( .A1(n119953), .A2(n118345), .B1(n119947), .B2(n118225), 
        .ZN(n117508) );
  AOI22_X1 U86552 ( .A1(n119977), .A2(n118932), .B1(n119971), .B2(n111017), 
        .ZN(n117483) );
  AOI22_X1 U86553 ( .A1(n120025), .A2(n118872), .B1(n120021), .B2(OUT2[21]), 
        .ZN(n117478) );
  AOI22_X1 U86554 ( .A1(n119953), .A2(n118346), .B1(n119947), .B2(n118226), 
        .ZN(n117485) );
  AOI22_X1 U86555 ( .A1(n119977), .A2(n118933), .B1(n119971), .B2(n111018), 
        .ZN(n117460) );
  AOI22_X1 U86556 ( .A1(n120025), .A2(n118873), .B1(n120021), .B2(OUT2[22]), 
        .ZN(n117455) );
  AOI22_X1 U86557 ( .A1(n119953), .A2(n118347), .B1(n119947), .B2(n118227), 
        .ZN(n117462) );
  AOI22_X1 U86558 ( .A1(n119977), .A2(n118934), .B1(n119971), .B2(n111019), 
        .ZN(n117437) );
  AOI22_X1 U86559 ( .A1(n120025), .A2(n118874), .B1(n120021), .B2(OUT2[23]), 
        .ZN(n117432) );
  AOI22_X1 U86560 ( .A1(n119953), .A2(n118348), .B1(n119947), .B2(n118228), 
        .ZN(n117439) );
  AOI22_X1 U86561 ( .A1(n119978), .A2(n118935), .B1(n119972), .B2(n111020), 
        .ZN(n117414) );
  AOI22_X1 U86562 ( .A1(n120026), .A2(n118875), .B1(n120021), .B2(OUT2[24]), 
        .ZN(n117409) );
  AOI22_X1 U86563 ( .A1(n119954), .A2(n118349), .B1(n119948), .B2(n118229), 
        .ZN(n117416) );
  AOI22_X1 U86564 ( .A1(n119978), .A2(n118936), .B1(n119972), .B2(n111021), 
        .ZN(n117391) );
  AOI22_X1 U86565 ( .A1(n120026), .A2(n118876), .B1(n120021), .B2(OUT2[25]), 
        .ZN(n117386) );
  AOI22_X1 U86566 ( .A1(n119954), .A2(n118350), .B1(n119948), .B2(n118230), 
        .ZN(n117393) );
  AOI22_X1 U86567 ( .A1(n119978), .A2(n118937), .B1(n119972), .B2(n111022), 
        .ZN(n117368) );
  AOI22_X1 U86568 ( .A1(n120026), .A2(n118877), .B1(n120021), .B2(OUT2[26]), 
        .ZN(n117363) );
  AOI22_X1 U86569 ( .A1(n119954), .A2(n118351), .B1(n119948), .B2(n118231), 
        .ZN(n117370) );
  AOI22_X1 U86570 ( .A1(n119978), .A2(n118938), .B1(n119972), .B2(n111023), 
        .ZN(n117345) );
  AOI22_X1 U86571 ( .A1(n120026), .A2(n118878), .B1(n120021), .B2(OUT2[27]), 
        .ZN(n117340) );
  AOI22_X1 U86572 ( .A1(n119954), .A2(n118352), .B1(n119948), .B2(n118232), 
        .ZN(n117347) );
  AOI22_X1 U86573 ( .A1(n119978), .A2(n118939), .B1(n119972), .B2(n111024), 
        .ZN(n117322) );
  AOI22_X1 U86574 ( .A1(n120026), .A2(n118879), .B1(n120021), .B2(OUT2[28]), 
        .ZN(n117317) );
  AOI22_X1 U86575 ( .A1(n119954), .A2(n118353), .B1(n119948), .B2(n118233), 
        .ZN(n117324) );
  AOI22_X1 U86576 ( .A1(n119978), .A2(n118940), .B1(n119972), .B2(n111025), 
        .ZN(n117299) );
  AOI22_X1 U86577 ( .A1(n120026), .A2(n118880), .B1(n120021), .B2(OUT2[29]), 
        .ZN(n117294) );
  AOI22_X1 U86578 ( .A1(n119954), .A2(n118354), .B1(n119948), .B2(n118234), 
        .ZN(n117301) );
  AOI22_X1 U86579 ( .A1(n119978), .A2(n118941), .B1(n119972), .B2(n111026), 
        .ZN(n117276) );
  AOI22_X1 U86580 ( .A1(n120026), .A2(n118881), .B1(n120020), .B2(OUT2[30]), 
        .ZN(n117271) );
  AOI22_X1 U86581 ( .A1(n119954), .A2(n118355), .B1(n119948), .B2(n118235), 
        .ZN(n117278) );
  AOI22_X1 U86582 ( .A1(n119978), .A2(n118942), .B1(n119972), .B2(n111027), 
        .ZN(n117253) );
  AOI22_X1 U86583 ( .A1(n120026), .A2(n118882), .B1(n120020), .B2(OUT2[31]), 
        .ZN(n117248) );
  AOI22_X1 U86584 ( .A1(n119954), .A2(n118356), .B1(n119948), .B2(n118236), 
        .ZN(n117255) );
  AOI22_X1 U86585 ( .A1(n119978), .A2(n118943), .B1(n119972), .B2(n111028), 
        .ZN(n117230) );
  AOI22_X1 U86586 ( .A1(n120026), .A2(n118883), .B1(n120020), .B2(OUT2[32]), 
        .ZN(n117225) );
  AOI22_X1 U86587 ( .A1(n119954), .A2(n118357), .B1(n119948), .B2(n118237), 
        .ZN(n117232) );
  AOI22_X1 U86588 ( .A1(n119978), .A2(n118944), .B1(n119972), .B2(n111029), 
        .ZN(n117207) );
  AOI22_X1 U86589 ( .A1(n120026), .A2(n118884), .B1(n120020), .B2(OUT2[33]), 
        .ZN(n117202) );
  AOI22_X1 U86590 ( .A1(n119954), .A2(n118358), .B1(n119948), .B2(n118238), 
        .ZN(n117209) );
  AOI22_X1 U86591 ( .A1(n119978), .A2(n118945), .B1(n119972), .B2(n111030), 
        .ZN(n117184) );
  AOI22_X1 U86592 ( .A1(n120026), .A2(n118885), .B1(n120020), .B2(OUT2[34]), 
        .ZN(n117179) );
  AOI22_X1 U86593 ( .A1(n119954), .A2(n118359), .B1(n119948), .B2(n118239), 
        .ZN(n117186) );
  AOI22_X1 U86594 ( .A1(n119978), .A2(n118946), .B1(n119972), .B2(n111031), 
        .ZN(n117161) );
  AOI22_X1 U86595 ( .A1(n120026), .A2(n118886), .B1(n120020), .B2(OUT2[35]), 
        .ZN(n117156) );
  AOI22_X1 U86596 ( .A1(n119954), .A2(n118360), .B1(n119948), .B2(n118240), 
        .ZN(n117163) );
  AOI22_X1 U86597 ( .A1(n119979), .A2(n118947), .B1(n119973), .B2(n111032), 
        .ZN(n117138) );
  AOI22_X1 U86598 ( .A1(n120027), .A2(n118887), .B1(n120020), .B2(OUT2[36]), 
        .ZN(n117133) );
  AOI22_X1 U86599 ( .A1(n119955), .A2(n118361), .B1(n119949), .B2(n118241), 
        .ZN(n117140) );
  AOI22_X1 U86600 ( .A1(n119979), .A2(n118948), .B1(n119973), .B2(n111033), 
        .ZN(n117115) );
  AOI22_X1 U86601 ( .A1(n120027), .A2(n118888), .B1(n120020), .B2(OUT2[37]), 
        .ZN(n117110) );
  AOI22_X1 U86602 ( .A1(n119955), .A2(n118362), .B1(n119949), .B2(n118242), 
        .ZN(n117117) );
  AOI22_X1 U86603 ( .A1(n119979), .A2(n118949), .B1(n119973), .B2(n111034), 
        .ZN(n117092) );
  AOI22_X1 U86604 ( .A1(n120027), .A2(n118889), .B1(n120020), .B2(OUT2[38]), 
        .ZN(n117087) );
  AOI22_X1 U86605 ( .A1(n119955), .A2(n118363), .B1(n119949), .B2(n118243), 
        .ZN(n117094) );
  AOI22_X1 U86606 ( .A1(n119979), .A2(n118950), .B1(n119973), .B2(n111035), 
        .ZN(n117069) );
  AOI22_X1 U86607 ( .A1(n120027), .A2(n118890), .B1(n120020), .B2(OUT2[39]), 
        .ZN(n117064) );
  AOI22_X1 U86608 ( .A1(n119955), .A2(n118364), .B1(n119949), .B2(n118244), 
        .ZN(n117071) );
  AOI22_X1 U86609 ( .A1(n119979), .A2(n118951), .B1(n119973), .B2(n111036), 
        .ZN(n117046) );
  AOI22_X1 U86610 ( .A1(n120027), .A2(n118891), .B1(n120020), .B2(OUT2[40]), 
        .ZN(n117041) );
  AOI22_X1 U86611 ( .A1(n119955), .A2(n118365), .B1(n119949), .B2(n118245), 
        .ZN(n117048) );
  AOI22_X1 U86612 ( .A1(n119979), .A2(n118952), .B1(n119973), .B2(n111037), 
        .ZN(n117023) );
  AOI22_X1 U86613 ( .A1(n120027), .A2(n118892), .B1(n120020), .B2(OUT2[41]), 
        .ZN(n117018) );
  AOI22_X1 U86614 ( .A1(n119955), .A2(n118366), .B1(n119949), .B2(n118246), 
        .ZN(n117025) );
  AOI22_X1 U86615 ( .A1(n119979), .A2(n118953), .B1(n119973), .B2(n111038), 
        .ZN(n117000) );
  AOI22_X1 U86616 ( .A1(n120027), .A2(n118893), .B1(n120019), .B2(OUT2[42]), 
        .ZN(n116995) );
  AOI22_X1 U86617 ( .A1(n119955), .A2(n118367), .B1(n119949), .B2(n118247), 
        .ZN(n117002) );
  AOI22_X1 U86618 ( .A1(n119979), .A2(n118954), .B1(n119973), .B2(n111039), 
        .ZN(n116977) );
  AOI22_X1 U86619 ( .A1(n120027), .A2(n118894), .B1(n120019), .B2(OUT2[43]), 
        .ZN(n116972) );
  AOI22_X1 U86620 ( .A1(n119955), .A2(n118368), .B1(n119949), .B2(n118248), 
        .ZN(n116979) );
  AOI22_X1 U86621 ( .A1(n119979), .A2(n118955), .B1(n119973), .B2(n111040), 
        .ZN(n116954) );
  AOI22_X1 U86622 ( .A1(n120027), .A2(n118895), .B1(n120019), .B2(OUT2[44]), 
        .ZN(n116949) );
  AOI22_X1 U86623 ( .A1(n119955), .A2(n118369), .B1(n119949), .B2(n118249), 
        .ZN(n116956) );
  AOI22_X1 U86624 ( .A1(n119979), .A2(n118956), .B1(n119973), .B2(n118070), 
        .ZN(n116931) );
  AOI22_X1 U86625 ( .A1(n120027), .A2(n118896), .B1(n120019), .B2(OUT2[45]), 
        .ZN(n116926) );
  AOI22_X1 U86626 ( .A1(n119955), .A2(n118370), .B1(n119949), .B2(n118250), 
        .ZN(n116933) );
  AOI22_X1 U86627 ( .A1(n119979), .A2(n118957), .B1(n119973), .B2(n118071), 
        .ZN(n116908) );
  AOI22_X1 U86628 ( .A1(n120027), .A2(n118897), .B1(n120019), .B2(OUT2[46]), 
        .ZN(n116903) );
  AOI22_X1 U86629 ( .A1(n119955), .A2(n118371), .B1(n119949), .B2(n118251), 
        .ZN(n116910) );
  AOI22_X1 U86630 ( .A1(n119979), .A2(n118958), .B1(n119973), .B2(n118072), 
        .ZN(n116885) );
  AOI22_X1 U86631 ( .A1(n120027), .A2(n118898), .B1(n120019), .B2(OUT2[47]), 
        .ZN(n116880) );
  AOI22_X1 U86632 ( .A1(n119955), .A2(n118372), .B1(n119949), .B2(n118252), 
        .ZN(n116887) );
  AOI22_X1 U86633 ( .A1(n119980), .A2(n118959), .B1(n119974), .B2(n118073), 
        .ZN(n116862) );
  AOI22_X1 U86634 ( .A1(n120028), .A2(n118899), .B1(n120019), .B2(OUT2[48]), 
        .ZN(n116857) );
  AOI22_X1 U86635 ( .A1(n119956), .A2(n118373), .B1(n119950), .B2(n118253), 
        .ZN(n116864) );
  AOI22_X1 U86636 ( .A1(n119980), .A2(n118960), .B1(n119974), .B2(n118074), 
        .ZN(n116839) );
  AOI22_X1 U86637 ( .A1(n120028), .A2(n118900), .B1(n120019), .B2(OUT2[49]), 
        .ZN(n116834) );
  AOI22_X1 U86638 ( .A1(n119956), .A2(n118374), .B1(n119950), .B2(n118254), 
        .ZN(n116841) );
  AOI22_X1 U86639 ( .A1(n119980), .A2(n118961), .B1(n119974), .B2(n118075), 
        .ZN(n116816) );
  AOI22_X1 U86640 ( .A1(n120028), .A2(n118901), .B1(n120019), .B2(OUT2[50]), 
        .ZN(n116811) );
  AOI22_X1 U86641 ( .A1(n119956), .A2(n118375), .B1(n119950), .B2(n118255), 
        .ZN(n116818) );
  AOI22_X1 U86642 ( .A1(n119980), .A2(n118962), .B1(n119974), .B2(n118076), 
        .ZN(n116793) );
  AOI22_X1 U86643 ( .A1(n120028), .A2(n118902), .B1(n120019), .B2(OUT2[51]), 
        .ZN(n116788) );
  AOI22_X1 U86644 ( .A1(n119956), .A2(n118376), .B1(n119950), .B2(n118256), 
        .ZN(n116795) );
  AOI22_X1 U86645 ( .A1(n119980), .A2(n118963), .B1(n119974), .B2(n118077), 
        .ZN(n116770) );
  AOI22_X1 U86646 ( .A1(n120028), .A2(n118903), .B1(n120019), .B2(OUT2[52]), 
        .ZN(n116765) );
  AOI22_X1 U86647 ( .A1(n119956), .A2(n118377), .B1(n119950), .B2(n118257), 
        .ZN(n116772) );
  AOI22_X1 U86648 ( .A1(n119980), .A2(n118964), .B1(n119974), .B2(n118078), 
        .ZN(n116747) );
  AOI22_X1 U86649 ( .A1(n120028), .A2(n118904), .B1(n120019), .B2(OUT2[53]), 
        .ZN(n116742) );
  AOI22_X1 U86650 ( .A1(n119956), .A2(n118378), .B1(n119950), .B2(n118258), 
        .ZN(n116749) );
  AOI22_X1 U86651 ( .A1(n119980), .A2(n118965), .B1(n119974), .B2(n118079), 
        .ZN(n116724) );
  AOI22_X1 U86652 ( .A1(n120028), .A2(n118905), .B1(n120019), .B2(OUT2[54]), 
        .ZN(n116719) );
  AOI22_X1 U86653 ( .A1(n119956), .A2(n118379), .B1(n119950), .B2(n118259), 
        .ZN(n116726) );
  AOI22_X1 U86654 ( .A1(n119980), .A2(n118966), .B1(n119974), .B2(n118080), 
        .ZN(n116701) );
  AOI22_X1 U86655 ( .A1(n120028), .A2(n118906), .B1(n120018), .B2(OUT2[55]), 
        .ZN(n116696) );
  AOI22_X1 U86656 ( .A1(n119956), .A2(n118380), .B1(n119950), .B2(n118260), 
        .ZN(n116703) );
  AOI22_X1 U86657 ( .A1(n119980), .A2(n118967), .B1(n119974), .B2(n118081), 
        .ZN(n116678) );
  AOI22_X1 U86658 ( .A1(n120028), .A2(n118907), .B1(n120018), .B2(OUT2[56]), 
        .ZN(n116673) );
  AOI22_X1 U86659 ( .A1(n119956), .A2(n118381), .B1(n119950), .B2(n118261), 
        .ZN(n116680) );
  AOI22_X1 U86660 ( .A1(n119980), .A2(n118968), .B1(n119974), .B2(n118082), 
        .ZN(n116655) );
  AOI22_X1 U86661 ( .A1(n120028), .A2(n118908), .B1(n120018), .B2(OUT2[57]), 
        .ZN(n116650) );
  AOI22_X1 U86662 ( .A1(n119956), .A2(n118382), .B1(n119950), .B2(n118262), 
        .ZN(n116657) );
  AOI22_X1 U86663 ( .A1(n119980), .A2(n118969), .B1(n119974), .B2(n118083), 
        .ZN(n116632) );
  AOI22_X1 U86664 ( .A1(n120028), .A2(n118909), .B1(n120018), .B2(OUT2[58]), 
        .ZN(n116627) );
  AOI22_X1 U86665 ( .A1(n119956), .A2(n118383), .B1(n119950), .B2(n118263), 
        .ZN(n116634) );
  AOI22_X1 U86666 ( .A1(n119980), .A2(n118970), .B1(n119974), .B2(n118084), 
        .ZN(n116609) );
  AOI22_X1 U86667 ( .A1(n120028), .A2(n118910), .B1(n120018), .B2(OUT2[59]), 
        .ZN(n116604) );
  AOI22_X1 U86668 ( .A1(n119956), .A2(n118384), .B1(n119950), .B2(n118264), 
        .ZN(n116611) );
  AOI22_X1 U86669 ( .A1(n120225), .A2(n118532), .B1(n120217), .B2(OUT1[46]), 
        .ZN(n115155) );
  AOI22_X1 U86670 ( .A1(n120177), .A2(n118251), .B1(n120171), .B2(n119114), 
        .ZN(n115160) );
  AOI22_X1 U86671 ( .A1(n120153), .A2(n118738), .B1(n120147), .B2(n119050), 
        .ZN(n115162) );
  AOI22_X1 U86672 ( .A1(n120225), .A2(n118533), .B1(n120217), .B2(OUT1[47]), 
        .ZN(n115127) );
  AOI22_X1 U86673 ( .A1(n120177), .A2(n118252), .B1(n120171), .B2(n119115), 
        .ZN(n115132) );
  AOI22_X1 U86674 ( .A1(n120153), .A2(n118739), .B1(n120147), .B2(n119051), 
        .ZN(n115134) );
  AOI22_X1 U86675 ( .A1(n120226), .A2(n118534), .B1(n120217), .B2(OUT1[48]), 
        .ZN(n115099) );
  AOI22_X1 U86676 ( .A1(n120178), .A2(n118253), .B1(n120172), .B2(n119116), 
        .ZN(n115104) );
  AOI22_X1 U86677 ( .A1(n120154), .A2(n118740), .B1(n120148), .B2(n119052), 
        .ZN(n115106) );
  AOI22_X1 U86678 ( .A1(n120226), .A2(n118535), .B1(n120217), .B2(OUT1[49]), 
        .ZN(n115071) );
  AOI22_X1 U86679 ( .A1(n120178), .A2(n118254), .B1(n120172), .B2(n119117), 
        .ZN(n115076) );
  AOI22_X1 U86680 ( .A1(n120154), .A2(n118741), .B1(n120148), .B2(n119053), 
        .ZN(n115078) );
  AOI22_X1 U86681 ( .A1(n120226), .A2(n118536), .B1(n120217), .B2(OUT1[50]), 
        .ZN(n115043) );
  AOI22_X1 U86682 ( .A1(n120178), .A2(n118255), .B1(n120172), .B2(n119118), 
        .ZN(n115048) );
  AOI22_X1 U86683 ( .A1(n120154), .A2(n118742), .B1(n120148), .B2(n119054), 
        .ZN(n115050) );
  AOI22_X1 U86684 ( .A1(n120226), .A2(n118537), .B1(n120217), .B2(OUT1[51]), 
        .ZN(n115015) );
  AOI22_X1 U86685 ( .A1(n120178), .A2(n118256), .B1(n120172), .B2(n119119), 
        .ZN(n115020) );
  AOI22_X1 U86686 ( .A1(n120154), .A2(n118743), .B1(n120148), .B2(n119055), 
        .ZN(n115022) );
  AOI22_X1 U86687 ( .A1(n120226), .A2(n118538), .B1(n120217), .B2(OUT1[52]), 
        .ZN(n114987) );
  AOI22_X1 U86688 ( .A1(n120178), .A2(n118257), .B1(n120172), .B2(n119120), 
        .ZN(n114992) );
  AOI22_X1 U86689 ( .A1(n120154), .A2(n118744), .B1(n120148), .B2(n119056), 
        .ZN(n114994) );
  AOI22_X1 U86690 ( .A1(n120226), .A2(n118539), .B1(n120217), .B2(OUT1[53]), 
        .ZN(n114959) );
  AOI22_X1 U86691 ( .A1(n120178), .A2(n118258), .B1(n120172), .B2(n119121), 
        .ZN(n114964) );
  AOI22_X1 U86692 ( .A1(n120154), .A2(n118745), .B1(n120148), .B2(n119057), 
        .ZN(n114966) );
  AOI22_X1 U86693 ( .A1(n120226), .A2(n118540), .B1(n120217), .B2(OUT1[54]), 
        .ZN(n114931) );
  AOI22_X1 U86694 ( .A1(n120178), .A2(n118259), .B1(n120172), .B2(n119122), 
        .ZN(n114936) );
  AOI22_X1 U86695 ( .A1(n120154), .A2(n118746), .B1(n120148), .B2(n119058), 
        .ZN(n114938) );
  AOI22_X1 U86696 ( .A1(n120226), .A2(n118541), .B1(n120216), .B2(OUT1[55]), 
        .ZN(n114903) );
  AOI22_X1 U86697 ( .A1(n120178), .A2(n118260), .B1(n120172), .B2(n119123), 
        .ZN(n114908) );
  AOI22_X1 U86698 ( .A1(n120154), .A2(n118747), .B1(n120148), .B2(n119059), 
        .ZN(n114910) );
  AOI22_X1 U86699 ( .A1(n120226), .A2(n118542), .B1(n120216), .B2(OUT1[56]), 
        .ZN(n114875) );
  AOI22_X1 U86700 ( .A1(n120178), .A2(n118261), .B1(n120172), .B2(n119124), 
        .ZN(n114880) );
  AOI22_X1 U86701 ( .A1(n120154), .A2(n118748), .B1(n120148), .B2(n119060), 
        .ZN(n114882) );
  AOI22_X1 U86702 ( .A1(n120226), .A2(n118543), .B1(n120216), .B2(OUT1[57]), 
        .ZN(n114847) );
  AOI22_X1 U86703 ( .A1(n120178), .A2(n118262), .B1(n120172), .B2(n119125), 
        .ZN(n114852) );
  AOI22_X1 U86704 ( .A1(n120154), .A2(n118749), .B1(n120148), .B2(n119061), 
        .ZN(n114854) );
  AOI22_X1 U86705 ( .A1(n120226), .A2(n118544), .B1(n120216), .B2(OUT1[58]), 
        .ZN(n114819) );
  AOI22_X1 U86706 ( .A1(n120178), .A2(n118263), .B1(n120172), .B2(n119126), 
        .ZN(n114824) );
  AOI22_X1 U86707 ( .A1(n120154), .A2(n118750), .B1(n120148), .B2(n119062), 
        .ZN(n114826) );
  AOI22_X1 U86708 ( .A1(n120226), .A2(n118545), .B1(n120216), .B2(OUT1[59]), 
        .ZN(n114791) );
  AOI22_X1 U86709 ( .A1(n120178), .A2(n118264), .B1(n120172), .B2(n119127), 
        .ZN(n114796) );
  AOI22_X1 U86710 ( .A1(n120154), .A2(n118751), .B1(n120148), .B2(n119063), 
        .ZN(n114798) );
  AOI22_X1 U86711 ( .A1(n120222), .A2(n118810), .B1(n120216), .B2(OUT1[0]), 
        .ZN(n116443) );
  AOI22_X1 U86712 ( .A1(n120174), .A2(n118205), .B1(n120168), .B2(n119128), 
        .ZN(n116455) );
  AOI22_X1 U86713 ( .A1(n120150), .A2(n118752), .B1(n120144), .B2(n119064), 
        .ZN(n116460) );
  AOI22_X1 U86714 ( .A1(n120222), .A2(n118811), .B1(n120221), .B2(OUT1[1]), 
        .ZN(n116415) );
  AOI22_X1 U86715 ( .A1(n120174), .A2(n118206), .B1(n120168), .B2(n119129), 
        .ZN(n116420) );
  AOI22_X1 U86716 ( .A1(n120150), .A2(n118753), .B1(n120144), .B2(n119065), 
        .ZN(n116422) );
  AOI22_X1 U86717 ( .A1(n120222), .A2(n118812), .B1(n120221), .B2(OUT1[2]), 
        .ZN(n116387) );
  AOI22_X1 U86718 ( .A1(n120174), .A2(n118207), .B1(n120168), .B2(n119130), 
        .ZN(n116392) );
  AOI22_X1 U86719 ( .A1(n120150), .A2(n118754), .B1(n120144), .B2(n119066), 
        .ZN(n116394) );
  AOI22_X1 U86720 ( .A1(n120222), .A2(n118813), .B1(n120221), .B2(OUT1[3]), 
        .ZN(n116359) );
  AOI22_X1 U86721 ( .A1(n120174), .A2(n118208), .B1(n120168), .B2(n119131), 
        .ZN(n116364) );
  AOI22_X1 U86722 ( .A1(n120150), .A2(n118755), .B1(n120144), .B2(n119067), 
        .ZN(n116366) );
  AOI22_X1 U86723 ( .A1(n119976), .A2(n118971), .B1(n119970), .B2(n111003), 
        .ZN(n117794) );
  AOI22_X1 U86724 ( .A1(n120024), .A2(n118911), .B1(n120022), .B2(OUT2[7]), 
        .ZN(n117789) );
  AOI22_X1 U86725 ( .A1(n119952), .A2(n118332), .B1(n119946), .B2(n118212), 
        .ZN(n117796) );
  AOI22_X1 U86726 ( .A1(n119976), .A2(n118972), .B1(n119970), .B2(n111004), 
        .ZN(n117772) );
  AOI22_X1 U86727 ( .A1(n120024), .A2(n118912), .B1(n120022), .B2(OUT2[8]), 
        .ZN(n117767) );
  AOI22_X1 U86728 ( .A1(n119952), .A2(n118333), .B1(n119946), .B2(n118213), 
        .ZN(n117774) );
  AOI22_X1 U86729 ( .A1(n119976), .A2(n118973), .B1(n119970), .B2(n111005), 
        .ZN(n117750) );
  AOI22_X1 U86730 ( .A1(n120024), .A2(n118913), .B1(n120022), .B2(OUT2[9]), 
        .ZN(n117745) );
  AOI22_X1 U86731 ( .A1(n119952), .A2(n118334), .B1(n119946), .B2(n118214), 
        .ZN(n117752) );
  AOI22_X1 U86732 ( .A1(n119976), .A2(n118974), .B1(n119970), .B2(n111006), 
        .ZN(n117728) );
  AOI22_X1 U86733 ( .A1(n120024), .A2(n118914), .B1(n120022), .B2(OUT2[10]), 
        .ZN(n117723) );
  AOI22_X1 U86734 ( .A1(n119952), .A2(n118335), .B1(n119946), .B2(n118215), 
        .ZN(n117730) );
  AOI22_X1 U86735 ( .A1(n119976), .A2(n118975), .B1(n119970), .B2(n110996), 
        .ZN(n117956) );
  AOI22_X1 U86736 ( .A1(n120024), .A2(n118915), .B1(n120018), .B2(OUT2[0]), 
        .ZN(n117943) );
  AOI22_X1 U86737 ( .A1(n119952), .A2(n118325), .B1(n119946), .B2(n118205), 
        .ZN(n117960) );
  AOI22_X1 U86738 ( .A1(n119976), .A2(n118976), .B1(n119970), .B2(n110997), 
        .ZN(n117926) );
  AOI22_X1 U86739 ( .A1(n120024), .A2(n118916), .B1(n120023), .B2(OUT2[1]), 
        .ZN(n117921) );
  AOI22_X1 U86740 ( .A1(n119952), .A2(n118326), .B1(n119946), .B2(n118206), 
        .ZN(n117928) );
  AOI22_X1 U86741 ( .A1(n119976), .A2(n118977), .B1(n119970), .B2(n110998), 
        .ZN(n117904) );
  AOI22_X1 U86742 ( .A1(n120024), .A2(n118917), .B1(n120023), .B2(OUT2[2]), 
        .ZN(n117899) );
  AOI22_X1 U86743 ( .A1(n119952), .A2(n118327), .B1(n119946), .B2(n118207), 
        .ZN(n117906) );
  AOI22_X1 U86744 ( .A1(n119976), .A2(n118978), .B1(n119970), .B2(n110999), 
        .ZN(n117882) );
  AOI22_X1 U86745 ( .A1(n120024), .A2(n118918), .B1(n120023), .B2(OUT2[3]), 
        .ZN(n117877) );
  AOI22_X1 U86746 ( .A1(n119952), .A2(n118328), .B1(n119946), .B2(n118208), 
        .ZN(n117884) );
  AOI22_X1 U86747 ( .A1(n119976), .A2(n118979), .B1(n119970), .B2(n111000), 
        .ZN(n117860) );
  AOI22_X1 U86748 ( .A1(n120024), .A2(n118919), .B1(n120022), .B2(OUT2[4]), 
        .ZN(n117855) );
  AOI22_X1 U86749 ( .A1(n119952), .A2(n118329), .B1(n119946), .B2(n118209), 
        .ZN(n117862) );
  AOI22_X1 U86750 ( .A1(n119976), .A2(n118980), .B1(n119970), .B2(n111001), 
        .ZN(n117838) );
  AOI22_X1 U86751 ( .A1(n120024), .A2(n118920), .B1(n120022), .B2(OUT2[5]), 
        .ZN(n117833) );
  AOI22_X1 U86752 ( .A1(n119952), .A2(n118330), .B1(n119946), .B2(n118210), 
        .ZN(n117840) );
  AOI22_X1 U86753 ( .A1(n119976), .A2(n118981), .B1(n119970), .B2(n111002), 
        .ZN(n117816) );
  AOI22_X1 U86754 ( .A1(n120024), .A2(n118921), .B1(n120022), .B2(OUT2[6]), 
        .ZN(n117811) );
  AOI22_X1 U86755 ( .A1(n119952), .A2(n118331), .B1(n119946), .B2(n118211), 
        .ZN(n117818) );
  AOI22_X1 U86756 ( .A1(n120222), .A2(n118814), .B1(n120220), .B2(OUT1[4]), 
        .ZN(n116331) );
  AOI22_X1 U86757 ( .A1(n120174), .A2(n118209), .B1(n120168), .B2(n119132), 
        .ZN(n116336) );
  AOI22_X1 U86758 ( .A1(n120150), .A2(n118756), .B1(n120144), .B2(n119068), 
        .ZN(n116338) );
  AOI22_X1 U86759 ( .A1(n120222), .A2(n118815), .B1(n120220), .B2(OUT1[5]), 
        .ZN(n116303) );
  AOI22_X1 U86760 ( .A1(n120174), .A2(n118210), .B1(n120168), .B2(n119133), 
        .ZN(n116308) );
  AOI22_X1 U86761 ( .A1(n120150), .A2(n118757), .B1(n120144), .B2(n119069), 
        .ZN(n116310) );
  AOI22_X1 U86762 ( .A1(n120222), .A2(n118816), .B1(n120220), .B2(OUT1[6]), 
        .ZN(n116275) );
  AOI22_X1 U86763 ( .A1(n120174), .A2(n118211), .B1(n120168), .B2(n119134), 
        .ZN(n116280) );
  AOI22_X1 U86764 ( .A1(n120150), .A2(n118758), .B1(n120144), .B2(n119070), 
        .ZN(n116282) );
  AOI22_X1 U86765 ( .A1(n120222), .A2(n118806), .B1(n120220), .B2(OUT1[7]), 
        .ZN(n116247) );
  AOI22_X1 U86766 ( .A1(n120174), .A2(n118212), .B1(n120168), .B2(n119135), 
        .ZN(n116252) );
  AOI22_X1 U86767 ( .A1(n120150), .A2(n118759), .B1(n120144), .B2(n119071), 
        .ZN(n116254) );
  AOI22_X1 U86768 ( .A1(n120222), .A2(n118807), .B1(n120220), .B2(OUT1[8]), 
        .ZN(n116219) );
  AOI22_X1 U86769 ( .A1(n120174), .A2(n118213), .B1(n120168), .B2(n119136), 
        .ZN(n116224) );
  AOI22_X1 U86770 ( .A1(n120150), .A2(n118760), .B1(n120144), .B2(n119072), 
        .ZN(n116226) );
  AOI22_X1 U86771 ( .A1(n120222), .A2(n118808), .B1(n120220), .B2(OUT1[9]), 
        .ZN(n116191) );
  AOI22_X1 U86772 ( .A1(n120174), .A2(n118214), .B1(n120168), .B2(n119137), 
        .ZN(n116196) );
  AOI22_X1 U86773 ( .A1(n120150), .A2(n118761), .B1(n120144), .B2(n119073), 
        .ZN(n116198) );
  AOI22_X1 U86774 ( .A1(n120222), .A2(n118809), .B1(n120220), .B2(OUT1[10]), 
        .ZN(n116163) );
  AOI22_X1 U86775 ( .A1(n120174), .A2(n118215), .B1(n120168), .B2(n119138), 
        .ZN(n116168) );
  AOI22_X1 U86776 ( .A1(n120150), .A2(n118762), .B1(n120144), .B2(n119074), 
        .ZN(n116170) );
  AOI22_X1 U86777 ( .A1(n120222), .A2(n118798), .B1(n120220), .B2(OUT1[11]), 
        .ZN(n116135) );
  AOI22_X1 U86778 ( .A1(n120174), .A2(n118216), .B1(n120168), .B2(n119139), 
        .ZN(n116140) );
  AOI22_X1 U86779 ( .A1(n120150), .A2(n118763), .B1(n120144), .B2(n119075), 
        .ZN(n116142) );
  AOI22_X1 U86780 ( .A1(n120223), .A2(n118799), .B1(n120220), .B2(OUT1[12]), 
        .ZN(n116107) );
  AOI22_X1 U86781 ( .A1(n120175), .A2(n118217), .B1(n120169), .B2(n119140), 
        .ZN(n116112) );
  AOI22_X1 U86782 ( .A1(n120151), .A2(n118764), .B1(n120145), .B2(n119076), 
        .ZN(n116114) );
  AOI22_X1 U86783 ( .A1(n120223), .A2(n118800), .B1(n120220), .B2(OUT1[13]), 
        .ZN(n116079) );
  AOI22_X1 U86784 ( .A1(n120175), .A2(n118218), .B1(n120169), .B2(n119141), 
        .ZN(n116084) );
  AOI22_X1 U86785 ( .A1(n120151), .A2(n118765), .B1(n120145), .B2(n119077), 
        .ZN(n116086) );
  AOI22_X1 U86786 ( .A1(n120223), .A2(n118801), .B1(n120220), .B2(OUT1[14]), 
        .ZN(n116051) );
  AOI22_X1 U86787 ( .A1(n120175), .A2(n118219), .B1(n120169), .B2(n119142), 
        .ZN(n116056) );
  AOI22_X1 U86788 ( .A1(n120151), .A2(n118766), .B1(n120145), .B2(n119078), 
        .ZN(n116058) );
  AOI22_X1 U86789 ( .A1(n120223), .A2(n118802), .B1(n120220), .B2(OUT1[15]), 
        .ZN(n116023) );
  AOI22_X1 U86790 ( .A1(n120175), .A2(n118220), .B1(n120169), .B2(n119143), 
        .ZN(n116028) );
  AOI22_X1 U86791 ( .A1(n120151), .A2(n118767), .B1(n120145), .B2(n119079), 
        .ZN(n116030) );
  AOI22_X1 U86792 ( .A1(n120223), .A2(n118803), .B1(n120220), .B2(OUT1[16]), 
        .ZN(n115995) );
  AOI22_X1 U86793 ( .A1(n120175), .A2(n118221), .B1(n120169), .B2(n119144), 
        .ZN(n116000) );
  AOI22_X1 U86794 ( .A1(n120151), .A2(n118768), .B1(n120145), .B2(n119080), 
        .ZN(n116002) );
  AOI22_X1 U86795 ( .A1(n120223), .A2(n118804), .B1(n120219), .B2(OUT1[17]), 
        .ZN(n115967) );
  AOI22_X1 U86796 ( .A1(n120175), .A2(n118222), .B1(n120169), .B2(n119145), 
        .ZN(n115972) );
  AOI22_X1 U86797 ( .A1(n120151), .A2(n118769), .B1(n120145), .B2(n119081), 
        .ZN(n115974) );
  AOI22_X1 U86798 ( .A1(n120223), .A2(n118805), .B1(n120219), .B2(OUT1[18]), 
        .ZN(n115939) );
  AOI22_X1 U86799 ( .A1(n120175), .A2(n118223), .B1(n120169), .B2(n119146), 
        .ZN(n115944) );
  AOI22_X1 U86800 ( .A1(n120151), .A2(n118770), .B1(n120145), .B2(n119082), 
        .ZN(n115946) );
  AOI22_X1 U86801 ( .A1(n120223), .A2(n118505), .B1(n120219), .B2(OUT1[19]), 
        .ZN(n115911) );
  AOI22_X1 U86802 ( .A1(n120175), .A2(n118224), .B1(n120169), .B2(n119147), 
        .ZN(n115916) );
  AOI22_X1 U86803 ( .A1(n120151), .A2(n118771), .B1(n120145), .B2(n119083), 
        .ZN(n115918) );
  AOI22_X1 U86804 ( .A1(n120223), .A2(n118506), .B1(n120219), .B2(OUT1[20]), 
        .ZN(n115883) );
  AOI22_X1 U86805 ( .A1(n120175), .A2(n118225), .B1(n120169), .B2(n119148), 
        .ZN(n115888) );
  AOI22_X1 U86806 ( .A1(n120151), .A2(n118772), .B1(n120145), .B2(n119084), 
        .ZN(n115890) );
  AOI22_X1 U86807 ( .A1(n120223), .A2(n118507), .B1(n120219), .B2(OUT1[21]), 
        .ZN(n115855) );
  AOI22_X1 U86808 ( .A1(n120175), .A2(n118226), .B1(n120169), .B2(n119149), 
        .ZN(n115860) );
  AOI22_X1 U86809 ( .A1(n120151), .A2(n118773), .B1(n120145), .B2(n119085), 
        .ZN(n115862) );
  AOI22_X1 U86810 ( .A1(n120223), .A2(n118508), .B1(n120219), .B2(OUT1[22]), 
        .ZN(n115827) );
  AOI22_X1 U86811 ( .A1(n120175), .A2(n118227), .B1(n120169), .B2(n119150), 
        .ZN(n115832) );
  AOI22_X1 U86812 ( .A1(n120151), .A2(n118774), .B1(n120145), .B2(n119086), 
        .ZN(n115834) );
  AOI22_X1 U86813 ( .A1(n120223), .A2(n118509), .B1(n120219), .B2(OUT1[23]), 
        .ZN(n115799) );
  AOI22_X1 U86814 ( .A1(n120175), .A2(n118228), .B1(n120169), .B2(n119151), 
        .ZN(n115804) );
  AOI22_X1 U86815 ( .A1(n120151), .A2(n118775), .B1(n120145), .B2(n119087), 
        .ZN(n115806) );
  AOI22_X1 U86816 ( .A1(n120224), .A2(n118510), .B1(n120219), .B2(OUT1[24]), 
        .ZN(n115771) );
  AOI22_X1 U86817 ( .A1(n120176), .A2(n118229), .B1(n120170), .B2(n119152), 
        .ZN(n115776) );
  AOI22_X1 U86818 ( .A1(n120152), .A2(n118776), .B1(n120146), .B2(n119088), 
        .ZN(n115778) );
  AOI22_X1 U86819 ( .A1(n120224), .A2(n118511), .B1(n120219), .B2(OUT1[25]), 
        .ZN(n115743) );
  AOI22_X1 U86820 ( .A1(n120176), .A2(n118230), .B1(n120170), .B2(n119153), 
        .ZN(n115748) );
  AOI22_X1 U86821 ( .A1(n120152), .A2(n118777), .B1(n120146), .B2(n119089), 
        .ZN(n115750) );
  AOI22_X1 U86822 ( .A1(n120224), .A2(n118512), .B1(n120219), .B2(OUT1[26]), 
        .ZN(n115715) );
  AOI22_X1 U86823 ( .A1(n120176), .A2(n118231), .B1(n120170), .B2(n119154), 
        .ZN(n115720) );
  AOI22_X1 U86824 ( .A1(n120152), .A2(n118778), .B1(n120146), .B2(n119090), 
        .ZN(n115722) );
  AOI22_X1 U86825 ( .A1(n120224), .A2(n118513), .B1(n120219), .B2(OUT1[27]), 
        .ZN(n115687) );
  AOI22_X1 U86826 ( .A1(n120176), .A2(n118232), .B1(n120170), .B2(n119155), 
        .ZN(n115692) );
  AOI22_X1 U86827 ( .A1(n120152), .A2(n118779), .B1(n120146), .B2(n119091), 
        .ZN(n115694) );
  AOI22_X1 U86828 ( .A1(n120224), .A2(n118514), .B1(n120219), .B2(OUT1[28]), 
        .ZN(n115659) );
  AOI22_X1 U86829 ( .A1(n120176), .A2(n118233), .B1(n120170), .B2(n119156), 
        .ZN(n115664) );
  AOI22_X1 U86830 ( .A1(n120152), .A2(n118780), .B1(n120146), .B2(n119092), 
        .ZN(n115666) );
  AOI22_X1 U86831 ( .A1(n120224), .A2(n118515), .B1(n120219), .B2(OUT1[29]), 
        .ZN(n115631) );
  AOI22_X1 U86832 ( .A1(n120176), .A2(n118234), .B1(n120170), .B2(n119157), 
        .ZN(n115636) );
  AOI22_X1 U86833 ( .A1(n120152), .A2(n118781), .B1(n120146), .B2(n119093), 
        .ZN(n115638) );
  AOI22_X1 U86834 ( .A1(n120224), .A2(n118516), .B1(n120218), .B2(OUT1[30]), 
        .ZN(n115603) );
  AOI22_X1 U86835 ( .A1(n120176), .A2(n118235), .B1(n120170), .B2(n119158), 
        .ZN(n115608) );
  AOI22_X1 U86836 ( .A1(n120152), .A2(n118782), .B1(n120146), .B2(n119094), 
        .ZN(n115610) );
  AOI22_X1 U86837 ( .A1(n120224), .A2(n118517), .B1(n120218), .B2(OUT1[31]), 
        .ZN(n115575) );
  AOI22_X1 U86838 ( .A1(n120176), .A2(n118236), .B1(n120170), .B2(n119159), 
        .ZN(n115580) );
  AOI22_X1 U86839 ( .A1(n120152), .A2(n118783), .B1(n120146), .B2(n119095), 
        .ZN(n115582) );
  AOI22_X1 U86840 ( .A1(n120224), .A2(n118518), .B1(n120218), .B2(OUT1[32]), 
        .ZN(n115547) );
  AOI22_X1 U86841 ( .A1(n120176), .A2(n118237), .B1(n120170), .B2(n119160), 
        .ZN(n115552) );
  AOI22_X1 U86842 ( .A1(n120152), .A2(n118784), .B1(n120146), .B2(n119096), 
        .ZN(n115554) );
  AOI22_X1 U86843 ( .A1(n120224), .A2(n118519), .B1(n120218), .B2(OUT1[33]), 
        .ZN(n115519) );
  AOI22_X1 U86844 ( .A1(n120176), .A2(n118238), .B1(n120170), .B2(n119161), 
        .ZN(n115524) );
  AOI22_X1 U86845 ( .A1(n120152), .A2(n118785), .B1(n120146), .B2(n119097), 
        .ZN(n115526) );
  AOI22_X1 U86846 ( .A1(n120224), .A2(n118520), .B1(n120218), .B2(OUT1[34]), 
        .ZN(n115491) );
  AOI22_X1 U86847 ( .A1(n120176), .A2(n118239), .B1(n120170), .B2(n119162), 
        .ZN(n115496) );
  AOI22_X1 U86848 ( .A1(n120152), .A2(n118786), .B1(n120146), .B2(n119098), 
        .ZN(n115498) );
  AOI22_X1 U86849 ( .A1(n120224), .A2(n118521), .B1(n120218), .B2(OUT1[35]), 
        .ZN(n115463) );
  AOI22_X1 U86850 ( .A1(n120176), .A2(n118240), .B1(n120170), .B2(n119163), 
        .ZN(n115468) );
  AOI22_X1 U86851 ( .A1(n120152), .A2(n118787), .B1(n120146), .B2(n119099), 
        .ZN(n115470) );
  AOI22_X1 U86852 ( .A1(n120225), .A2(n118522), .B1(n120218), .B2(OUT1[36]), 
        .ZN(n115435) );
  AOI22_X1 U86853 ( .A1(n120177), .A2(n118241), .B1(n120171), .B2(n119164), 
        .ZN(n115440) );
  AOI22_X1 U86854 ( .A1(n120153), .A2(n118788), .B1(n120147), .B2(n119100), 
        .ZN(n115442) );
  AOI22_X1 U86855 ( .A1(n120225), .A2(n118523), .B1(n120218), .B2(OUT1[37]), 
        .ZN(n115407) );
  AOI22_X1 U86856 ( .A1(n120177), .A2(n118242), .B1(n120171), .B2(n119165), 
        .ZN(n115412) );
  AOI22_X1 U86857 ( .A1(n120153), .A2(n118789), .B1(n120147), .B2(n119101), 
        .ZN(n115414) );
  AOI22_X1 U86858 ( .A1(n120225), .A2(n118524), .B1(n120218), .B2(OUT1[38]), 
        .ZN(n115379) );
  AOI22_X1 U86859 ( .A1(n120177), .A2(n118243), .B1(n120171), .B2(n119166), 
        .ZN(n115384) );
  AOI22_X1 U86860 ( .A1(n120153), .A2(n118790), .B1(n120147), .B2(n119102), 
        .ZN(n115386) );
  AOI22_X1 U86861 ( .A1(n120225), .A2(n118525), .B1(n120218), .B2(OUT1[39]), 
        .ZN(n115351) );
  AOI22_X1 U86862 ( .A1(n120177), .A2(n118244), .B1(n120171), .B2(n119167), 
        .ZN(n115356) );
  AOI22_X1 U86863 ( .A1(n120153), .A2(n118791), .B1(n120147), .B2(n119103), 
        .ZN(n115358) );
  AOI22_X1 U86864 ( .A1(n120225), .A2(n118526), .B1(n120218), .B2(OUT1[40]), 
        .ZN(n115323) );
  AOI22_X1 U86865 ( .A1(n120177), .A2(n118245), .B1(n120171), .B2(n119168), 
        .ZN(n115328) );
  AOI22_X1 U86866 ( .A1(n120153), .A2(n118792), .B1(n120147), .B2(n119104), 
        .ZN(n115330) );
  AOI22_X1 U86867 ( .A1(n120225), .A2(n118527), .B1(n120218), .B2(OUT1[41]), 
        .ZN(n115295) );
  AOI22_X1 U86868 ( .A1(n120177), .A2(n118246), .B1(n120171), .B2(n119169), 
        .ZN(n115300) );
  AOI22_X1 U86869 ( .A1(n120153), .A2(n118793), .B1(n120147), .B2(n119105), 
        .ZN(n115302) );
  AOI22_X1 U86870 ( .A1(n120225), .A2(n118528), .B1(n120217), .B2(OUT1[42]), 
        .ZN(n115267) );
  AOI22_X1 U86871 ( .A1(n120177), .A2(n118247), .B1(n120171), .B2(n119170), 
        .ZN(n115272) );
  AOI22_X1 U86872 ( .A1(n120153), .A2(n118794), .B1(n120147), .B2(n119106), 
        .ZN(n115274) );
  AOI22_X1 U86873 ( .A1(n120225), .A2(n118529), .B1(n120217), .B2(OUT1[43]), 
        .ZN(n115239) );
  AOI22_X1 U86874 ( .A1(n120177), .A2(n118248), .B1(n120171), .B2(n119171), 
        .ZN(n115244) );
  AOI22_X1 U86875 ( .A1(n120153), .A2(n118795), .B1(n120147), .B2(n119107), 
        .ZN(n115246) );
  AOI22_X1 U86876 ( .A1(n120225), .A2(n118530), .B1(n120217), .B2(OUT1[44]), 
        .ZN(n115211) );
  AOI22_X1 U86877 ( .A1(n120177), .A2(n118249), .B1(n120171), .B2(n119172), 
        .ZN(n115216) );
  AOI22_X1 U86878 ( .A1(n120153), .A2(n118796), .B1(n120147), .B2(n119108), 
        .ZN(n115218) );
  AOI22_X1 U86879 ( .A1(n120225), .A2(n118531), .B1(n120217), .B2(OUT1[45]), 
        .ZN(n115183) );
  AOI22_X1 U86880 ( .A1(n120177), .A2(n118250), .B1(n120171), .B2(n119173), 
        .ZN(n115188) );
  AOI22_X1 U86881 ( .A1(n120153), .A2(n118797), .B1(n120147), .B2(n119109), 
        .ZN(n115190) );
  OAI221_X1 U86882 ( .B1(n99967), .B2(n120012), .C1(n114431), .C2(n120006), 
        .A(n117703), .ZN(n117699) );
  AOI22_X1 U86883 ( .A1(n120000), .A2(n118670), .B1(n119994), .B2(n119302), 
        .ZN(n117703) );
  OAI221_X1 U86884 ( .B1(n99966), .B2(n120013), .C1(n114430), .C2(n120007), 
        .A(n117681), .ZN(n117677) );
  AOI22_X1 U86885 ( .A1(n120001), .A2(n118671), .B1(n119995), .B2(n119303), 
        .ZN(n117681) );
  OAI221_X1 U86886 ( .B1(n99965), .B2(n120013), .C1(n114429), .C2(n120007), 
        .A(n117659), .ZN(n117655) );
  AOI22_X1 U86887 ( .A1(n120001), .A2(n118672), .B1(n119995), .B2(n119304), 
        .ZN(n117659) );
  OAI221_X1 U86888 ( .B1(n99964), .B2(n120013), .C1(n114428), .C2(n120007), 
        .A(n117637), .ZN(n117633) );
  AOI22_X1 U86889 ( .A1(n120001), .A2(n118673), .B1(n119995), .B2(n119305), 
        .ZN(n117637) );
  OAI221_X1 U86890 ( .B1(n99963), .B2(n120013), .C1(n114427), .C2(n120007), 
        .A(n117615), .ZN(n117611) );
  AOI22_X1 U86891 ( .A1(n120001), .A2(n118674), .B1(n119995), .B2(n119306), 
        .ZN(n117615) );
  OAI221_X1 U86892 ( .B1(n99962), .B2(n120013), .C1(n114426), .C2(n120007), 
        .A(n117593), .ZN(n117589) );
  AOI22_X1 U86893 ( .A1(n120001), .A2(n118675), .B1(n119995), .B2(n119307), 
        .ZN(n117593) );
  OAI221_X1 U86894 ( .B1(n99961), .B2(n120013), .C1(n114425), .C2(n120007), 
        .A(n117571), .ZN(n117567) );
  AOI22_X1 U86895 ( .A1(n120001), .A2(n118676), .B1(n119995), .B2(n119308), 
        .ZN(n117571) );
  OAI221_X1 U86896 ( .B1(n99960), .B2(n120013), .C1(n114424), .C2(n120007), 
        .A(n117549), .ZN(n117545) );
  AOI22_X1 U86897 ( .A1(n120001), .A2(n118677), .B1(n119995), .B2(n119309), 
        .ZN(n117549) );
  OAI221_X1 U86898 ( .B1(n99959), .B2(n120013), .C1(n114423), .C2(n120007), 
        .A(n117526), .ZN(n117522) );
  AOI22_X1 U86899 ( .A1(n120001), .A2(n118678), .B1(n119995), .B2(n119310), 
        .ZN(n117526) );
  OAI221_X1 U86900 ( .B1(n99958), .B2(n120013), .C1(n114422), .C2(n120007), 
        .A(n117503), .ZN(n117499) );
  AOI22_X1 U86901 ( .A1(n120001), .A2(n118679), .B1(n119995), .B2(n119311), 
        .ZN(n117503) );
  OAI221_X1 U86902 ( .B1(n99957), .B2(n120013), .C1(n114421), .C2(n120007), 
        .A(n117480), .ZN(n117476) );
  AOI22_X1 U86903 ( .A1(n120001), .A2(n118680), .B1(n119995), .B2(n119312), 
        .ZN(n117480) );
  OAI221_X1 U86904 ( .B1(n99956), .B2(n120013), .C1(n114420), .C2(n120007), 
        .A(n117457), .ZN(n117453) );
  AOI22_X1 U86905 ( .A1(n120001), .A2(n118681), .B1(n119995), .B2(n119313), 
        .ZN(n117457) );
  OAI221_X1 U86906 ( .B1(n99955), .B2(n120013), .C1(n114419), .C2(n120007), 
        .A(n117434), .ZN(n117430) );
  AOI22_X1 U86907 ( .A1(n120001), .A2(n118682), .B1(n119995), .B2(n119314), 
        .ZN(n117434) );
  OAI221_X1 U86908 ( .B1(n99954), .B2(n120014), .C1(n114418), .C2(n120008), 
        .A(n117411), .ZN(n117407) );
  AOI22_X1 U86909 ( .A1(n120002), .A2(n118683), .B1(n119996), .B2(n119315), 
        .ZN(n117411) );
  OAI221_X1 U86910 ( .B1(n99953), .B2(n120014), .C1(n114417), .C2(n120008), 
        .A(n117388), .ZN(n117384) );
  AOI22_X1 U86911 ( .A1(n120002), .A2(n118684), .B1(n119996), .B2(n119316), 
        .ZN(n117388) );
  OAI221_X1 U86912 ( .B1(n99952), .B2(n120014), .C1(n114416), .C2(n120008), 
        .A(n117365), .ZN(n117361) );
  AOI22_X1 U86913 ( .A1(n120002), .A2(n118685), .B1(n119996), .B2(n119317), 
        .ZN(n117365) );
  OAI221_X1 U86914 ( .B1(n99951), .B2(n120014), .C1(n114415), .C2(n120008), 
        .A(n117342), .ZN(n117338) );
  AOI22_X1 U86915 ( .A1(n120002), .A2(n118686), .B1(n119996), .B2(n119318), 
        .ZN(n117342) );
  OAI221_X1 U86916 ( .B1(n99950), .B2(n120014), .C1(n114414), .C2(n120008), 
        .A(n117319), .ZN(n117315) );
  AOI22_X1 U86917 ( .A1(n120002), .A2(n118687), .B1(n119996), .B2(n119319), 
        .ZN(n117319) );
  OAI221_X1 U86918 ( .B1(n99949), .B2(n120014), .C1(n114413), .C2(n120008), 
        .A(n117296), .ZN(n117292) );
  AOI22_X1 U86919 ( .A1(n120002), .A2(n118688), .B1(n119996), .B2(n119320), 
        .ZN(n117296) );
  OAI221_X1 U86920 ( .B1(n99948), .B2(n120014), .C1(n114412), .C2(n120008), 
        .A(n117273), .ZN(n117269) );
  AOI22_X1 U86921 ( .A1(n120002), .A2(n118689), .B1(n119996), .B2(n119321), 
        .ZN(n117273) );
  OAI221_X1 U86922 ( .B1(n99947), .B2(n120014), .C1(n114411), .C2(n120008), 
        .A(n117250), .ZN(n117246) );
  AOI22_X1 U86923 ( .A1(n120002), .A2(n118690), .B1(n119996), .B2(n119322), 
        .ZN(n117250) );
  OAI221_X1 U86924 ( .B1(n99946), .B2(n120014), .C1(n114410), .C2(n120008), 
        .A(n117227), .ZN(n117223) );
  AOI22_X1 U86925 ( .A1(n120002), .A2(n118691), .B1(n119996), .B2(n119323), 
        .ZN(n117227) );
  OAI221_X1 U86926 ( .B1(n99945), .B2(n120014), .C1(n114409), .C2(n120008), 
        .A(n117204), .ZN(n117200) );
  AOI22_X1 U86927 ( .A1(n120002), .A2(n118692), .B1(n119996), .B2(n119324), 
        .ZN(n117204) );
  OAI221_X1 U86928 ( .B1(n99944), .B2(n120014), .C1(n114408), .C2(n120008), 
        .A(n117181), .ZN(n117177) );
  AOI22_X1 U86929 ( .A1(n120002), .A2(n118693), .B1(n119996), .B2(n119325), 
        .ZN(n117181) );
  OAI221_X1 U86930 ( .B1(n99943), .B2(n120014), .C1(n114407), .C2(n120008), 
        .A(n117158), .ZN(n117154) );
  AOI22_X1 U86931 ( .A1(n120002), .A2(n118694), .B1(n119996), .B2(n119326), 
        .ZN(n117158) );
  OAI221_X1 U86932 ( .B1(n99942), .B2(n120015), .C1(n114406), .C2(n120009), 
        .A(n117135), .ZN(n117131) );
  AOI22_X1 U86933 ( .A1(n120003), .A2(n118695), .B1(n119997), .B2(n119327), 
        .ZN(n117135) );
  OAI221_X1 U86934 ( .B1(n99941), .B2(n120015), .C1(n114405), .C2(n120009), 
        .A(n117112), .ZN(n117108) );
  AOI22_X1 U86935 ( .A1(n120003), .A2(n118696), .B1(n119997), .B2(n119328), 
        .ZN(n117112) );
  OAI221_X1 U86936 ( .B1(n99940), .B2(n120015), .C1(n114404), .C2(n120009), 
        .A(n117089), .ZN(n117085) );
  AOI22_X1 U86937 ( .A1(n120003), .A2(n118697), .B1(n119997), .B2(n119329), 
        .ZN(n117089) );
  OAI221_X1 U86938 ( .B1(n99939), .B2(n120015), .C1(n114403), .C2(n120009), 
        .A(n117066), .ZN(n117062) );
  AOI22_X1 U86939 ( .A1(n120003), .A2(n118698), .B1(n119997), .B2(n119330), 
        .ZN(n117066) );
  OAI221_X1 U86940 ( .B1(n99938), .B2(n120015), .C1(n114402), .C2(n120009), 
        .A(n117043), .ZN(n117039) );
  AOI22_X1 U86941 ( .A1(n120003), .A2(n118699), .B1(n119997), .B2(n119331), 
        .ZN(n117043) );
  OAI221_X1 U86942 ( .B1(n99937), .B2(n120015), .C1(n114401), .C2(n120009), 
        .A(n117020), .ZN(n117016) );
  AOI22_X1 U86943 ( .A1(n120003), .A2(n118700), .B1(n119997), .B2(n119332), 
        .ZN(n117020) );
  OAI221_X1 U86944 ( .B1(n99936), .B2(n120015), .C1(n114400), .C2(n120009), 
        .A(n116997), .ZN(n116993) );
  AOI22_X1 U86945 ( .A1(n120003), .A2(n118701), .B1(n119997), .B2(n119333), 
        .ZN(n116997) );
  OAI221_X1 U86946 ( .B1(n99935), .B2(n120015), .C1(n114399), .C2(n120009), 
        .A(n116974), .ZN(n116970) );
  AOI22_X1 U86947 ( .A1(n120003), .A2(n118702), .B1(n119997), .B2(n119334), 
        .ZN(n116974) );
  OAI221_X1 U86948 ( .B1(n99934), .B2(n120015), .C1(n114398), .C2(n120009), 
        .A(n116951), .ZN(n116947) );
  AOI22_X1 U86949 ( .A1(n120003), .A2(n118703), .B1(n119997), .B2(n119335), 
        .ZN(n116951) );
  OAI221_X1 U86950 ( .B1(n99933), .B2(n120015), .C1(n114397), .C2(n120009), 
        .A(n116928), .ZN(n116924) );
  AOI22_X1 U86951 ( .A1(n120003), .A2(n118704), .B1(n119997), .B2(n119336), 
        .ZN(n116928) );
  OAI221_X1 U86952 ( .B1(n99932), .B2(n120015), .C1(n114396), .C2(n120009), 
        .A(n116905), .ZN(n116901) );
  AOI22_X1 U86953 ( .A1(n120003), .A2(n118705), .B1(n119997), .B2(n119337), 
        .ZN(n116905) );
  OAI221_X1 U86954 ( .B1(n99931), .B2(n120015), .C1(n114395), .C2(n120009), 
        .A(n116882), .ZN(n116878) );
  AOI22_X1 U86955 ( .A1(n120003), .A2(n118706), .B1(n119997), .B2(n119338), 
        .ZN(n116882) );
  OAI221_X1 U86956 ( .B1(n99930), .B2(n120016), .C1(n114394), .C2(n120010), 
        .A(n116859), .ZN(n116855) );
  AOI22_X1 U86957 ( .A1(n120004), .A2(n118707), .B1(n119998), .B2(n119339), 
        .ZN(n116859) );
  OAI221_X1 U86958 ( .B1(n99929), .B2(n120016), .C1(n114393), .C2(n120010), 
        .A(n116836), .ZN(n116832) );
  AOI22_X1 U86959 ( .A1(n120004), .A2(n118708), .B1(n119998), .B2(n119340), 
        .ZN(n116836) );
  OAI221_X1 U86960 ( .B1(n99928), .B2(n120016), .C1(n114392), .C2(n120010), 
        .A(n116813), .ZN(n116809) );
  AOI22_X1 U86961 ( .A1(n120004), .A2(n118709), .B1(n119998), .B2(n119341), 
        .ZN(n116813) );
  OAI221_X1 U86962 ( .B1(n99927), .B2(n120016), .C1(n114391), .C2(n120010), 
        .A(n116790), .ZN(n116786) );
  AOI22_X1 U86963 ( .A1(n120004), .A2(n118710), .B1(n119998), .B2(n119342), 
        .ZN(n116790) );
  OAI221_X1 U86964 ( .B1(n99926), .B2(n120016), .C1(n114390), .C2(n120010), 
        .A(n116767), .ZN(n116763) );
  AOI22_X1 U86965 ( .A1(n120004), .A2(n118711), .B1(n119998), .B2(n119343), 
        .ZN(n116767) );
  OAI221_X1 U86966 ( .B1(n99925), .B2(n120016), .C1(n114389), .C2(n120010), 
        .A(n116744), .ZN(n116740) );
  AOI22_X1 U86967 ( .A1(n120004), .A2(n118712), .B1(n119998), .B2(n119344), 
        .ZN(n116744) );
  OAI221_X1 U86968 ( .B1(n99924), .B2(n120016), .C1(n114388), .C2(n120010), 
        .A(n116721), .ZN(n116717) );
  AOI22_X1 U86969 ( .A1(n120004), .A2(n118713), .B1(n119998), .B2(n119345), 
        .ZN(n116721) );
  OAI221_X1 U86970 ( .B1(n99923), .B2(n120016), .C1(n114387), .C2(n120010), 
        .A(n116698), .ZN(n116694) );
  AOI22_X1 U86971 ( .A1(n120004), .A2(n118714), .B1(n119998), .B2(n119346), 
        .ZN(n116698) );
  OAI221_X1 U86972 ( .B1(n99922), .B2(n120016), .C1(n114386), .C2(n120010), 
        .A(n116675), .ZN(n116671) );
  AOI22_X1 U86973 ( .A1(n120004), .A2(n118715), .B1(n119998), .B2(n119347), 
        .ZN(n116675) );
  OAI221_X1 U86974 ( .B1(n99921), .B2(n120016), .C1(n114385), .C2(n120010), 
        .A(n116652), .ZN(n116648) );
  AOI22_X1 U86975 ( .A1(n120004), .A2(n118716), .B1(n119998), .B2(n119348), 
        .ZN(n116652) );
  OAI221_X1 U86976 ( .B1(n99920), .B2(n120016), .C1(n114384), .C2(n120010), 
        .A(n116629), .ZN(n116625) );
  AOI22_X1 U86977 ( .A1(n120004), .A2(n118717), .B1(n119998), .B2(n119349), 
        .ZN(n116629) );
  OAI221_X1 U86978 ( .B1(n99919), .B2(n120016), .C1(n114383), .C2(n120010), 
        .A(n116606), .ZN(n116602) );
  AOI22_X1 U86979 ( .A1(n120004), .A2(n118718), .B1(n119998), .B2(n119350), 
        .ZN(n116606) );
  OAI221_X1 U86980 ( .B1(n114150), .B2(n120215), .C1(n98652), .C2(n120209), 
        .A(n114766), .ZN(n114763) );
  AOI22_X1 U86981 ( .A1(n120203), .A2(n118719), .B1(n120197), .B2(n119298), 
        .ZN(n114766) );
  OAI221_X1 U86982 ( .B1(n114149), .B2(n120215), .C1(n98651), .C2(n120209), 
        .A(n114740), .ZN(n114737) );
  AOI22_X1 U86983 ( .A1(n120203), .A2(n118720), .B1(n120197), .B2(n119299), 
        .ZN(n114740) );
  OAI221_X1 U86984 ( .B1(n114148), .B2(n120215), .C1(n98650), .C2(n120209), 
        .A(n114714), .ZN(n114711) );
  AOI22_X1 U86985 ( .A1(n120203), .A2(n118721), .B1(n120197), .B2(n119300), 
        .ZN(n114714) );
  OAI221_X1 U86986 ( .B1(n114146), .B2(n120215), .C1(n98648), .C2(n120209), 
        .A(n114661), .ZN(n114652) );
  AOI22_X1 U86987 ( .A1(n120203), .A2(n118722), .B1(n120197), .B2(n119301), 
        .ZN(n114661) );
  OAI221_X1 U86988 ( .B1(n99918), .B2(n120017), .C1(n114382), .C2(n120011), 
        .A(n116584), .ZN(n116581) );
  AOI22_X1 U86989 ( .A1(n120005), .A2(n118723), .B1(n119999), .B2(n119351), 
        .ZN(n116584) );
  OAI221_X1 U86990 ( .B1(n99917), .B2(n120017), .C1(n114381), .C2(n120011), 
        .A(n116563), .ZN(n116560) );
  AOI22_X1 U86991 ( .A1(n120005), .A2(n118724), .B1(n119999), .B2(n119352), 
        .ZN(n116563) );
  OAI221_X1 U86992 ( .B1(n99916), .B2(n120017), .C1(n114380), .C2(n120011), 
        .A(n116542), .ZN(n116539) );
  AOI22_X1 U86993 ( .A1(n120005), .A2(n118725), .B1(n119999), .B2(n119353), 
        .ZN(n116542) );
  OAI221_X1 U86994 ( .B1(n99914), .B2(n120017), .C1(n114378), .C2(n120011), 
        .A(n116494), .ZN(n116485) );
  AOI22_X1 U86995 ( .A1(n120005), .A2(n118726), .B1(n119999), .B2(n119354), 
        .ZN(n116494) );
  OAI221_X1 U86996 ( .B1(n99971), .B2(n120012), .C1(n114435), .C2(n120006), 
        .A(n117791), .ZN(n117787) );
  AOI22_X1 U86997 ( .A1(n120000), .A2(n118727), .B1(n119994), .B2(n119355), 
        .ZN(n117791) );
  OAI221_X1 U86998 ( .B1(n99970), .B2(n120012), .C1(n114434), .C2(n120006), 
        .A(n117769), .ZN(n117765) );
  AOI22_X1 U86999 ( .A1(n120000), .A2(n118728), .B1(n119994), .B2(n119356), 
        .ZN(n117769) );
  OAI221_X1 U87000 ( .B1(n99969), .B2(n120012), .C1(n114433), .C2(n120006), 
        .A(n117747), .ZN(n117743) );
  AOI22_X1 U87001 ( .A1(n120000), .A2(n118729), .B1(n119994), .B2(n119357), 
        .ZN(n117747) );
  OAI221_X1 U87002 ( .B1(n99968), .B2(n120012), .C1(n114432), .C2(n120006), 
        .A(n117725), .ZN(n117721) );
  AOI22_X1 U87003 ( .A1(n120000), .A2(n118730), .B1(n119994), .B2(n119358), 
        .ZN(n117725) );
  OAI221_X1 U87004 ( .B1(n99978), .B2(n120012), .C1(n114442), .C2(n120006), 
        .A(n117950), .ZN(n117941) );
  AOI22_X1 U87005 ( .A1(n120000), .A2(n118731), .B1(n119994), .B2(n119359), 
        .ZN(n117950) );
  OAI221_X1 U87006 ( .B1(n99977), .B2(n120012), .C1(n114441), .C2(n120006), 
        .A(n117923), .ZN(n117919) );
  AOI22_X1 U87007 ( .A1(n120000), .A2(n118732), .B1(n119994), .B2(n119360), 
        .ZN(n117923) );
  OAI221_X1 U87008 ( .B1(n99976), .B2(n120012), .C1(n114440), .C2(n120006), 
        .A(n117901), .ZN(n117897) );
  AOI22_X1 U87009 ( .A1(n120000), .A2(n118733), .B1(n119994), .B2(n119361), 
        .ZN(n117901) );
  OAI221_X1 U87010 ( .B1(n99975), .B2(n120012), .C1(n114439), .C2(n120006), 
        .A(n117879), .ZN(n117875) );
  AOI22_X1 U87011 ( .A1(n120000), .A2(n118734), .B1(n119994), .B2(n119362), 
        .ZN(n117879) );
  OAI221_X1 U87012 ( .B1(n99974), .B2(n120012), .C1(n114438), .C2(n120006), 
        .A(n117857), .ZN(n117853) );
  AOI22_X1 U87013 ( .A1(n120000), .A2(n118735), .B1(n119994), .B2(n119363), 
        .ZN(n117857) );
  OAI221_X1 U87014 ( .B1(n99973), .B2(n120012), .C1(n114437), .C2(n120006), 
        .A(n117835), .ZN(n117831) );
  AOI22_X1 U87015 ( .A1(n120000), .A2(n118736), .B1(n119994), .B2(n119364), 
        .ZN(n117835) );
  OAI221_X1 U87016 ( .B1(n99972), .B2(n120012), .C1(n114436), .C2(n120006), 
        .A(n117813), .ZN(n117809) );
  AOI22_X1 U87017 ( .A1(n120000), .A2(n118737), .B1(n119994), .B2(n119365), 
        .ZN(n117813) );
  OAI22_X1 U87018 ( .A1(n99780), .A2(n120323), .B1(n120631), .B2(n120317), 
        .ZN(n5823) );
  OAI22_X1 U87019 ( .A1(n99779), .A2(n120323), .B1(n120634), .B2(n120317), 
        .ZN(n5824) );
  OAI22_X1 U87020 ( .A1(n99778), .A2(n120323), .B1(n120637), .B2(n120317), 
        .ZN(n5825) );
  OAI22_X1 U87021 ( .A1(n99777), .A2(n120323), .B1(n120640), .B2(n120317), 
        .ZN(n5826) );
  OAI22_X1 U87022 ( .A1(n99776), .A2(n120323), .B1(n120643), .B2(n120317), 
        .ZN(n5827) );
  OAI22_X1 U87023 ( .A1(n99775), .A2(n120323), .B1(n120646), .B2(n120317), 
        .ZN(n5828) );
  OAI22_X1 U87024 ( .A1(n99774), .A2(n120323), .B1(n120649), .B2(n120317), 
        .ZN(n5829) );
  OAI22_X1 U87025 ( .A1(n99773), .A2(n120323), .B1(n120652), .B2(n120317), 
        .ZN(n5830) );
  OAI22_X1 U87026 ( .A1(n99772), .A2(n120323), .B1(n120655), .B2(n120317), 
        .ZN(n5831) );
  OAI22_X1 U87027 ( .A1(n99771), .A2(n120323), .B1(n120658), .B2(n120317), 
        .ZN(n5832) );
  OAI22_X1 U87028 ( .A1(n99770), .A2(n120323), .B1(n120661), .B2(n120317), 
        .ZN(n5833) );
  OAI22_X1 U87029 ( .A1(n99769), .A2(n120324), .B1(n120664), .B2(n120317), 
        .ZN(n5834) );
  OAI22_X1 U87030 ( .A1(n99768), .A2(n120324), .B1(n120667), .B2(n120318), 
        .ZN(n5835) );
  OAI22_X1 U87031 ( .A1(n99767), .A2(n120324), .B1(n120670), .B2(n120318), 
        .ZN(n5836) );
  OAI22_X1 U87032 ( .A1(n99766), .A2(n120324), .B1(n120673), .B2(n120318), 
        .ZN(n5837) );
  OAI22_X1 U87033 ( .A1(n99765), .A2(n120324), .B1(n120676), .B2(n120318), 
        .ZN(n5838) );
  OAI22_X1 U87034 ( .A1(n99764), .A2(n120324), .B1(n120679), .B2(n120318), 
        .ZN(n5839) );
  OAI22_X1 U87035 ( .A1(n99763), .A2(n120324), .B1(n120682), .B2(n120318), 
        .ZN(n5840) );
  OAI22_X1 U87036 ( .A1(n99762), .A2(n120324), .B1(n120685), .B2(n120318), 
        .ZN(n5841) );
  OAI22_X1 U87037 ( .A1(n99761), .A2(n120324), .B1(n120688), .B2(n120318), 
        .ZN(n5842) );
  OAI22_X1 U87038 ( .A1(n99760), .A2(n120324), .B1(n120691), .B2(n120318), 
        .ZN(n5843) );
  OAI22_X1 U87039 ( .A1(n99759), .A2(n120324), .B1(n120694), .B2(n120318), 
        .ZN(n5844) );
  OAI22_X1 U87040 ( .A1(n99758), .A2(n120324), .B1(n120697), .B2(n120318), 
        .ZN(n5845) );
  OAI22_X1 U87041 ( .A1(n99757), .A2(n120325), .B1(n120700), .B2(n120318), 
        .ZN(n5846) );
  OAI22_X1 U87042 ( .A1(n99756), .A2(n120325), .B1(n120703), .B2(n120319), 
        .ZN(n5847) );
  OAI22_X1 U87043 ( .A1(n99755), .A2(n120325), .B1(n120706), .B2(n120319), 
        .ZN(n5848) );
  OAI22_X1 U87044 ( .A1(n99754), .A2(n120325), .B1(n120709), .B2(n120319), 
        .ZN(n5849) );
  OAI22_X1 U87045 ( .A1(n99753), .A2(n120325), .B1(n120712), .B2(n120319), 
        .ZN(n5850) );
  OAI22_X1 U87046 ( .A1(n99752), .A2(n120325), .B1(n120715), .B2(n120319), 
        .ZN(n5851) );
  OAI22_X1 U87047 ( .A1(n99751), .A2(n120325), .B1(n120718), .B2(n120319), 
        .ZN(n5852) );
  OAI22_X1 U87048 ( .A1(n99750), .A2(n120325), .B1(n120721), .B2(n120319), 
        .ZN(n5853) );
  OAI22_X1 U87049 ( .A1(n99749), .A2(n120325), .B1(n120724), .B2(n120319), 
        .ZN(n5854) );
  OAI22_X1 U87050 ( .A1(n99748), .A2(n120325), .B1(n120727), .B2(n120319), 
        .ZN(n5855) );
  OAI22_X1 U87051 ( .A1(n99747), .A2(n120325), .B1(n120730), .B2(n120319), 
        .ZN(n5856) );
  OAI22_X1 U87052 ( .A1(n99746), .A2(n120325), .B1(n120733), .B2(n120319), 
        .ZN(n5857) );
  OAI22_X1 U87053 ( .A1(n99745), .A2(n120326), .B1(n120736), .B2(n120319), 
        .ZN(n5858) );
  OAI22_X1 U87054 ( .A1(n99744), .A2(n120326), .B1(n120739), .B2(n120320), 
        .ZN(n5859) );
  OAI22_X1 U87055 ( .A1(n99743), .A2(n120326), .B1(n120742), .B2(n120320), 
        .ZN(n5860) );
  OAI22_X1 U87056 ( .A1(n99742), .A2(n120326), .B1(n120745), .B2(n120320), 
        .ZN(n5861) );
  OAI22_X1 U87057 ( .A1(n99741), .A2(n120326), .B1(n120748), .B2(n120320), 
        .ZN(n5862) );
  OAI22_X1 U87058 ( .A1(n99740), .A2(n120326), .B1(n120751), .B2(n120320), 
        .ZN(n5863) );
  OAI22_X1 U87059 ( .A1(n99739), .A2(n120326), .B1(n120754), .B2(n120320), 
        .ZN(n5864) );
  OAI22_X1 U87060 ( .A1(n99738), .A2(n120326), .B1(n120757), .B2(n120320), 
        .ZN(n5865) );
  OAI22_X1 U87061 ( .A1(n99737), .A2(n120326), .B1(n120760), .B2(n120320), 
        .ZN(n5866) );
  OAI22_X1 U87062 ( .A1(n99736), .A2(n120326), .B1(n120763), .B2(n120320), 
        .ZN(n5867) );
  OAI22_X1 U87063 ( .A1(n99735), .A2(n120326), .B1(n120766), .B2(n120320), 
        .ZN(n5868) );
  OAI22_X1 U87064 ( .A1(n99734), .A2(n120326), .B1(n120769), .B2(n120320), 
        .ZN(n5869) );
  OAI22_X1 U87065 ( .A1(n99733), .A2(n120327), .B1(n120772), .B2(n120320), 
        .ZN(n5870) );
  OAI22_X1 U87066 ( .A1(n99732), .A2(n120327), .B1(n120775), .B2(n120321), 
        .ZN(n5871) );
  OAI22_X1 U87067 ( .A1(n99731), .A2(n120327), .B1(n120778), .B2(n120321), 
        .ZN(n5872) );
  OAI22_X1 U87068 ( .A1(n99730), .A2(n120327), .B1(n120781), .B2(n120321), 
        .ZN(n5873) );
  OAI22_X1 U87069 ( .A1(n99729), .A2(n120327), .B1(n120784), .B2(n120321), 
        .ZN(n5874) );
  OAI22_X1 U87070 ( .A1(n99728), .A2(n120327), .B1(n120787), .B2(n120321), 
        .ZN(n5875) );
  OAI22_X1 U87071 ( .A1(n99727), .A2(n120327), .B1(n120790), .B2(n120321), 
        .ZN(n5876) );
  OAI22_X1 U87072 ( .A1(n99726), .A2(n120327), .B1(n120793), .B2(n120321), 
        .ZN(n5877) );
  OAI22_X1 U87073 ( .A1(n99725), .A2(n120327), .B1(n120796), .B2(n120321), 
        .ZN(n5878) );
  OAI22_X1 U87074 ( .A1(n99724), .A2(n120327), .B1(n120799), .B2(n120321), 
        .ZN(n5879) );
  OAI22_X1 U87075 ( .A1(n99723), .A2(n120327), .B1(n120802), .B2(n120321), 
        .ZN(n5880) );
  OAI22_X1 U87076 ( .A1(n99722), .A2(n120327), .B1(n120805), .B2(n120321), 
        .ZN(n5881) );
  OAI22_X1 U87077 ( .A1(n99721), .A2(n120328), .B1(n120808), .B2(n120321), 
        .ZN(n5882) );
  OAI22_X1 U87078 ( .A1(n99978), .A2(n120272), .B1(n120631), .B2(n120266), 
        .ZN(n5567) );
  OAI22_X1 U87079 ( .A1(n99977), .A2(n120272), .B1(n120634), .B2(n120266), 
        .ZN(n5568) );
  OAI22_X1 U87080 ( .A1(n99976), .A2(n120272), .B1(n120637), .B2(n120266), 
        .ZN(n5569) );
  OAI22_X1 U87081 ( .A1(n99975), .A2(n120272), .B1(n120640), .B2(n120266), 
        .ZN(n5570) );
  OAI22_X1 U87082 ( .A1(n99974), .A2(n120272), .B1(n120643), .B2(n120266), 
        .ZN(n5571) );
  OAI22_X1 U87083 ( .A1(n99973), .A2(n120272), .B1(n120646), .B2(n120266), 
        .ZN(n5572) );
  OAI22_X1 U87084 ( .A1(n99972), .A2(n120272), .B1(n120649), .B2(n120266), 
        .ZN(n5573) );
  OAI22_X1 U87085 ( .A1(n99971), .A2(n120272), .B1(n120652), .B2(n120266), 
        .ZN(n5574) );
  OAI22_X1 U87086 ( .A1(n99970), .A2(n120272), .B1(n120655), .B2(n120266), 
        .ZN(n5575) );
  OAI22_X1 U87087 ( .A1(n99969), .A2(n120272), .B1(n120658), .B2(n120266), 
        .ZN(n5576) );
  OAI22_X1 U87088 ( .A1(n99968), .A2(n120272), .B1(n120661), .B2(n120266), 
        .ZN(n5577) );
  OAI22_X1 U87089 ( .A1(n99967), .A2(n120273), .B1(n120664), .B2(n120266), 
        .ZN(n5578) );
  OAI22_X1 U87090 ( .A1(n99966), .A2(n120273), .B1(n120667), .B2(n120267), 
        .ZN(n5579) );
  OAI22_X1 U87091 ( .A1(n99965), .A2(n120273), .B1(n120670), .B2(n120267), 
        .ZN(n5580) );
  OAI22_X1 U87092 ( .A1(n99964), .A2(n120273), .B1(n120673), .B2(n120267), 
        .ZN(n5581) );
  OAI22_X1 U87093 ( .A1(n99963), .A2(n120273), .B1(n120676), .B2(n120267), 
        .ZN(n5582) );
  OAI22_X1 U87094 ( .A1(n99962), .A2(n120273), .B1(n120679), .B2(n120267), 
        .ZN(n5583) );
  OAI22_X1 U87095 ( .A1(n99961), .A2(n120273), .B1(n120682), .B2(n120267), 
        .ZN(n5584) );
  OAI22_X1 U87096 ( .A1(n99960), .A2(n120273), .B1(n120685), .B2(n120267), 
        .ZN(n5585) );
  OAI22_X1 U87097 ( .A1(n99959), .A2(n120273), .B1(n120688), .B2(n120267), 
        .ZN(n5586) );
  OAI22_X1 U87098 ( .A1(n99958), .A2(n120273), .B1(n120691), .B2(n120267), 
        .ZN(n5587) );
  OAI22_X1 U87099 ( .A1(n99957), .A2(n120273), .B1(n120694), .B2(n120267), 
        .ZN(n5588) );
  OAI22_X1 U87100 ( .A1(n99956), .A2(n120273), .B1(n120697), .B2(n120267), 
        .ZN(n5589) );
  OAI22_X1 U87101 ( .A1(n99955), .A2(n120274), .B1(n120700), .B2(n120267), 
        .ZN(n5590) );
  OAI22_X1 U87102 ( .A1(n99954), .A2(n120274), .B1(n120703), .B2(n120268), 
        .ZN(n5591) );
  OAI22_X1 U87103 ( .A1(n99953), .A2(n120274), .B1(n120706), .B2(n120268), 
        .ZN(n5592) );
  OAI22_X1 U87104 ( .A1(n99952), .A2(n120274), .B1(n120709), .B2(n120268), 
        .ZN(n5593) );
  OAI22_X1 U87105 ( .A1(n99951), .A2(n120274), .B1(n120712), .B2(n120268), 
        .ZN(n5594) );
  OAI22_X1 U87106 ( .A1(n99950), .A2(n120274), .B1(n120715), .B2(n120268), 
        .ZN(n5595) );
  OAI22_X1 U87107 ( .A1(n99949), .A2(n120274), .B1(n120718), .B2(n120268), 
        .ZN(n5596) );
  OAI22_X1 U87108 ( .A1(n99948), .A2(n120274), .B1(n120721), .B2(n120268), 
        .ZN(n5597) );
  OAI22_X1 U87109 ( .A1(n99947), .A2(n120274), .B1(n120724), .B2(n120268), 
        .ZN(n5598) );
  OAI22_X1 U87110 ( .A1(n99946), .A2(n120274), .B1(n120727), .B2(n120268), 
        .ZN(n5599) );
  OAI22_X1 U87111 ( .A1(n99945), .A2(n120274), .B1(n120730), .B2(n120268), 
        .ZN(n5600) );
  OAI22_X1 U87112 ( .A1(n99944), .A2(n120274), .B1(n120733), .B2(n120268), 
        .ZN(n5601) );
  OAI22_X1 U87113 ( .A1(n99943), .A2(n120275), .B1(n120736), .B2(n120268), 
        .ZN(n5602) );
  OAI22_X1 U87114 ( .A1(n99942), .A2(n120275), .B1(n120739), .B2(n120269), 
        .ZN(n5603) );
  OAI22_X1 U87115 ( .A1(n99941), .A2(n120275), .B1(n120742), .B2(n120269), 
        .ZN(n5604) );
  OAI22_X1 U87116 ( .A1(n99940), .A2(n120275), .B1(n120745), .B2(n120269), 
        .ZN(n5605) );
  OAI22_X1 U87117 ( .A1(n99939), .A2(n120275), .B1(n120748), .B2(n120269), 
        .ZN(n5606) );
  OAI22_X1 U87118 ( .A1(n99938), .A2(n120275), .B1(n120751), .B2(n120269), 
        .ZN(n5607) );
  OAI22_X1 U87119 ( .A1(n99937), .A2(n120275), .B1(n120754), .B2(n120269), 
        .ZN(n5608) );
  OAI22_X1 U87120 ( .A1(n99936), .A2(n120275), .B1(n120757), .B2(n120269), 
        .ZN(n5609) );
  OAI22_X1 U87121 ( .A1(n99935), .A2(n120275), .B1(n120760), .B2(n120269), 
        .ZN(n5610) );
  OAI22_X1 U87122 ( .A1(n99934), .A2(n120275), .B1(n120763), .B2(n120269), 
        .ZN(n5611) );
  OAI22_X1 U87123 ( .A1(n99933), .A2(n120275), .B1(n120766), .B2(n120269), 
        .ZN(n5612) );
  OAI22_X1 U87124 ( .A1(n99932), .A2(n120275), .B1(n120769), .B2(n120269), 
        .ZN(n5613) );
  OAI22_X1 U87125 ( .A1(n99931), .A2(n120276), .B1(n120772), .B2(n120269), 
        .ZN(n5614) );
  OAI22_X1 U87126 ( .A1(n99930), .A2(n120276), .B1(n120775), .B2(n120270), 
        .ZN(n5615) );
  OAI22_X1 U87127 ( .A1(n99929), .A2(n120276), .B1(n120778), .B2(n120270), 
        .ZN(n5616) );
  OAI22_X1 U87128 ( .A1(n99928), .A2(n120276), .B1(n120781), .B2(n120270), 
        .ZN(n5617) );
  OAI22_X1 U87129 ( .A1(n99927), .A2(n120276), .B1(n120784), .B2(n120270), 
        .ZN(n5618) );
  OAI22_X1 U87130 ( .A1(n99926), .A2(n120276), .B1(n120787), .B2(n120270), 
        .ZN(n5619) );
  OAI22_X1 U87131 ( .A1(n99925), .A2(n120276), .B1(n120790), .B2(n120270), 
        .ZN(n5620) );
  OAI22_X1 U87132 ( .A1(n99924), .A2(n120276), .B1(n120793), .B2(n120270), 
        .ZN(n5621) );
  OAI22_X1 U87133 ( .A1(n99923), .A2(n120276), .B1(n120796), .B2(n120270), 
        .ZN(n5622) );
  OAI22_X1 U87134 ( .A1(n99922), .A2(n120276), .B1(n120799), .B2(n120270), 
        .ZN(n5623) );
  OAI22_X1 U87135 ( .A1(n99921), .A2(n120276), .B1(n120802), .B2(n120270), 
        .ZN(n5624) );
  OAI22_X1 U87136 ( .A1(n99920), .A2(n120276), .B1(n120805), .B2(n120270), 
        .ZN(n5625) );
  OAI22_X1 U87137 ( .A1(n99919), .A2(n120277), .B1(n120808), .B2(n120270), 
        .ZN(n5626) );
  OAI22_X1 U87138 ( .A1(n99243), .A2(n120470), .B1(n120630), .B2(n120464), 
        .ZN(n6591) );
  OAI22_X1 U87139 ( .A1(n99242), .A2(n120470), .B1(n120633), .B2(n120464), 
        .ZN(n6592) );
  OAI22_X1 U87140 ( .A1(n99241), .A2(n120470), .B1(n120636), .B2(n120464), 
        .ZN(n6593) );
  OAI22_X1 U87141 ( .A1(n99240), .A2(n120470), .B1(n120639), .B2(n120464), 
        .ZN(n6594) );
  OAI22_X1 U87142 ( .A1(n99239), .A2(n120470), .B1(n120642), .B2(n120464), 
        .ZN(n6595) );
  OAI22_X1 U87143 ( .A1(n99238), .A2(n120470), .B1(n120645), .B2(n120464), 
        .ZN(n6596) );
  OAI22_X1 U87144 ( .A1(n99237), .A2(n120470), .B1(n120648), .B2(n120464), 
        .ZN(n6597) );
  OAI22_X1 U87145 ( .A1(n99236), .A2(n120470), .B1(n120651), .B2(n120464), 
        .ZN(n6598) );
  OAI22_X1 U87146 ( .A1(n99235), .A2(n120470), .B1(n120654), .B2(n120464), 
        .ZN(n6599) );
  OAI22_X1 U87147 ( .A1(n99234), .A2(n120470), .B1(n120657), .B2(n120464), 
        .ZN(n6600) );
  OAI22_X1 U87148 ( .A1(n99233), .A2(n120470), .B1(n120660), .B2(n120464), 
        .ZN(n6601) );
  OAI22_X1 U87149 ( .A1(n99232), .A2(n120471), .B1(n120663), .B2(n120464), 
        .ZN(n6602) );
  OAI22_X1 U87150 ( .A1(n99231), .A2(n120471), .B1(n120666), .B2(n120465), 
        .ZN(n6603) );
  OAI22_X1 U87151 ( .A1(n99230), .A2(n120471), .B1(n120669), .B2(n120465), 
        .ZN(n6604) );
  OAI22_X1 U87152 ( .A1(n99229), .A2(n120471), .B1(n120672), .B2(n120465), 
        .ZN(n6605) );
  OAI22_X1 U87153 ( .A1(n99228), .A2(n120471), .B1(n120675), .B2(n120465), 
        .ZN(n6606) );
  OAI22_X1 U87154 ( .A1(n99227), .A2(n120471), .B1(n120678), .B2(n120465), 
        .ZN(n6607) );
  OAI22_X1 U87155 ( .A1(n99226), .A2(n120471), .B1(n120681), .B2(n120465), 
        .ZN(n6608) );
  OAI22_X1 U87156 ( .A1(n99225), .A2(n120471), .B1(n120684), .B2(n120465), 
        .ZN(n6609) );
  OAI22_X1 U87157 ( .A1(n99224), .A2(n120471), .B1(n120687), .B2(n120465), 
        .ZN(n6610) );
  OAI22_X1 U87158 ( .A1(n99223), .A2(n120471), .B1(n120690), .B2(n120465), 
        .ZN(n6611) );
  OAI22_X1 U87159 ( .A1(n99222), .A2(n120471), .B1(n120693), .B2(n120465), 
        .ZN(n6612) );
  OAI22_X1 U87160 ( .A1(n99221), .A2(n120471), .B1(n120696), .B2(n120465), 
        .ZN(n6613) );
  OAI22_X1 U87161 ( .A1(n99220), .A2(n120472), .B1(n120699), .B2(n120465), 
        .ZN(n6614) );
  OAI22_X1 U87162 ( .A1(n99219), .A2(n120472), .B1(n120702), .B2(n120466), 
        .ZN(n6615) );
  OAI22_X1 U87163 ( .A1(n99218), .A2(n120472), .B1(n120705), .B2(n120466), 
        .ZN(n6616) );
  OAI22_X1 U87164 ( .A1(n99217), .A2(n120472), .B1(n120708), .B2(n120466), 
        .ZN(n6617) );
  OAI22_X1 U87165 ( .A1(n99216), .A2(n120472), .B1(n120711), .B2(n120466), 
        .ZN(n6618) );
  OAI22_X1 U87166 ( .A1(n99215), .A2(n120472), .B1(n120714), .B2(n120466), 
        .ZN(n6619) );
  OAI22_X1 U87167 ( .A1(n99214), .A2(n120472), .B1(n120717), .B2(n120466), 
        .ZN(n6620) );
  OAI22_X1 U87168 ( .A1(n99213), .A2(n120472), .B1(n120720), .B2(n120466), 
        .ZN(n6621) );
  OAI22_X1 U87169 ( .A1(n99212), .A2(n120472), .B1(n120723), .B2(n120466), 
        .ZN(n6622) );
  OAI22_X1 U87170 ( .A1(n99211), .A2(n120472), .B1(n120726), .B2(n120466), 
        .ZN(n6623) );
  OAI22_X1 U87171 ( .A1(n99210), .A2(n120472), .B1(n120729), .B2(n120466), 
        .ZN(n6624) );
  OAI22_X1 U87172 ( .A1(n99209), .A2(n120472), .B1(n120732), .B2(n120466), 
        .ZN(n6625) );
  OAI22_X1 U87173 ( .A1(n99208), .A2(n120473), .B1(n120735), .B2(n120466), 
        .ZN(n6626) );
  OAI22_X1 U87174 ( .A1(n99207), .A2(n120473), .B1(n120738), .B2(n120467), 
        .ZN(n6627) );
  OAI22_X1 U87175 ( .A1(n99206), .A2(n120473), .B1(n120741), .B2(n120467), 
        .ZN(n6628) );
  OAI22_X1 U87176 ( .A1(n99205), .A2(n120473), .B1(n120744), .B2(n120467), 
        .ZN(n6629) );
  OAI22_X1 U87177 ( .A1(n99204), .A2(n120473), .B1(n120747), .B2(n120467), 
        .ZN(n6630) );
  OAI22_X1 U87178 ( .A1(n99203), .A2(n120473), .B1(n120750), .B2(n120467), 
        .ZN(n6631) );
  OAI22_X1 U87179 ( .A1(n99202), .A2(n120473), .B1(n120753), .B2(n120467), 
        .ZN(n6632) );
  OAI22_X1 U87180 ( .A1(n99201), .A2(n120473), .B1(n120756), .B2(n120467), 
        .ZN(n6633) );
  OAI22_X1 U87181 ( .A1(n99200), .A2(n120473), .B1(n120759), .B2(n120467), 
        .ZN(n6634) );
  OAI22_X1 U87182 ( .A1(n99199), .A2(n120473), .B1(n120762), .B2(n120467), 
        .ZN(n6635) );
  OAI22_X1 U87183 ( .A1(n99198), .A2(n120473), .B1(n120765), .B2(n120467), 
        .ZN(n6636) );
  OAI22_X1 U87184 ( .A1(n99197), .A2(n120473), .B1(n120768), .B2(n120467), 
        .ZN(n6637) );
  OAI22_X1 U87185 ( .A1(n99196), .A2(n120474), .B1(n120771), .B2(n120467), 
        .ZN(n6638) );
  OAI22_X1 U87186 ( .A1(n99195), .A2(n120474), .B1(n120774), .B2(n120468), 
        .ZN(n6639) );
  OAI22_X1 U87187 ( .A1(n99194), .A2(n120474), .B1(n120777), .B2(n120468), 
        .ZN(n6640) );
  OAI22_X1 U87188 ( .A1(n99193), .A2(n120474), .B1(n120780), .B2(n120468), 
        .ZN(n6641) );
  OAI22_X1 U87189 ( .A1(n99192), .A2(n120474), .B1(n120783), .B2(n120468), 
        .ZN(n6642) );
  OAI22_X1 U87190 ( .A1(n99191), .A2(n120474), .B1(n120786), .B2(n120468), 
        .ZN(n6643) );
  OAI22_X1 U87191 ( .A1(n99190), .A2(n120474), .B1(n120789), .B2(n120468), 
        .ZN(n6644) );
  OAI22_X1 U87192 ( .A1(n99189), .A2(n120474), .B1(n120792), .B2(n120468), 
        .ZN(n6645) );
  OAI22_X1 U87193 ( .A1(n99188), .A2(n120474), .B1(n120795), .B2(n120468), 
        .ZN(n6646) );
  OAI22_X1 U87194 ( .A1(n99187), .A2(n120474), .B1(n120798), .B2(n120468), 
        .ZN(n6647) );
  OAI22_X1 U87195 ( .A1(n99186), .A2(n120474), .B1(n120801), .B2(n120468), 
        .ZN(n6648) );
  OAI22_X1 U87196 ( .A1(n99185), .A2(n120474), .B1(n120804), .B2(n120468), 
        .ZN(n6649) );
  OAI22_X1 U87197 ( .A1(n99184), .A2(n120475), .B1(n120807), .B2(n120468), 
        .ZN(n6650) );
  OAI22_X1 U87198 ( .A1(n99375), .A2(n120446), .B1(n120630), .B2(n120440), 
        .ZN(n6463) );
  OAI22_X1 U87199 ( .A1(n99374), .A2(n120446), .B1(n120633), .B2(n120440), 
        .ZN(n6464) );
  OAI22_X1 U87200 ( .A1(n99373), .A2(n120446), .B1(n120636), .B2(n120440), 
        .ZN(n6465) );
  OAI22_X1 U87201 ( .A1(n99372), .A2(n120446), .B1(n120639), .B2(n120440), 
        .ZN(n6466) );
  OAI22_X1 U87202 ( .A1(n99371), .A2(n120446), .B1(n120642), .B2(n120440), 
        .ZN(n6467) );
  OAI22_X1 U87203 ( .A1(n99370), .A2(n120446), .B1(n120645), .B2(n120440), 
        .ZN(n6468) );
  OAI22_X1 U87204 ( .A1(n99369), .A2(n120446), .B1(n120648), .B2(n120440), 
        .ZN(n6469) );
  OAI22_X1 U87205 ( .A1(n99368), .A2(n120446), .B1(n120651), .B2(n120440), 
        .ZN(n6470) );
  OAI22_X1 U87206 ( .A1(n99367), .A2(n120446), .B1(n120654), .B2(n120440), 
        .ZN(n6471) );
  OAI22_X1 U87207 ( .A1(n99366), .A2(n120446), .B1(n120657), .B2(n120440), 
        .ZN(n6472) );
  OAI22_X1 U87208 ( .A1(n99365), .A2(n120446), .B1(n120660), .B2(n120440), 
        .ZN(n6473) );
  OAI22_X1 U87209 ( .A1(n99364), .A2(n120447), .B1(n120663), .B2(n120440), 
        .ZN(n6474) );
  OAI22_X1 U87210 ( .A1(n99363), .A2(n120447), .B1(n120666), .B2(n120441), 
        .ZN(n6475) );
  OAI22_X1 U87211 ( .A1(n99362), .A2(n120447), .B1(n120669), .B2(n120441), 
        .ZN(n6476) );
  OAI22_X1 U87212 ( .A1(n99361), .A2(n120447), .B1(n120672), .B2(n120441), 
        .ZN(n6477) );
  OAI22_X1 U87213 ( .A1(n99360), .A2(n120447), .B1(n120675), .B2(n120441), 
        .ZN(n6478) );
  OAI22_X1 U87214 ( .A1(n99359), .A2(n120447), .B1(n120678), .B2(n120441), 
        .ZN(n6479) );
  OAI22_X1 U87215 ( .A1(n99358), .A2(n120447), .B1(n120681), .B2(n120441), 
        .ZN(n6480) );
  OAI22_X1 U87216 ( .A1(n99357), .A2(n120447), .B1(n120684), .B2(n120441), 
        .ZN(n6481) );
  OAI22_X1 U87217 ( .A1(n99356), .A2(n120447), .B1(n120687), .B2(n120441), 
        .ZN(n6482) );
  OAI22_X1 U87218 ( .A1(n99355), .A2(n120447), .B1(n120690), .B2(n120441), 
        .ZN(n6483) );
  OAI22_X1 U87219 ( .A1(n99354), .A2(n120447), .B1(n120693), .B2(n120441), 
        .ZN(n6484) );
  OAI22_X1 U87220 ( .A1(n99353), .A2(n120447), .B1(n120696), .B2(n120441), 
        .ZN(n6485) );
  OAI22_X1 U87221 ( .A1(n99352), .A2(n120448), .B1(n120699), .B2(n120441), 
        .ZN(n6486) );
  OAI22_X1 U87222 ( .A1(n99351), .A2(n120448), .B1(n120702), .B2(n120442), 
        .ZN(n6487) );
  OAI22_X1 U87223 ( .A1(n99350), .A2(n120448), .B1(n120705), .B2(n120442), 
        .ZN(n6488) );
  OAI22_X1 U87224 ( .A1(n99349), .A2(n120448), .B1(n120708), .B2(n120442), 
        .ZN(n6489) );
  OAI22_X1 U87225 ( .A1(n99348), .A2(n120448), .B1(n120711), .B2(n120442), 
        .ZN(n6490) );
  OAI22_X1 U87226 ( .A1(n99347), .A2(n120448), .B1(n120714), .B2(n120442), 
        .ZN(n6491) );
  OAI22_X1 U87227 ( .A1(n99346), .A2(n120448), .B1(n120717), .B2(n120442), 
        .ZN(n6492) );
  OAI22_X1 U87228 ( .A1(n99345), .A2(n120448), .B1(n120720), .B2(n120442), 
        .ZN(n6493) );
  OAI22_X1 U87229 ( .A1(n99344), .A2(n120448), .B1(n120723), .B2(n120442), 
        .ZN(n6494) );
  OAI22_X1 U87230 ( .A1(n99343), .A2(n120448), .B1(n120726), .B2(n120442), 
        .ZN(n6495) );
  OAI22_X1 U87231 ( .A1(n99342), .A2(n120448), .B1(n120729), .B2(n120442), 
        .ZN(n6496) );
  OAI22_X1 U87232 ( .A1(n99341), .A2(n120448), .B1(n120732), .B2(n120442), 
        .ZN(n6497) );
  OAI22_X1 U87233 ( .A1(n99340), .A2(n120449), .B1(n120735), .B2(n120442), 
        .ZN(n6498) );
  OAI22_X1 U87234 ( .A1(n99339), .A2(n120449), .B1(n120738), .B2(n120443), 
        .ZN(n6499) );
  OAI22_X1 U87235 ( .A1(n99338), .A2(n120449), .B1(n120741), .B2(n120443), 
        .ZN(n6500) );
  OAI22_X1 U87236 ( .A1(n99337), .A2(n120449), .B1(n120744), .B2(n120443), 
        .ZN(n6501) );
  OAI22_X1 U87237 ( .A1(n99336), .A2(n120449), .B1(n120747), .B2(n120443), 
        .ZN(n6502) );
  OAI22_X1 U87238 ( .A1(n99335), .A2(n120449), .B1(n120750), .B2(n120443), 
        .ZN(n6503) );
  OAI22_X1 U87239 ( .A1(n99334), .A2(n120449), .B1(n120753), .B2(n120443), 
        .ZN(n6504) );
  OAI22_X1 U87240 ( .A1(n99333), .A2(n120449), .B1(n120756), .B2(n120443), 
        .ZN(n6505) );
  OAI22_X1 U87241 ( .A1(n99332), .A2(n120449), .B1(n120759), .B2(n120443), 
        .ZN(n6506) );
  OAI22_X1 U87242 ( .A1(n99331), .A2(n120449), .B1(n120762), .B2(n120443), 
        .ZN(n6507) );
  OAI22_X1 U87243 ( .A1(n99330), .A2(n120449), .B1(n120765), .B2(n120443), 
        .ZN(n6508) );
  OAI22_X1 U87244 ( .A1(n99329), .A2(n120449), .B1(n120768), .B2(n120443), 
        .ZN(n6509) );
  OAI22_X1 U87245 ( .A1(n99328), .A2(n120450), .B1(n120771), .B2(n120443), 
        .ZN(n6510) );
  OAI22_X1 U87246 ( .A1(n99327), .A2(n120450), .B1(n120774), .B2(n120444), 
        .ZN(n6511) );
  OAI22_X1 U87247 ( .A1(n99326), .A2(n120450), .B1(n120777), .B2(n120444), 
        .ZN(n6512) );
  OAI22_X1 U87248 ( .A1(n99325), .A2(n120450), .B1(n120780), .B2(n120444), 
        .ZN(n6513) );
  OAI22_X1 U87249 ( .A1(n99324), .A2(n120450), .B1(n120783), .B2(n120444), 
        .ZN(n6514) );
  OAI22_X1 U87250 ( .A1(n99323), .A2(n120450), .B1(n120786), .B2(n120444), 
        .ZN(n6515) );
  OAI22_X1 U87251 ( .A1(n99322), .A2(n120450), .B1(n120789), .B2(n120444), 
        .ZN(n6516) );
  OAI22_X1 U87252 ( .A1(n99321), .A2(n120450), .B1(n120792), .B2(n120444), 
        .ZN(n6517) );
  OAI22_X1 U87253 ( .A1(n99320), .A2(n120450), .B1(n120795), .B2(n120444), 
        .ZN(n6518) );
  OAI22_X1 U87254 ( .A1(n99319), .A2(n120450), .B1(n120798), .B2(n120444), 
        .ZN(n6519) );
  OAI22_X1 U87255 ( .A1(n99318), .A2(n120450), .B1(n120801), .B2(n120444), 
        .ZN(n6520) );
  OAI22_X1 U87256 ( .A1(n99317), .A2(n120450), .B1(n120804), .B2(n120444), 
        .ZN(n6521) );
  OAI22_X1 U87257 ( .A1(n99316), .A2(n120451), .B1(n120807), .B2(n120444), 
        .ZN(n6522) );
  OAI22_X1 U87258 ( .A1(n120520), .A2(n114120), .B1(n120629), .B2(n120512), 
        .ZN(n6847) );
  OAI22_X1 U87259 ( .A1(n120520), .A2(n114119), .B1(n120632), .B2(n120512), 
        .ZN(n6848) );
  OAI22_X1 U87260 ( .A1(n120520), .A2(n114118), .B1(n120635), .B2(n120512), 
        .ZN(n6849) );
  OAI22_X1 U87261 ( .A1(n120520), .A2(n114117), .B1(n120638), .B2(n120512), 
        .ZN(n6850) );
  OAI22_X1 U87262 ( .A1(n120520), .A2(n114116), .B1(n120641), .B2(n120512), 
        .ZN(n6851) );
  OAI22_X1 U87263 ( .A1(n120520), .A2(n114115), .B1(n120644), .B2(n120512), 
        .ZN(n6852) );
  OAI22_X1 U87264 ( .A1(n120520), .A2(n114114), .B1(n120647), .B2(n120512), 
        .ZN(n6853) );
  OAI22_X1 U87265 ( .A1(n120520), .A2(n114113), .B1(n120650), .B2(n120512), 
        .ZN(n6854) );
  OAI22_X1 U87266 ( .A1(n120520), .A2(n114112), .B1(n120653), .B2(n120512), 
        .ZN(n6855) );
  OAI22_X1 U87267 ( .A1(n120520), .A2(n114111), .B1(n120656), .B2(n120512), 
        .ZN(n6856) );
  OAI22_X1 U87268 ( .A1(n120520), .A2(n114110), .B1(n120659), .B2(n120512), 
        .ZN(n6857) );
  OAI22_X1 U87269 ( .A1(n120520), .A2(n114109), .B1(n120662), .B2(n120512), 
        .ZN(n6858) );
  OAI22_X1 U87270 ( .A1(n120521), .A2(n114108), .B1(n120665), .B2(n120513), 
        .ZN(n6859) );
  OAI22_X1 U87271 ( .A1(n120521), .A2(n114107), .B1(n120668), .B2(n120513), 
        .ZN(n6860) );
  OAI22_X1 U87272 ( .A1(n120521), .A2(n114106), .B1(n120671), .B2(n120513), 
        .ZN(n6861) );
  OAI22_X1 U87273 ( .A1(n120521), .A2(n114105), .B1(n120674), .B2(n120513), 
        .ZN(n6862) );
  OAI22_X1 U87274 ( .A1(n120521), .A2(n114104), .B1(n120677), .B2(n120513), 
        .ZN(n6863) );
  OAI22_X1 U87275 ( .A1(n120521), .A2(n114103), .B1(n120680), .B2(n120513), 
        .ZN(n6864) );
  OAI22_X1 U87276 ( .A1(n120521), .A2(n114102), .B1(n120683), .B2(n120513), 
        .ZN(n6865) );
  OAI22_X1 U87277 ( .A1(n120521), .A2(n114101), .B1(n120686), .B2(n120513), 
        .ZN(n6866) );
  OAI22_X1 U87278 ( .A1(n120521), .A2(n114100), .B1(n120689), .B2(n120513), 
        .ZN(n6867) );
  OAI22_X1 U87279 ( .A1(n120521), .A2(n114099), .B1(n120692), .B2(n120513), 
        .ZN(n6868) );
  OAI22_X1 U87280 ( .A1(n120521), .A2(n114098), .B1(n120695), .B2(n120513), 
        .ZN(n6869) );
  OAI22_X1 U87281 ( .A1(n120521), .A2(n114097), .B1(n120698), .B2(n120513), 
        .ZN(n6870) );
  OAI22_X1 U87282 ( .A1(n120521), .A2(n114096), .B1(n120701), .B2(n120514), 
        .ZN(n6871) );
  OAI22_X1 U87283 ( .A1(n120522), .A2(n114095), .B1(n120704), .B2(n120514), 
        .ZN(n6872) );
  OAI22_X1 U87284 ( .A1(n120522), .A2(n114094), .B1(n120707), .B2(n120514), 
        .ZN(n6873) );
  OAI22_X1 U87285 ( .A1(n120522), .A2(n114093), .B1(n120710), .B2(n120514), 
        .ZN(n6874) );
  OAI22_X1 U87286 ( .A1(n120522), .A2(n114092), .B1(n120713), .B2(n120514), 
        .ZN(n6875) );
  OAI22_X1 U87287 ( .A1(n120522), .A2(n114091), .B1(n120716), .B2(n120514), 
        .ZN(n6876) );
  OAI22_X1 U87288 ( .A1(n120522), .A2(n114090), .B1(n120719), .B2(n120514), 
        .ZN(n6877) );
  OAI22_X1 U87289 ( .A1(n120522), .A2(n114089), .B1(n120722), .B2(n120514), 
        .ZN(n6878) );
  OAI22_X1 U87290 ( .A1(n120522), .A2(n114088), .B1(n120725), .B2(n120514), 
        .ZN(n6879) );
  OAI22_X1 U87291 ( .A1(n120522), .A2(n114087), .B1(n120728), .B2(n120514), 
        .ZN(n6880) );
  OAI22_X1 U87292 ( .A1(n120522), .A2(n114086), .B1(n120731), .B2(n120514), 
        .ZN(n6881) );
  OAI22_X1 U87293 ( .A1(n120522), .A2(n114085), .B1(n120734), .B2(n120514), 
        .ZN(n6882) );
  OAI22_X1 U87294 ( .A1(n120522), .A2(n114084), .B1(n120737), .B2(n120515), 
        .ZN(n6883) );
  OAI22_X1 U87295 ( .A1(n120522), .A2(n114083), .B1(n120740), .B2(n120515), 
        .ZN(n6884) );
  OAI22_X1 U87296 ( .A1(n120523), .A2(n114082), .B1(n120743), .B2(n120515), 
        .ZN(n6885) );
  OAI22_X1 U87297 ( .A1(n120523), .A2(n114081), .B1(n120746), .B2(n120515), 
        .ZN(n6886) );
  OAI22_X1 U87298 ( .A1(n120523), .A2(n114080), .B1(n120749), .B2(n120515), 
        .ZN(n6887) );
  OAI22_X1 U87299 ( .A1(n120523), .A2(n114079), .B1(n120752), .B2(n120515), 
        .ZN(n6888) );
  OAI22_X1 U87300 ( .A1(n120523), .A2(n114078), .B1(n120755), .B2(n120515), 
        .ZN(n6889) );
  OAI22_X1 U87301 ( .A1(n120523), .A2(n114077), .B1(n120758), .B2(n120515), 
        .ZN(n6890) );
  OAI22_X1 U87302 ( .A1(n120523), .A2(n114076), .B1(n120761), .B2(n120515), 
        .ZN(n6891) );
  OAI22_X1 U87303 ( .A1(n120523), .A2(n114075), .B1(n120764), .B2(n120515), 
        .ZN(n6892) );
  OAI22_X1 U87304 ( .A1(n120523), .A2(n114074), .B1(n120767), .B2(n120515), 
        .ZN(n6893) );
  OAI22_X1 U87305 ( .A1(n120523), .A2(n114073), .B1(n120770), .B2(n120515), 
        .ZN(n6894) );
  OAI22_X1 U87306 ( .A1(n120523), .A2(n114072), .B1(n120773), .B2(n120516), 
        .ZN(n6895) );
  OAI22_X1 U87307 ( .A1(n120523), .A2(n114071), .B1(n120776), .B2(n120516), 
        .ZN(n6896) );
  OAI22_X1 U87308 ( .A1(n120523), .A2(n114070), .B1(n120779), .B2(n120516), 
        .ZN(n6897) );
  OAI22_X1 U87309 ( .A1(n120524), .A2(n114069), .B1(n120782), .B2(n120516), 
        .ZN(n6898) );
  OAI22_X1 U87310 ( .A1(n120524), .A2(n114068), .B1(n120785), .B2(n120516), 
        .ZN(n6899) );
  OAI22_X1 U87311 ( .A1(n120524), .A2(n114067), .B1(n120788), .B2(n120516), 
        .ZN(n6900) );
  OAI22_X1 U87312 ( .A1(n120524), .A2(n114066), .B1(n120791), .B2(n120516), 
        .ZN(n6901) );
  OAI22_X1 U87313 ( .A1(n120524), .A2(n114065), .B1(n120794), .B2(n120516), 
        .ZN(n6902) );
  OAI22_X1 U87314 ( .A1(n120524), .A2(n114064), .B1(n120797), .B2(n120516), 
        .ZN(n6903) );
  OAI22_X1 U87315 ( .A1(n120524), .A2(n114063), .B1(n120800), .B2(n120516), 
        .ZN(n6904) );
  OAI22_X1 U87316 ( .A1(n120524), .A2(n114062), .B1(n120803), .B2(n120516), 
        .ZN(n6905) );
  OAI22_X1 U87317 ( .A1(n120524), .A2(n114061), .B1(n120806), .B2(n120516), 
        .ZN(n6906) );
  OAI22_X1 U87318 ( .A1(n99111), .A2(n120494), .B1(n120629), .B2(n120488), 
        .ZN(n6719) );
  OAI22_X1 U87319 ( .A1(n99110), .A2(n120494), .B1(n120632), .B2(n120488), 
        .ZN(n6720) );
  OAI22_X1 U87320 ( .A1(n99109), .A2(n120494), .B1(n120635), .B2(n120488), 
        .ZN(n6721) );
  OAI22_X1 U87321 ( .A1(n99108), .A2(n120494), .B1(n120638), .B2(n120488), 
        .ZN(n6722) );
  OAI22_X1 U87322 ( .A1(n99107), .A2(n120494), .B1(n120641), .B2(n120488), 
        .ZN(n6723) );
  OAI22_X1 U87323 ( .A1(n99106), .A2(n120494), .B1(n120644), .B2(n120488), 
        .ZN(n6724) );
  OAI22_X1 U87324 ( .A1(n99105), .A2(n120494), .B1(n120647), .B2(n120488), 
        .ZN(n6725) );
  OAI22_X1 U87325 ( .A1(n99104), .A2(n120494), .B1(n120650), .B2(n120488), 
        .ZN(n6726) );
  OAI22_X1 U87326 ( .A1(n99103), .A2(n120494), .B1(n120653), .B2(n120488), 
        .ZN(n6727) );
  OAI22_X1 U87327 ( .A1(n99102), .A2(n120494), .B1(n120656), .B2(n120488), 
        .ZN(n6728) );
  OAI22_X1 U87328 ( .A1(n99101), .A2(n120494), .B1(n120659), .B2(n120488), 
        .ZN(n6729) );
  OAI22_X1 U87329 ( .A1(n99100), .A2(n120495), .B1(n120662), .B2(n120488), 
        .ZN(n6730) );
  OAI22_X1 U87330 ( .A1(n99099), .A2(n120495), .B1(n120665), .B2(n120489), 
        .ZN(n6731) );
  OAI22_X1 U87331 ( .A1(n99098), .A2(n120495), .B1(n120668), .B2(n120489), 
        .ZN(n6732) );
  OAI22_X1 U87332 ( .A1(n99097), .A2(n120495), .B1(n120671), .B2(n120489), 
        .ZN(n6733) );
  OAI22_X1 U87333 ( .A1(n99096), .A2(n120495), .B1(n120674), .B2(n120489), 
        .ZN(n6734) );
  OAI22_X1 U87334 ( .A1(n99095), .A2(n120495), .B1(n120677), .B2(n120489), 
        .ZN(n6735) );
  OAI22_X1 U87335 ( .A1(n99094), .A2(n120495), .B1(n120680), .B2(n120489), 
        .ZN(n6736) );
  OAI22_X1 U87336 ( .A1(n99093), .A2(n120495), .B1(n120683), .B2(n120489), 
        .ZN(n6737) );
  OAI22_X1 U87337 ( .A1(n99092), .A2(n120495), .B1(n120686), .B2(n120489), 
        .ZN(n6738) );
  OAI22_X1 U87338 ( .A1(n99091), .A2(n120495), .B1(n120689), .B2(n120489), 
        .ZN(n6739) );
  OAI22_X1 U87339 ( .A1(n99090), .A2(n120495), .B1(n120692), .B2(n120489), 
        .ZN(n6740) );
  OAI22_X1 U87340 ( .A1(n99089), .A2(n120495), .B1(n120695), .B2(n120489), 
        .ZN(n6741) );
  OAI22_X1 U87341 ( .A1(n99088), .A2(n120496), .B1(n120698), .B2(n120489), 
        .ZN(n6742) );
  OAI22_X1 U87342 ( .A1(n99087), .A2(n120496), .B1(n120701), .B2(n120490), 
        .ZN(n6743) );
  OAI22_X1 U87343 ( .A1(n99086), .A2(n120496), .B1(n120704), .B2(n120490), 
        .ZN(n6744) );
  OAI22_X1 U87344 ( .A1(n99085), .A2(n120496), .B1(n120707), .B2(n120490), 
        .ZN(n6745) );
  OAI22_X1 U87345 ( .A1(n99084), .A2(n120496), .B1(n120710), .B2(n120490), 
        .ZN(n6746) );
  OAI22_X1 U87346 ( .A1(n99083), .A2(n120496), .B1(n120713), .B2(n120490), 
        .ZN(n6747) );
  OAI22_X1 U87347 ( .A1(n99082), .A2(n120496), .B1(n120716), .B2(n120490), 
        .ZN(n6748) );
  OAI22_X1 U87348 ( .A1(n99081), .A2(n120496), .B1(n120719), .B2(n120490), 
        .ZN(n6749) );
  OAI22_X1 U87349 ( .A1(n99080), .A2(n120496), .B1(n120722), .B2(n120490), 
        .ZN(n6750) );
  OAI22_X1 U87350 ( .A1(n99079), .A2(n120496), .B1(n120725), .B2(n120490), 
        .ZN(n6751) );
  OAI22_X1 U87351 ( .A1(n99078), .A2(n120496), .B1(n120728), .B2(n120490), 
        .ZN(n6752) );
  OAI22_X1 U87352 ( .A1(n99077), .A2(n120496), .B1(n120731), .B2(n120490), 
        .ZN(n6753) );
  OAI22_X1 U87353 ( .A1(n99076), .A2(n120497), .B1(n120734), .B2(n120490), 
        .ZN(n6754) );
  OAI22_X1 U87354 ( .A1(n99075), .A2(n120497), .B1(n120737), .B2(n120491), 
        .ZN(n6755) );
  OAI22_X1 U87355 ( .A1(n99074), .A2(n120497), .B1(n120740), .B2(n120491), 
        .ZN(n6756) );
  OAI22_X1 U87356 ( .A1(n99073), .A2(n120497), .B1(n120743), .B2(n120491), 
        .ZN(n6757) );
  OAI22_X1 U87357 ( .A1(n99072), .A2(n120497), .B1(n120746), .B2(n120491), 
        .ZN(n6758) );
  OAI22_X1 U87358 ( .A1(n99071), .A2(n120497), .B1(n120749), .B2(n120491), 
        .ZN(n6759) );
  OAI22_X1 U87359 ( .A1(n99070), .A2(n120497), .B1(n120752), .B2(n120491), 
        .ZN(n6760) );
  OAI22_X1 U87360 ( .A1(n99069), .A2(n120497), .B1(n120755), .B2(n120491), 
        .ZN(n6761) );
  OAI22_X1 U87361 ( .A1(n99068), .A2(n120497), .B1(n120758), .B2(n120491), 
        .ZN(n6762) );
  OAI22_X1 U87362 ( .A1(n99067), .A2(n120497), .B1(n120761), .B2(n120491), 
        .ZN(n6763) );
  OAI22_X1 U87363 ( .A1(n99066), .A2(n120497), .B1(n120764), .B2(n120491), 
        .ZN(n6764) );
  OAI22_X1 U87364 ( .A1(n99065), .A2(n120497), .B1(n120767), .B2(n120491), 
        .ZN(n6765) );
  OAI22_X1 U87365 ( .A1(n99064), .A2(n120498), .B1(n120770), .B2(n120491), 
        .ZN(n6766) );
  OAI22_X1 U87366 ( .A1(n99063), .A2(n120498), .B1(n120773), .B2(n120492), 
        .ZN(n6767) );
  OAI22_X1 U87367 ( .A1(n99062), .A2(n120498), .B1(n120776), .B2(n120492), 
        .ZN(n6768) );
  OAI22_X1 U87368 ( .A1(n99061), .A2(n120498), .B1(n120779), .B2(n120492), 
        .ZN(n6769) );
  OAI22_X1 U87369 ( .A1(n99060), .A2(n120498), .B1(n120782), .B2(n120492), 
        .ZN(n6770) );
  OAI22_X1 U87370 ( .A1(n99059), .A2(n120498), .B1(n120785), .B2(n120492), 
        .ZN(n6771) );
  OAI22_X1 U87371 ( .A1(n99058), .A2(n120498), .B1(n120788), .B2(n120492), 
        .ZN(n6772) );
  OAI22_X1 U87372 ( .A1(n99057), .A2(n120498), .B1(n120791), .B2(n120492), 
        .ZN(n6773) );
  OAI22_X1 U87373 ( .A1(n99056), .A2(n120498), .B1(n120794), .B2(n120492), 
        .ZN(n6774) );
  OAI22_X1 U87374 ( .A1(n99055), .A2(n120498), .B1(n120797), .B2(n120492), 
        .ZN(n6775) );
  OAI22_X1 U87375 ( .A1(n99054), .A2(n120498), .B1(n120800), .B2(n120492), 
        .ZN(n6776) );
  OAI22_X1 U87376 ( .A1(n99053), .A2(n120498), .B1(n120803), .B2(n120492), 
        .ZN(n6777) );
  OAI22_X1 U87377 ( .A1(n99052), .A2(n120499), .B1(n120806), .B2(n120492), 
        .ZN(n6778) );
  OAI22_X1 U87378 ( .A1(n99177), .A2(n120482), .B1(n120630), .B2(n120476), 
        .ZN(n6655) );
  OAI22_X1 U87379 ( .A1(n99176), .A2(n120482), .B1(n120633), .B2(n120476), 
        .ZN(n6656) );
  OAI22_X1 U87380 ( .A1(n99175), .A2(n120482), .B1(n120636), .B2(n120476), 
        .ZN(n6657) );
  OAI22_X1 U87381 ( .A1(n99174), .A2(n120482), .B1(n120639), .B2(n120476), 
        .ZN(n6658) );
  OAI22_X1 U87382 ( .A1(n99173), .A2(n120482), .B1(n120642), .B2(n120476), 
        .ZN(n6659) );
  OAI22_X1 U87383 ( .A1(n99172), .A2(n120482), .B1(n120645), .B2(n120476), 
        .ZN(n6660) );
  OAI22_X1 U87384 ( .A1(n99171), .A2(n120482), .B1(n120648), .B2(n120476), 
        .ZN(n6661) );
  OAI22_X1 U87385 ( .A1(n99170), .A2(n120482), .B1(n120651), .B2(n120476), 
        .ZN(n6662) );
  OAI22_X1 U87386 ( .A1(n99169), .A2(n120482), .B1(n120654), .B2(n120476), 
        .ZN(n6663) );
  OAI22_X1 U87387 ( .A1(n99168), .A2(n120482), .B1(n120657), .B2(n120476), 
        .ZN(n6664) );
  OAI22_X1 U87388 ( .A1(n99167), .A2(n120482), .B1(n120660), .B2(n120476), 
        .ZN(n6665) );
  OAI22_X1 U87389 ( .A1(n99166), .A2(n120483), .B1(n120663), .B2(n120476), 
        .ZN(n6666) );
  OAI22_X1 U87390 ( .A1(n99165), .A2(n120483), .B1(n120666), .B2(n120477), 
        .ZN(n6667) );
  OAI22_X1 U87391 ( .A1(n99164), .A2(n120483), .B1(n120669), .B2(n120477), 
        .ZN(n6668) );
  OAI22_X1 U87392 ( .A1(n99163), .A2(n120483), .B1(n120672), .B2(n120477), 
        .ZN(n6669) );
  OAI22_X1 U87393 ( .A1(n99162), .A2(n120483), .B1(n120675), .B2(n120477), 
        .ZN(n6670) );
  OAI22_X1 U87394 ( .A1(n99161), .A2(n120483), .B1(n120678), .B2(n120477), 
        .ZN(n6671) );
  OAI22_X1 U87395 ( .A1(n99160), .A2(n120483), .B1(n120681), .B2(n120477), 
        .ZN(n6672) );
  OAI22_X1 U87396 ( .A1(n99159), .A2(n120483), .B1(n120684), .B2(n120477), 
        .ZN(n6673) );
  OAI22_X1 U87397 ( .A1(n99158), .A2(n120483), .B1(n120687), .B2(n120477), 
        .ZN(n6674) );
  OAI22_X1 U87398 ( .A1(n99157), .A2(n120483), .B1(n120690), .B2(n120477), 
        .ZN(n6675) );
  OAI22_X1 U87399 ( .A1(n99156), .A2(n120483), .B1(n120693), .B2(n120477), 
        .ZN(n6676) );
  OAI22_X1 U87400 ( .A1(n99155), .A2(n120483), .B1(n120696), .B2(n120477), 
        .ZN(n6677) );
  OAI22_X1 U87401 ( .A1(n99154), .A2(n120484), .B1(n120699), .B2(n120477), 
        .ZN(n6678) );
  OAI22_X1 U87402 ( .A1(n99153), .A2(n120484), .B1(n120702), .B2(n120478), 
        .ZN(n6679) );
  OAI22_X1 U87403 ( .A1(n99152), .A2(n120484), .B1(n120705), .B2(n120478), 
        .ZN(n6680) );
  OAI22_X1 U87404 ( .A1(n99151), .A2(n120484), .B1(n120708), .B2(n120478), 
        .ZN(n6681) );
  OAI22_X1 U87405 ( .A1(n99150), .A2(n120484), .B1(n120711), .B2(n120478), 
        .ZN(n6682) );
  OAI22_X1 U87406 ( .A1(n99149), .A2(n120484), .B1(n120714), .B2(n120478), 
        .ZN(n6683) );
  OAI22_X1 U87407 ( .A1(n99148), .A2(n120484), .B1(n120717), .B2(n120478), 
        .ZN(n6684) );
  OAI22_X1 U87408 ( .A1(n99147), .A2(n120484), .B1(n120720), .B2(n120478), 
        .ZN(n6685) );
  OAI22_X1 U87409 ( .A1(n99146), .A2(n120484), .B1(n120723), .B2(n120478), 
        .ZN(n6686) );
  OAI22_X1 U87410 ( .A1(n99145), .A2(n120484), .B1(n120726), .B2(n120478), 
        .ZN(n6687) );
  OAI22_X1 U87411 ( .A1(n99144), .A2(n120484), .B1(n120729), .B2(n120478), 
        .ZN(n6688) );
  OAI22_X1 U87412 ( .A1(n99143), .A2(n120484), .B1(n120732), .B2(n120478), 
        .ZN(n6689) );
  OAI22_X1 U87413 ( .A1(n99142), .A2(n120485), .B1(n120735), .B2(n120478), 
        .ZN(n6690) );
  OAI22_X1 U87414 ( .A1(n99141), .A2(n120485), .B1(n120738), .B2(n120479), 
        .ZN(n6691) );
  OAI22_X1 U87415 ( .A1(n99140), .A2(n120485), .B1(n120741), .B2(n120479), 
        .ZN(n6692) );
  OAI22_X1 U87416 ( .A1(n99139), .A2(n120485), .B1(n120744), .B2(n120479), 
        .ZN(n6693) );
  OAI22_X1 U87417 ( .A1(n99138), .A2(n120485), .B1(n120747), .B2(n120479), 
        .ZN(n6694) );
  OAI22_X1 U87418 ( .A1(n99137), .A2(n120485), .B1(n120750), .B2(n120479), 
        .ZN(n6695) );
  OAI22_X1 U87419 ( .A1(n99136), .A2(n120485), .B1(n120753), .B2(n120479), 
        .ZN(n6696) );
  OAI22_X1 U87420 ( .A1(n99135), .A2(n120485), .B1(n120756), .B2(n120479), 
        .ZN(n6697) );
  OAI22_X1 U87421 ( .A1(n99134), .A2(n120485), .B1(n120759), .B2(n120479), 
        .ZN(n6698) );
  OAI22_X1 U87422 ( .A1(n99133), .A2(n120485), .B1(n120762), .B2(n120479), 
        .ZN(n6699) );
  OAI22_X1 U87423 ( .A1(n99132), .A2(n120485), .B1(n120765), .B2(n120479), 
        .ZN(n6700) );
  OAI22_X1 U87424 ( .A1(n99131), .A2(n120485), .B1(n120768), .B2(n120479), 
        .ZN(n6701) );
  OAI22_X1 U87425 ( .A1(n99130), .A2(n120486), .B1(n120771), .B2(n120479), 
        .ZN(n6702) );
  OAI22_X1 U87426 ( .A1(n99129), .A2(n120486), .B1(n120774), .B2(n120480), 
        .ZN(n6703) );
  OAI22_X1 U87427 ( .A1(n99128), .A2(n120486), .B1(n120777), .B2(n120480), 
        .ZN(n6704) );
  OAI22_X1 U87428 ( .A1(n99127), .A2(n120486), .B1(n120780), .B2(n120480), 
        .ZN(n6705) );
  OAI22_X1 U87429 ( .A1(n99126), .A2(n120486), .B1(n120783), .B2(n120480), 
        .ZN(n6706) );
  OAI22_X1 U87430 ( .A1(n99125), .A2(n120486), .B1(n120786), .B2(n120480), 
        .ZN(n6707) );
  OAI22_X1 U87431 ( .A1(n99124), .A2(n120486), .B1(n120789), .B2(n120480), 
        .ZN(n6708) );
  OAI22_X1 U87432 ( .A1(n99123), .A2(n120486), .B1(n120792), .B2(n120480), 
        .ZN(n6709) );
  OAI22_X1 U87433 ( .A1(n99122), .A2(n120486), .B1(n120795), .B2(n120480), 
        .ZN(n6710) );
  OAI22_X1 U87434 ( .A1(n99121), .A2(n120486), .B1(n120798), .B2(n120480), 
        .ZN(n6711) );
  OAI22_X1 U87435 ( .A1(n99120), .A2(n120486), .B1(n120801), .B2(n120480), 
        .ZN(n6712) );
  OAI22_X1 U87436 ( .A1(n99119), .A2(n120486), .B1(n120804), .B2(n120480), 
        .ZN(n6713) );
  OAI22_X1 U87437 ( .A1(n99118), .A2(n120487), .B1(n120807), .B2(n120480), 
        .ZN(n6714) );
  OAI22_X1 U87438 ( .A1(n99309), .A2(n120458), .B1(n120630), .B2(n120452), 
        .ZN(n6527) );
  OAI22_X1 U87439 ( .A1(n99308), .A2(n120458), .B1(n120633), .B2(n120452), 
        .ZN(n6528) );
  OAI22_X1 U87440 ( .A1(n99307), .A2(n120458), .B1(n120636), .B2(n120452), 
        .ZN(n6529) );
  OAI22_X1 U87441 ( .A1(n99306), .A2(n120458), .B1(n120639), .B2(n120452), 
        .ZN(n6530) );
  OAI22_X1 U87442 ( .A1(n99305), .A2(n120458), .B1(n120642), .B2(n120452), 
        .ZN(n6531) );
  OAI22_X1 U87443 ( .A1(n99304), .A2(n120458), .B1(n120645), .B2(n120452), 
        .ZN(n6532) );
  OAI22_X1 U87444 ( .A1(n99303), .A2(n120458), .B1(n120648), .B2(n120452), 
        .ZN(n6533) );
  OAI22_X1 U87445 ( .A1(n99302), .A2(n120458), .B1(n120651), .B2(n120452), 
        .ZN(n6534) );
  OAI22_X1 U87446 ( .A1(n99301), .A2(n120458), .B1(n120654), .B2(n120452), 
        .ZN(n6535) );
  OAI22_X1 U87447 ( .A1(n99300), .A2(n120458), .B1(n120657), .B2(n120452), 
        .ZN(n6536) );
  OAI22_X1 U87448 ( .A1(n99299), .A2(n120458), .B1(n120660), .B2(n120452), 
        .ZN(n6537) );
  OAI22_X1 U87449 ( .A1(n99298), .A2(n120459), .B1(n120663), .B2(n120452), 
        .ZN(n6538) );
  OAI22_X1 U87450 ( .A1(n99297), .A2(n120459), .B1(n120666), .B2(n120453), 
        .ZN(n6539) );
  OAI22_X1 U87451 ( .A1(n99296), .A2(n120459), .B1(n120669), .B2(n120453), 
        .ZN(n6540) );
  OAI22_X1 U87452 ( .A1(n99295), .A2(n120459), .B1(n120672), .B2(n120453), 
        .ZN(n6541) );
  OAI22_X1 U87453 ( .A1(n99294), .A2(n120459), .B1(n120675), .B2(n120453), 
        .ZN(n6542) );
  OAI22_X1 U87454 ( .A1(n99293), .A2(n120459), .B1(n120678), .B2(n120453), 
        .ZN(n6543) );
  OAI22_X1 U87455 ( .A1(n99292), .A2(n120459), .B1(n120681), .B2(n120453), 
        .ZN(n6544) );
  OAI22_X1 U87456 ( .A1(n99291), .A2(n120459), .B1(n120684), .B2(n120453), 
        .ZN(n6545) );
  OAI22_X1 U87457 ( .A1(n99290), .A2(n120459), .B1(n120687), .B2(n120453), 
        .ZN(n6546) );
  OAI22_X1 U87458 ( .A1(n99289), .A2(n120459), .B1(n120690), .B2(n120453), 
        .ZN(n6547) );
  OAI22_X1 U87459 ( .A1(n99288), .A2(n120459), .B1(n120693), .B2(n120453), 
        .ZN(n6548) );
  OAI22_X1 U87460 ( .A1(n99287), .A2(n120459), .B1(n120696), .B2(n120453), 
        .ZN(n6549) );
  OAI22_X1 U87461 ( .A1(n99286), .A2(n120460), .B1(n120699), .B2(n120453), 
        .ZN(n6550) );
  OAI22_X1 U87462 ( .A1(n99285), .A2(n120460), .B1(n120702), .B2(n120454), 
        .ZN(n6551) );
  OAI22_X1 U87463 ( .A1(n99284), .A2(n120460), .B1(n120705), .B2(n120454), 
        .ZN(n6552) );
  OAI22_X1 U87464 ( .A1(n99283), .A2(n120460), .B1(n120708), .B2(n120454), 
        .ZN(n6553) );
  OAI22_X1 U87465 ( .A1(n99282), .A2(n120460), .B1(n120711), .B2(n120454), 
        .ZN(n6554) );
  OAI22_X1 U87466 ( .A1(n99281), .A2(n120460), .B1(n120714), .B2(n120454), 
        .ZN(n6555) );
  OAI22_X1 U87467 ( .A1(n99280), .A2(n120460), .B1(n120717), .B2(n120454), 
        .ZN(n6556) );
  OAI22_X1 U87468 ( .A1(n99279), .A2(n120460), .B1(n120720), .B2(n120454), 
        .ZN(n6557) );
  OAI22_X1 U87469 ( .A1(n99278), .A2(n120460), .B1(n120723), .B2(n120454), 
        .ZN(n6558) );
  OAI22_X1 U87470 ( .A1(n99277), .A2(n120460), .B1(n120726), .B2(n120454), 
        .ZN(n6559) );
  OAI22_X1 U87471 ( .A1(n99276), .A2(n120460), .B1(n120729), .B2(n120454), 
        .ZN(n6560) );
  OAI22_X1 U87472 ( .A1(n99275), .A2(n120460), .B1(n120732), .B2(n120454), 
        .ZN(n6561) );
  OAI22_X1 U87473 ( .A1(n99274), .A2(n120461), .B1(n120735), .B2(n120454), 
        .ZN(n6562) );
  OAI22_X1 U87474 ( .A1(n99273), .A2(n120461), .B1(n120738), .B2(n120455), 
        .ZN(n6563) );
  OAI22_X1 U87475 ( .A1(n99272), .A2(n120461), .B1(n120741), .B2(n120455), 
        .ZN(n6564) );
  OAI22_X1 U87476 ( .A1(n99271), .A2(n120461), .B1(n120744), .B2(n120455), 
        .ZN(n6565) );
  OAI22_X1 U87477 ( .A1(n99270), .A2(n120461), .B1(n120747), .B2(n120455), 
        .ZN(n6566) );
  OAI22_X1 U87478 ( .A1(n99269), .A2(n120461), .B1(n120750), .B2(n120455), 
        .ZN(n6567) );
  OAI22_X1 U87479 ( .A1(n99268), .A2(n120461), .B1(n120753), .B2(n120455), 
        .ZN(n6568) );
  OAI22_X1 U87480 ( .A1(n99267), .A2(n120461), .B1(n120756), .B2(n120455), 
        .ZN(n6569) );
  OAI22_X1 U87481 ( .A1(n99266), .A2(n120461), .B1(n120759), .B2(n120455), 
        .ZN(n6570) );
  OAI22_X1 U87482 ( .A1(n99265), .A2(n120461), .B1(n120762), .B2(n120455), 
        .ZN(n6571) );
  OAI22_X1 U87483 ( .A1(n99264), .A2(n120461), .B1(n120765), .B2(n120455), 
        .ZN(n6572) );
  OAI22_X1 U87484 ( .A1(n99263), .A2(n120461), .B1(n120768), .B2(n120455), 
        .ZN(n6573) );
  OAI22_X1 U87485 ( .A1(n99262), .A2(n120462), .B1(n120771), .B2(n120455), 
        .ZN(n6574) );
  OAI22_X1 U87486 ( .A1(n99261), .A2(n120462), .B1(n120774), .B2(n120456), 
        .ZN(n6575) );
  OAI22_X1 U87487 ( .A1(n99260), .A2(n120462), .B1(n120777), .B2(n120456), 
        .ZN(n6576) );
  OAI22_X1 U87488 ( .A1(n99259), .A2(n120462), .B1(n120780), .B2(n120456), 
        .ZN(n6577) );
  OAI22_X1 U87489 ( .A1(n99258), .A2(n120462), .B1(n120783), .B2(n120456), 
        .ZN(n6578) );
  OAI22_X1 U87490 ( .A1(n99257), .A2(n120462), .B1(n120786), .B2(n120456), 
        .ZN(n6579) );
  OAI22_X1 U87491 ( .A1(n99256), .A2(n120462), .B1(n120789), .B2(n120456), 
        .ZN(n6580) );
  OAI22_X1 U87492 ( .A1(n99255), .A2(n120462), .B1(n120792), .B2(n120456), 
        .ZN(n6581) );
  OAI22_X1 U87493 ( .A1(n99254), .A2(n120462), .B1(n120795), .B2(n120456), 
        .ZN(n6582) );
  OAI22_X1 U87494 ( .A1(n99253), .A2(n120462), .B1(n120798), .B2(n120456), 
        .ZN(n6583) );
  OAI22_X1 U87495 ( .A1(n99252), .A2(n120462), .B1(n120801), .B2(n120456), 
        .ZN(n6584) );
  OAI22_X1 U87496 ( .A1(n99251), .A2(n120462), .B1(n120804), .B2(n120456), 
        .ZN(n6585) );
  OAI22_X1 U87497 ( .A1(n99250), .A2(n120463), .B1(n120807), .B2(n120456), 
        .ZN(n6586) );
  OAI22_X1 U87498 ( .A1(n98778), .A2(n120581), .B1(n120629), .B2(n120575), 
        .ZN(n7167) );
  OAI22_X1 U87499 ( .A1(n98777), .A2(n120581), .B1(n120632), .B2(n120575), 
        .ZN(n7168) );
  OAI22_X1 U87500 ( .A1(n98776), .A2(n120581), .B1(n120635), .B2(n120575), 
        .ZN(n7169) );
  OAI22_X1 U87501 ( .A1(n98775), .A2(n120581), .B1(n120638), .B2(n120575), 
        .ZN(n7170) );
  OAI22_X1 U87502 ( .A1(n98774), .A2(n120581), .B1(n120641), .B2(n120575), 
        .ZN(n7171) );
  OAI22_X1 U87503 ( .A1(n98773), .A2(n120581), .B1(n120644), .B2(n120575), 
        .ZN(n7172) );
  OAI22_X1 U87504 ( .A1(n98772), .A2(n120581), .B1(n120647), .B2(n120575), 
        .ZN(n7173) );
  OAI22_X1 U87505 ( .A1(n98771), .A2(n120581), .B1(n120650), .B2(n120575), 
        .ZN(n7174) );
  OAI22_X1 U87506 ( .A1(n98770), .A2(n120581), .B1(n120653), .B2(n120575), 
        .ZN(n7175) );
  OAI22_X1 U87507 ( .A1(n98769), .A2(n120581), .B1(n120656), .B2(n120575), 
        .ZN(n7176) );
  OAI22_X1 U87508 ( .A1(n98768), .A2(n120581), .B1(n120659), .B2(n120575), 
        .ZN(n7177) );
  OAI22_X1 U87509 ( .A1(n98767), .A2(n120582), .B1(n120662), .B2(n120575), 
        .ZN(n7178) );
  OAI22_X1 U87510 ( .A1(n98766), .A2(n120582), .B1(n120665), .B2(n120576), 
        .ZN(n7179) );
  OAI22_X1 U87511 ( .A1(n98765), .A2(n120582), .B1(n120668), .B2(n120576), 
        .ZN(n7180) );
  OAI22_X1 U87512 ( .A1(n98764), .A2(n120582), .B1(n120671), .B2(n120576), 
        .ZN(n7181) );
  OAI22_X1 U87513 ( .A1(n98763), .A2(n120582), .B1(n120674), .B2(n120576), 
        .ZN(n7182) );
  OAI22_X1 U87514 ( .A1(n98762), .A2(n120582), .B1(n120677), .B2(n120576), 
        .ZN(n7183) );
  OAI22_X1 U87515 ( .A1(n98761), .A2(n120582), .B1(n120680), .B2(n120576), 
        .ZN(n7184) );
  OAI22_X1 U87516 ( .A1(n98760), .A2(n120582), .B1(n120683), .B2(n120576), 
        .ZN(n7185) );
  OAI22_X1 U87517 ( .A1(n98759), .A2(n120582), .B1(n120686), .B2(n120576), 
        .ZN(n7186) );
  OAI22_X1 U87518 ( .A1(n98758), .A2(n120582), .B1(n120689), .B2(n120576), 
        .ZN(n7187) );
  OAI22_X1 U87519 ( .A1(n98757), .A2(n120582), .B1(n120692), .B2(n120576), 
        .ZN(n7188) );
  OAI22_X1 U87520 ( .A1(n98756), .A2(n120582), .B1(n120695), .B2(n120576), 
        .ZN(n7189) );
  OAI22_X1 U87521 ( .A1(n98755), .A2(n120583), .B1(n120698), .B2(n120576), 
        .ZN(n7190) );
  OAI22_X1 U87522 ( .A1(n98754), .A2(n120583), .B1(n120701), .B2(n120577), 
        .ZN(n7191) );
  OAI22_X1 U87523 ( .A1(n98753), .A2(n120583), .B1(n120704), .B2(n120577), 
        .ZN(n7192) );
  OAI22_X1 U87524 ( .A1(n98752), .A2(n120583), .B1(n120707), .B2(n120577), 
        .ZN(n7193) );
  OAI22_X1 U87525 ( .A1(n98751), .A2(n120583), .B1(n120710), .B2(n120577), 
        .ZN(n7194) );
  OAI22_X1 U87526 ( .A1(n98750), .A2(n120583), .B1(n120713), .B2(n120577), 
        .ZN(n7195) );
  OAI22_X1 U87527 ( .A1(n98749), .A2(n120583), .B1(n120716), .B2(n120577), 
        .ZN(n7196) );
  OAI22_X1 U87528 ( .A1(n98748), .A2(n120583), .B1(n120719), .B2(n120577), 
        .ZN(n7197) );
  OAI22_X1 U87529 ( .A1(n98747), .A2(n120583), .B1(n120722), .B2(n120577), 
        .ZN(n7198) );
  OAI22_X1 U87530 ( .A1(n98746), .A2(n120583), .B1(n120725), .B2(n120577), 
        .ZN(n7199) );
  OAI22_X1 U87531 ( .A1(n98745), .A2(n120583), .B1(n120728), .B2(n120577), 
        .ZN(n7200) );
  OAI22_X1 U87532 ( .A1(n98744), .A2(n120583), .B1(n120731), .B2(n120577), 
        .ZN(n7201) );
  OAI22_X1 U87533 ( .A1(n98743), .A2(n120584), .B1(n120734), .B2(n120577), 
        .ZN(n7202) );
  OAI22_X1 U87534 ( .A1(n98742), .A2(n120584), .B1(n120737), .B2(n120578), 
        .ZN(n7203) );
  OAI22_X1 U87535 ( .A1(n98741), .A2(n120584), .B1(n120740), .B2(n120578), 
        .ZN(n7204) );
  OAI22_X1 U87536 ( .A1(n98740), .A2(n120584), .B1(n120743), .B2(n120578), 
        .ZN(n7205) );
  OAI22_X1 U87537 ( .A1(n98739), .A2(n120584), .B1(n120746), .B2(n120578), 
        .ZN(n7206) );
  OAI22_X1 U87538 ( .A1(n98738), .A2(n120584), .B1(n120749), .B2(n120578), 
        .ZN(n7207) );
  OAI22_X1 U87539 ( .A1(n98737), .A2(n120584), .B1(n120752), .B2(n120578), 
        .ZN(n7208) );
  OAI22_X1 U87540 ( .A1(n98736), .A2(n120584), .B1(n120755), .B2(n120578), 
        .ZN(n7209) );
  OAI22_X1 U87541 ( .A1(n98735), .A2(n120584), .B1(n120758), .B2(n120578), 
        .ZN(n7210) );
  OAI22_X1 U87542 ( .A1(n98734), .A2(n120584), .B1(n120761), .B2(n120578), 
        .ZN(n7211) );
  OAI22_X1 U87543 ( .A1(n98733), .A2(n120584), .B1(n120764), .B2(n120578), 
        .ZN(n7212) );
  OAI22_X1 U87544 ( .A1(n98732), .A2(n120584), .B1(n120767), .B2(n120578), 
        .ZN(n7213) );
  OAI22_X1 U87545 ( .A1(n98731), .A2(n120585), .B1(n120770), .B2(n120578), 
        .ZN(n7214) );
  OAI22_X1 U87546 ( .A1(n98730), .A2(n120585), .B1(n120773), .B2(n120579), 
        .ZN(n7215) );
  OAI22_X1 U87547 ( .A1(n98729), .A2(n120585), .B1(n120776), .B2(n120579), 
        .ZN(n7216) );
  OAI22_X1 U87548 ( .A1(n98728), .A2(n120585), .B1(n120779), .B2(n120579), 
        .ZN(n7217) );
  OAI22_X1 U87549 ( .A1(n98727), .A2(n120585), .B1(n120782), .B2(n120579), 
        .ZN(n7218) );
  OAI22_X1 U87550 ( .A1(n98726), .A2(n120585), .B1(n120785), .B2(n120579), 
        .ZN(n7219) );
  OAI22_X1 U87551 ( .A1(n98725), .A2(n120585), .B1(n120788), .B2(n120579), 
        .ZN(n7220) );
  OAI22_X1 U87552 ( .A1(n98724), .A2(n120585), .B1(n120791), .B2(n120579), 
        .ZN(n7221) );
  OAI22_X1 U87553 ( .A1(n98723), .A2(n120585), .B1(n120794), .B2(n120579), 
        .ZN(n7222) );
  OAI22_X1 U87554 ( .A1(n98722), .A2(n120585), .B1(n120797), .B2(n120579), 
        .ZN(n7223) );
  OAI22_X1 U87555 ( .A1(n98721), .A2(n120585), .B1(n120800), .B2(n120579), 
        .ZN(n7224) );
  OAI22_X1 U87556 ( .A1(n98720), .A2(n120585), .B1(n120803), .B2(n120579), 
        .ZN(n7225) );
  OAI22_X1 U87557 ( .A1(n98719), .A2(n120586), .B1(n120806), .B2(n120579), 
        .ZN(n7226) );
  OAI22_X1 U87558 ( .A1(n99045), .A2(n120506), .B1(n120629), .B2(n120500), 
        .ZN(n6783) );
  OAI22_X1 U87559 ( .A1(n99044), .A2(n120506), .B1(n120632), .B2(n120500), 
        .ZN(n6784) );
  OAI22_X1 U87560 ( .A1(n99043), .A2(n120506), .B1(n120635), .B2(n120500), 
        .ZN(n6785) );
  OAI22_X1 U87561 ( .A1(n99042), .A2(n120506), .B1(n120638), .B2(n120500), 
        .ZN(n6786) );
  OAI22_X1 U87562 ( .A1(n99041), .A2(n120506), .B1(n120641), .B2(n120500), 
        .ZN(n6787) );
  OAI22_X1 U87563 ( .A1(n99040), .A2(n120506), .B1(n120644), .B2(n120500), 
        .ZN(n6788) );
  OAI22_X1 U87564 ( .A1(n99039), .A2(n120506), .B1(n120647), .B2(n120500), 
        .ZN(n6789) );
  OAI22_X1 U87565 ( .A1(n99038), .A2(n120506), .B1(n120650), .B2(n120500), 
        .ZN(n6790) );
  OAI22_X1 U87566 ( .A1(n99037), .A2(n120506), .B1(n120653), .B2(n120500), 
        .ZN(n6791) );
  OAI22_X1 U87567 ( .A1(n99036), .A2(n120506), .B1(n120656), .B2(n120500), 
        .ZN(n6792) );
  OAI22_X1 U87568 ( .A1(n99035), .A2(n120506), .B1(n120659), .B2(n120500), 
        .ZN(n6793) );
  OAI22_X1 U87569 ( .A1(n99034), .A2(n120507), .B1(n120662), .B2(n120500), 
        .ZN(n6794) );
  OAI22_X1 U87570 ( .A1(n99033), .A2(n120507), .B1(n120665), .B2(n120501), 
        .ZN(n6795) );
  OAI22_X1 U87571 ( .A1(n99032), .A2(n120507), .B1(n120668), .B2(n120501), 
        .ZN(n6796) );
  OAI22_X1 U87572 ( .A1(n99031), .A2(n120507), .B1(n120671), .B2(n120501), 
        .ZN(n6797) );
  OAI22_X1 U87573 ( .A1(n99030), .A2(n120507), .B1(n120674), .B2(n120501), 
        .ZN(n6798) );
  OAI22_X1 U87574 ( .A1(n99029), .A2(n120507), .B1(n120677), .B2(n120501), 
        .ZN(n6799) );
  OAI22_X1 U87575 ( .A1(n99028), .A2(n120507), .B1(n120680), .B2(n120501), 
        .ZN(n6800) );
  OAI22_X1 U87576 ( .A1(n99027), .A2(n120507), .B1(n120683), .B2(n120501), 
        .ZN(n6801) );
  OAI22_X1 U87577 ( .A1(n99026), .A2(n120507), .B1(n120686), .B2(n120501), 
        .ZN(n6802) );
  OAI22_X1 U87578 ( .A1(n99025), .A2(n120507), .B1(n120689), .B2(n120501), 
        .ZN(n6803) );
  OAI22_X1 U87579 ( .A1(n99024), .A2(n120507), .B1(n120692), .B2(n120501), 
        .ZN(n6804) );
  OAI22_X1 U87580 ( .A1(n99023), .A2(n120507), .B1(n120695), .B2(n120501), 
        .ZN(n6805) );
  OAI22_X1 U87581 ( .A1(n99022), .A2(n120508), .B1(n120698), .B2(n120501), 
        .ZN(n6806) );
  OAI22_X1 U87582 ( .A1(n99021), .A2(n120508), .B1(n120701), .B2(n120502), 
        .ZN(n6807) );
  OAI22_X1 U87583 ( .A1(n99020), .A2(n120508), .B1(n120704), .B2(n120502), 
        .ZN(n6808) );
  OAI22_X1 U87584 ( .A1(n99019), .A2(n120508), .B1(n120707), .B2(n120502), 
        .ZN(n6809) );
  OAI22_X1 U87585 ( .A1(n99018), .A2(n120508), .B1(n120710), .B2(n120502), 
        .ZN(n6810) );
  OAI22_X1 U87586 ( .A1(n99017), .A2(n120508), .B1(n120713), .B2(n120502), 
        .ZN(n6811) );
  OAI22_X1 U87587 ( .A1(n99016), .A2(n120508), .B1(n120716), .B2(n120502), 
        .ZN(n6812) );
  OAI22_X1 U87588 ( .A1(n99015), .A2(n120508), .B1(n120719), .B2(n120502), 
        .ZN(n6813) );
  OAI22_X1 U87589 ( .A1(n99014), .A2(n120508), .B1(n120722), .B2(n120502), 
        .ZN(n6814) );
  OAI22_X1 U87590 ( .A1(n99013), .A2(n120508), .B1(n120725), .B2(n120502), 
        .ZN(n6815) );
  OAI22_X1 U87591 ( .A1(n99012), .A2(n120508), .B1(n120728), .B2(n120502), 
        .ZN(n6816) );
  OAI22_X1 U87592 ( .A1(n99011), .A2(n120508), .B1(n120731), .B2(n120502), 
        .ZN(n6817) );
  OAI22_X1 U87593 ( .A1(n99010), .A2(n120509), .B1(n120734), .B2(n120502), 
        .ZN(n6818) );
  OAI22_X1 U87594 ( .A1(n99009), .A2(n120509), .B1(n120737), .B2(n120503), 
        .ZN(n6819) );
  OAI22_X1 U87595 ( .A1(n99008), .A2(n120509), .B1(n120740), .B2(n120503), 
        .ZN(n6820) );
  OAI22_X1 U87596 ( .A1(n99007), .A2(n120509), .B1(n120743), .B2(n120503), 
        .ZN(n6821) );
  OAI22_X1 U87597 ( .A1(n99006), .A2(n120509), .B1(n120746), .B2(n120503), 
        .ZN(n6822) );
  OAI22_X1 U87598 ( .A1(n99005), .A2(n120509), .B1(n120749), .B2(n120503), 
        .ZN(n6823) );
  OAI22_X1 U87599 ( .A1(n99004), .A2(n120509), .B1(n120752), .B2(n120503), 
        .ZN(n6824) );
  OAI22_X1 U87600 ( .A1(n99003), .A2(n120509), .B1(n120755), .B2(n120503), 
        .ZN(n6825) );
  OAI22_X1 U87601 ( .A1(n99002), .A2(n120509), .B1(n120758), .B2(n120503), 
        .ZN(n6826) );
  OAI22_X1 U87602 ( .A1(n99001), .A2(n120509), .B1(n120761), .B2(n120503), 
        .ZN(n6827) );
  OAI22_X1 U87603 ( .A1(n99000), .A2(n120509), .B1(n120764), .B2(n120503), 
        .ZN(n6828) );
  OAI22_X1 U87604 ( .A1(n98999), .A2(n120509), .B1(n120767), .B2(n120503), 
        .ZN(n6829) );
  OAI22_X1 U87605 ( .A1(n98998), .A2(n120510), .B1(n120770), .B2(n120503), 
        .ZN(n6830) );
  OAI22_X1 U87606 ( .A1(n98997), .A2(n120510), .B1(n120773), .B2(n120504), 
        .ZN(n6831) );
  OAI22_X1 U87607 ( .A1(n98996), .A2(n120510), .B1(n120776), .B2(n120504), 
        .ZN(n6832) );
  OAI22_X1 U87608 ( .A1(n98995), .A2(n120510), .B1(n120779), .B2(n120504), 
        .ZN(n6833) );
  OAI22_X1 U87609 ( .A1(n98994), .A2(n120510), .B1(n120782), .B2(n120504), 
        .ZN(n6834) );
  OAI22_X1 U87610 ( .A1(n98993), .A2(n120510), .B1(n120785), .B2(n120504), 
        .ZN(n6835) );
  OAI22_X1 U87611 ( .A1(n98992), .A2(n120510), .B1(n120788), .B2(n120504), 
        .ZN(n6836) );
  OAI22_X1 U87612 ( .A1(n98991), .A2(n120510), .B1(n120791), .B2(n120504), 
        .ZN(n6837) );
  OAI22_X1 U87613 ( .A1(n98990), .A2(n120510), .B1(n120794), .B2(n120504), 
        .ZN(n6838) );
  OAI22_X1 U87614 ( .A1(n98989), .A2(n120510), .B1(n120797), .B2(n120504), 
        .ZN(n6839) );
  OAI22_X1 U87615 ( .A1(n98988), .A2(n120510), .B1(n120800), .B2(n120504), 
        .ZN(n6840) );
  OAI22_X1 U87616 ( .A1(n98987), .A2(n120510), .B1(n120803), .B2(n120504), 
        .ZN(n6841) );
  OAI22_X1 U87617 ( .A1(n98986), .A2(n120511), .B1(n120806), .B2(n120504), 
        .ZN(n6842) );
  OAI22_X1 U87618 ( .A1(n98907), .A2(n120556), .B1(n120629), .B2(n120550), 
        .ZN(n7039) );
  OAI22_X1 U87619 ( .A1(n98906), .A2(n120556), .B1(n120632), .B2(n120550), 
        .ZN(n7040) );
  OAI22_X1 U87620 ( .A1(n98905), .A2(n120556), .B1(n120635), .B2(n120550), 
        .ZN(n7041) );
  OAI22_X1 U87621 ( .A1(n98904), .A2(n120556), .B1(n120638), .B2(n120550), 
        .ZN(n7042) );
  OAI22_X1 U87622 ( .A1(n98903), .A2(n120556), .B1(n120641), .B2(n120550), 
        .ZN(n7043) );
  OAI22_X1 U87623 ( .A1(n98902), .A2(n120556), .B1(n120644), .B2(n120550), 
        .ZN(n7044) );
  OAI22_X1 U87624 ( .A1(n98901), .A2(n120556), .B1(n120647), .B2(n120550), 
        .ZN(n7045) );
  OAI22_X1 U87625 ( .A1(n98900), .A2(n120556), .B1(n120650), .B2(n120550), 
        .ZN(n7046) );
  OAI22_X1 U87626 ( .A1(n98899), .A2(n120556), .B1(n120653), .B2(n120550), 
        .ZN(n7047) );
  OAI22_X1 U87627 ( .A1(n98898), .A2(n120556), .B1(n120656), .B2(n120550), 
        .ZN(n7048) );
  OAI22_X1 U87628 ( .A1(n98897), .A2(n120556), .B1(n120659), .B2(n120550), 
        .ZN(n7049) );
  OAI22_X1 U87629 ( .A1(n98896), .A2(n120557), .B1(n120662), .B2(n120550), 
        .ZN(n7050) );
  OAI22_X1 U87630 ( .A1(n98895), .A2(n120557), .B1(n120665), .B2(n120551), 
        .ZN(n7051) );
  OAI22_X1 U87631 ( .A1(n98894), .A2(n120557), .B1(n120668), .B2(n120551), 
        .ZN(n7052) );
  OAI22_X1 U87632 ( .A1(n98893), .A2(n120557), .B1(n120671), .B2(n120551), 
        .ZN(n7053) );
  OAI22_X1 U87633 ( .A1(n98892), .A2(n120557), .B1(n120674), .B2(n120551), 
        .ZN(n7054) );
  OAI22_X1 U87634 ( .A1(n98891), .A2(n120557), .B1(n120677), .B2(n120551), 
        .ZN(n7055) );
  OAI22_X1 U87635 ( .A1(n98890), .A2(n120557), .B1(n120680), .B2(n120551), 
        .ZN(n7056) );
  OAI22_X1 U87636 ( .A1(n98889), .A2(n120557), .B1(n120683), .B2(n120551), 
        .ZN(n7057) );
  OAI22_X1 U87637 ( .A1(n98888), .A2(n120557), .B1(n120686), .B2(n120551), 
        .ZN(n7058) );
  OAI22_X1 U87638 ( .A1(n98887), .A2(n120557), .B1(n120689), .B2(n120551), 
        .ZN(n7059) );
  OAI22_X1 U87639 ( .A1(n98886), .A2(n120557), .B1(n120692), .B2(n120551), 
        .ZN(n7060) );
  OAI22_X1 U87640 ( .A1(n98885), .A2(n120557), .B1(n120695), .B2(n120551), 
        .ZN(n7061) );
  OAI22_X1 U87641 ( .A1(n98884), .A2(n120558), .B1(n120698), .B2(n120551), 
        .ZN(n7062) );
  OAI22_X1 U87642 ( .A1(n98883), .A2(n120558), .B1(n120701), .B2(n120552), 
        .ZN(n7063) );
  OAI22_X1 U87643 ( .A1(n98882), .A2(n120558), .B1(n120704), .B2(n120552), 
        .ZN(n7064) );
  OAI22_X1 U87644 ( .A1(n98881), .A2(n120558), .B1(n120707), .B2(n120552), 
        .ZN(n7065) );
  OAI22_X1 U87645 ( .A1(n98880), .A2(n120558), .B1(n120710), .B2(n120552), 
        .ZN(n7066) );
  OAI22_X1 U87646 ( .A1(n98879), .A2(n120558), .B1(n120713), .B2(n120552), 
        .ZN(n7067) );
  OAI22_X1 U87647 ( .A1(n98878), .A2(n120558), .B1(n120716), .B2(n120552), 
        .ZN(n7068) );
  OAI22_X1 U87648 ( .A1(n98877), .A2(n120558), .B1(n120719), .B2(n120552), 
        .ZN(n7069) );
  OAI22_X1 U87649 ( .A1(n98876), .A2(n120558), .B1(n120722), .B2(n120552), 
        .ZN(n7070) );
  OAI22_X1 U87650 ( .A1(n98875), .A2(n120558), .B1(n120725), .B2(n120552), 
        .ZN(n7071) );
  OAI22_X1 U87651 ( .A1(n98874), .A2(n120558), .B1(n120728), .B2(n120552), 
        .ZN(n7072) );
  OAI22_X1 U87652 ( .A1(n98873), .A2(n120558), .B1(n120731), .B2(n120552), 
        .ZN(n7073) );
  OAI22_X1 U87653 ( .A1(n98872), .A2(n120559), .B1(n120734), .B2(n120552), 
        .ZN(n7074) );
  OAI22_X1 U87654 ( .A1(n98871), .A2(n120559), .B1(n120737), .B2(n120553), 
        .ZN(n7075) );
  OAI22_X1 U87655 ( .A1(n98870), .A2(n120559), .B1(n120740), .B2(n120553), 
        .ZN(n7076) );
  OAI22_X1 U87656 ( .A1(n98869), .A2(n120559), .B1(n120743), .B2(n120553), 
        .ZN(n7077) );
  OAI22_X1 U87657 ( .A1(n98868), .A2(n120559), .B1(n120746), .B2(n120553), 
        .ZN(n7078) );
  OAI22_X1 U87658 ( .A1(n98867), .A2(n120559), .B1(n120749), .B2(n120553), 
        .ZN(n7079) );
  OAI22_X1 U87659 ( .A1(n98866), .A2(n120559), .B1(n120752), .B2(n120553), 
        .ZN(n7080) );
  OAI22_X1 U87660 ( .A1(n98865), .A2(n120559), .B1(n120755), .B2(n120553), 
        .ZN(n7081) );
  OAI22_X1 U87661 ( .A1(n98864), .A2(n120559), .B1(n120758), .B2(n120553), 
        .ZN(n7082) );
  OAI22_X1 U87662 ( .A1(n98863), .A2(n120559), .B1(n120761), .B2(n120553), 
        .ZN(n7083) );
  OAI22_X1 U87663 ( .A1(n98862), .A2(n120559), .B1(n120764), .B2(n120553), 
        .ZN(n7084) );
  OAI22_X1 U87664 ( .A1(n98861), .A2(n120559), .B1(n120767), .B2(n120553), 
        .ZN(n7085) );
  OAI22_X1 U87665 ( .A1(n98860), .A2(n120560), .B1(n120770), .B2(n120553), 
        .ZN(n7086) );
  OAI22_X1 U87666 ( .A1(n98859), .A2(n120560), .B1(n120773), .B2(n120554), 
        .ZN(n7087) );
  OAI22_X1 U87667 ( .A1(n98858), .A2(n120560), .B1(n120776), .B2(n120554), 
        .ZN(n7088) );
  OAI22_X1 U87668 ( .A1(n98857), .A2(n120560), .B1(n120779), .B2(n120554), 
        .ZN(n7089) );
  OAI22_X1 U87669 ( .A1(n98856), .A2(n120560), .B1(n120782), .B2(n120554), 
        .ZN(n7090) );
  OAI22_X1 U87670 ( .A1(n98855), .A2(n120560), .B1(n120785), .B2(n120554), 
        .ZN(n7091) );
  OAI22_X1 U87671 ( .A1(n98854), .A2(n120560), .B1(n120788), .B2(n120554), 
        .ZN(n7092) );
  OAI22_X1 U87672 ( .A1(n98853), .A2(n120560), .B1(n120791), .B2(n120554), 
        .ZN(n7093) );
  OAI22_X1 U87673 ( .A1(n98852), .A2(n120560), .B1(n120794), .B2(n120554), 
        .ZN(n7094) );
  OAI22_X1 U87674 ( .A1(n98851), .A2(n120560), .B1(n120797), .B2(n120554), 
        .ZN(n7095) );
  OAI22_X1 U87675 ( .A1(n98850), .A2(n120560), .B1(n120800), .B2(n120554), 
        .ZN(n7096) );
  OAI22_X1 U87676 ( .A1(n98849), .A2(n120560), .B1(n120803), .B2(n120554), 
        .ZN(n7097) );
  OAI22_X1 U87677 ( .A1(n98848), .A2(n120561), .B1(n120806), .B2(n120554), 
        .ZN(n7098) );
  OAI22_X1 U87678 ( .A1(n98582), .A2(n120617), .B1(n120629), .B2(n120611), 
        .ZN(n7359) );
  OAI22_X1 U87679 ( .A1(n98581), .A2(n120617), .B1(n120632), .B2(n120611), 
        .ZN(n7360) );
  OAI22_X1 U87680 ( .A1(n98580), .A2(n120617), .B1(n120635), .B2(n120611), 
        .ZN(n7361) );
  OAI22_X1 U87681 ( .A1(n98579), .A2(n120617), .B1(n120638), .B2(n120611), 
        .ZN(n7362) );
  OAI22_X1 U87682 ( .A1(n98578), .A2(n120617), .B1(n120641), .B2(n120611), 
        .ZN(n7363) );
  OAI22_X1 U87683 ( .A1(n98577), .A2(n120617), .B1(n120644), .B2(n120611), 
        .ZN(n7364) );
  OAI22_X1 U87684 ( .A1(n98576), .A2(n120617), .B1(n120647), .B2(n120611), 
        .ZN(n7365) );
  OAI22_X1 U87685 ( .A1(n98575), .A2(n120617), .B1(n120650), .B2(n120611), 
        .ZN(n7366) );
  OAI22_X1 U87686 ( .A1(n98574), .A2(n120617), .B1(n120653), .B2(n120611), 
        .ZN(n7367) );
  OAI22_X1 U87687 ( .A1(n98573), .A2(n120617), .B1(n120656), .B2(n120611), 
        .ZN(n7368) );
  OAI22_X1 U87688 ( .A1(n98572), .A2(n120617), .B1(n120659), .B2(n120611), 
        .ZN(n7369) );
  OAI22_X1 U87689 ( .A1(n98571), .A2(n120618), .B1(n120662), .B2(n120611), 
        .ZN(n7370) );
  OAI22_X1 U87690 ( .A1(n98570), .A2(n120618), .B1(n120665), .B2(n120612), 
        .ZN(n7371) );
  OAI22_X1 U87691 ( .A1(n98569), .A2(n120618), .B1(n120668), .B2(n120612), 
        .ZN(n7372) );
  OAI22_X1 U87692 ( .A1(n98568), .A2(n120618), .B1(n120671), .B2(n120612), 
        .ZN(n7373) );
  OAI22_X1 U87693 ( .A1(n98567), .A2(n120618), .B1(n120674), .B2(n120612), 
        .ZN(n7374) );
  OAI22_X1 U87694 ( .A1(n98566), .A2(n120618), .B1(n120677), .B2(n120612), 
        .ZN(n7375) );
  OAI22_X1 U87695 ( .A1(n98565), .A2(n120618), .B1(n120680), .B2(n120612), 
        .ZN(n7376) );
  OAI22_X1 U87696 ( .A1(n98564), .A2(n120618), .B1(n120683), .B2(n120612), 
        .ZN(n7377) );
  OAI22_X1 U87697 ( .A1(n98563), .A2(n120618), .B1(n120686), .B2(n120612), 
        .ZN(n7378) );
  OAI22_X1 U87698 ( .A1(n98562), .A2(n120618), .B1(n120689), .B2(n120612), 
        .ZN(n7379) );
  OAI22_X1 U87699 ( .A1(n98561), .A2(n120618), .B1(n120692), .B2(n120612), 
        .ZN(n7380) );
  OAI22_X1 U87700 ( .A1(n98560), .A2(n120618), .B1(n120695), .B2(n120612), 
        .ZN(n7381) );
  OAI22_X1 U87701 ( .A1(n98559), .A2(n120619), .B1(n120698), .B2(n120612), 
        .ZN(n7382) );
  OAI22_X1 U87702 ( .A1(n98558), .A2(n120619), .B1(n120701), .B2(n120613), 
        .ZN(n7383) );
  OAI22_X1 U87703 ( .A1(n98557), .A2(n120619), .B1(n120704), .B2(n120613), 
        .ZN(n7384) );
  OAI22_X1 U87704 ( .A1(n98556), .A2(n120619), .B1(n120707), .B2(n120613), 
        .ZN(n7385) );
  OAI22_X1 U87705 ( .A1(n98555), .A2(n120619), .B1(n120710), .B2(n120613), 
        .ZN(n7386) );
  OAI22_X1 U87706 ( .A1(n98554), .A2(n120619), .B1(n120713), .B2(n120613), 
        .ZN(n7387) );
  OAI22_X1 U87707 ( .A1(n98553), .A2(n120619), .B1(n120716), .B2(n120613), 
        .ZN(n7388) );
  OAI22_X1 U87708 ( .A1(n98552), .A2(n120619), .B1(n120719), .B2(n120613), 
        .ZN(n7389) );
  OAI22_X1 U87709 ( .A1(n98551), .A2(n120619), .B1(n120722), .B2(n120613), 
        .ZN(n7390) );
  OAI22_X1 U87710 ( .A1(n98550), .A2(n120619), .B1(n120725), .B2(n120613), 
        .ZN(n7391) );
  OAI22_X1 U87711 ( .A1(n98549), .A2(n120619), .B1(n120728), .B2(n120613), 
        .ZN(n7392) );
  OAI22_X1 U87712 ( .A1(n98548), .A2(n120619), .B1(n120731), .B2(n120613), 
        .ZN(n7393) );
  OAI22_X1 U87713 ( .A1(n98547), .A2(n120620), .B1(n120734), .B2(n120613), 
        .ZN(n7394) );
  OAI22_X1 U87714 ( .A1(n98546), .A2(n120620), .B1(n120737), .B2(n120614), 
        .ZN(n7395) );
  OAI22_X1 U87715 ( .A1(n98545), .A2(n120620), .B1(n120740), .B2(n120614), 
        .ZN(n7396) );
  OAI22_X1 U87716 ( .A1(n98544), .A2(n120620), .B1(n120743), .B2(n120614), 
        .ZN(n7397) );
  OAI22_X1 U87717 ( .A1(n98543), .A2(n120620), .B1(n120746), .B2(n120614), 
        .ZN(n7398) );
  OAI22_X1 U87718 ( .A1(n98542), .A2(n120620), .B1(n120749), .B2(n120614), 
        .ZN(n7399) );
  OAI22_X1 U87719 ( .A1(n98541), .A2(n120620), .B1(n120752), .B2(n120614), 
        .ZN(n7400) );
  OAI22_X1 U87720 ( .A1(n98540), .A2(n120620), .B1(n120755), .B2(n120614), 
        .ZN(n7401) );
  OAI22_X1 U87721 ( .A1(n98539), .A2(n120620), .B1(n120758), .B2(n120614), 
        .ZN(n7402) );
  OAI22_X1 U87722 ( .A1(n98538), .A2(n120620), .B1(n120761), .B2(n120614), 
        .ZN(n7403) );
  OAI22_X1 U87723 ( .A1(n98537), .A2(n120620), .B1(n120764), .B2(n120614), 
        .ZN(n7404) );
  OAI22_X1 U87724 ( .A1(n98536), .A2(n120620), .B1(n120767), .B2(n120614), 
        .ZN(n7405) );
  OAI22_X1 U87725 ( .A1(n98535), .A2(n120621), .B1(n120770), .B2(n120614), 
        .ZN(n7406) );
  OAI22_X1 U87726 ( .A1(n98534), .A2(n120621), .B1(n120773), .B2(n120615), 
        .ZN(n7407) );
  OAI22_X1 U87727 ( .A1(n98533), .A2(n120621), .B1(n120776), .B2(n120615), 
        .ZN(n7408) );
  OAI22_X1 U87728 ( .A1(n98532), .A2(n120621), .B1(n120779), .B2(n120615), 
        .ZN(n7409) );
  OAI22_X1 U87729 ( .A1(n98531), .A2(n120621), .B1(n120782), .B2(n120615), 
        .ZN(n7410) );
  OAI22_X1 U87730 ( .A1(n98530), .A2(n120621), .B1(n120785), .B2(n120615), 
        .ZN(n7411) );
  OAI22_X1 U87731 ( .A1(n98529), .A2(n120621), .B1(n120788), .B2(n120615), 
        .ZN(n7412) );
  OAI22_X1 U87732 ( .A1(n98528), .A2(n120621), .B1(n120791), .B2(n120615), 
        .ZN(n7413) );
  OAI22_X1 U87733 ( .A1(n98527), .A2(n120621), .B1(n120794), .B2(n120615), 
        .ZN(n7414) );
  OAI22_X1 U87734 ( .A1(n98526), .A2(n120621), .B1(n120797), .B2(n120615), 
        .ZN(n7415) );
  OAI22_X1 U87735 ( .A1(n98525), .A2(n120621), .B1(n120800), .B2(n120615), 
        .ZN(n7416) );
  OAI22_X1 U87736 ( .A1(n98524), .A2(n120621), .B1(n120803), .B2(n120615), 
        .ZN(n7417) );
  OAI22_X1 U87737 ( .A1(n98523), .A2(n120622), .B1(n120806), .B2(n120615), 
        .ZN(n7418) );
  OAI22_X1 U87738 ( .A1(n98712), .A2(n120593), .B1(n120629), .B2(n120587), 
        .ZN(n7231) );
  OAI22_X1 U87739 ( .A1(n98711), .A2(n120593), .B1(n120632), .B2(n120587), 
        .ZN(n7232) );
  OAI22_X1 U87740 ( .A1(n98710), .A2(n120593), .B1(n120635), .B2(n120587), 
        .ZN(n7233) );
  OAI22_X1 U87741 ( .A1(n98709), .A2(n120593), .B1(n120638), .B2(n120587), 
        .ZN(n7234) );
  OAI22_X1 U87742 ( .A1(n98708), .A2(n120593), .B1(n120641), .B2(n120587), 
        .ZN(n7235) );
  OAI22_X1 U87743 ( .A1(n98707), .A2(n120593), .B1(n120644), .B2(n120587), 
        .ZN(n7236) );
  OAI22_X1 U87744 ( .A1(n98706), .A2(n120593), .B1(n120647), .B2(n120587), 
        .ZN(n7237) );
  OAI22_X1 U87745 ( .A1(n98705), .A2(n120593), .B1(n120650), .B2(n120587), 
        .ZN(n7238) );
  OAI22_X1 U87746 ( .A1(n98704), .A2(n120593), .B1(n120653), .B2(n120587), 
        .ZN(n7239) );
  OAI22_X1 U87747 ( .A1(n98703), .A2(n120593), .B1(n120656), .B2(n120587), 
        .ZN(n7240) );
  OAI22_X1 U87748 ( .A1(n98702), .A2(n120593), .B1(n120659), .B2(n120587), 
        .ZN(n7241) );
  OAI22_X1 U87749 ( .A1(n98701), .A2(n120594), .B1(n120662), .B2(n120587), 
        .ZN(n7242) );
  OAI22_X1 U87750 ( .A1(n98700), .A2(n120594), .B1(n120665), .B2(n120588), 
        .ZN(n7243) );
  OAI22_X1 U87751 ( .A1(n98699), .A2(n120594), .B1(n120668), .B2(n120588), 
        .ZN(n7244) );
  OAI22_X1 U87752 ( .A1(n98698), .A2(n120594), .B1(n120671), .B2(n120588), 
        .ZN(n7245) );
  OAI22_X1 U87753 ( .A1(n98697), .A2(n120594), .B1(n120674), .B2(n120588), 
        .ZN(n7246) );
  OAI22_X1 U87754 ( .A1(n98696), .A2(n120594), .B1(n120677), .B2(n120588), 
        .ZN(n7247) );
  OAI22_X1 U87755 ( .A1(n98695), .A2(n120594), .B1(n120680), .B2(n120588), 
        .ZN(n7248) );
  OAI22_X1 U87756 ( .A1(n98694), .A2(n120594), .B1(n120683), .B2(n120588), 
        .ZN(n7249) );
  OAI22_X1 U87757 ( .A1(n98693), .A2(n120594), .B1(n120686), .B2(n120588), 
        .ZN(n7250) );
  OAI22_X1 U87758 ( .A1(n98692), .A2(n120594), .B1(n120689), .B2(n120588), 
        .ZN(n7251) );
  OAI22_X1 U87759 ( .A1(n98691), .A2(n120594), .B1(n120692), .B2(n120588), 
        .ZN(n7252) );
  OAI22_X1 U87760 ( .A1(n98690), .A2(n120594), .B1(n120695), .B2(n120588), 
        .ZN(n7253) );
  OAI22_X1 U87761 ( .A1(n98689), .A2(n120595), .B1(n120698), .B2(n120588), 
        .ZN(n7254) );
  OAI22_X1 U87762 ( .A1(n98688), .A2(n120595), .B1(n120701), .B2(n120589), 
        .ZN(n7255) );
  OAI22_X1 U87763 ( .A1(n98687), .A2(n120595), .B1(n120704), .B2(n120589), 
        .ZN(n7256) );
  OAI22_X1 U87764 ( .A1(n98686), .A2(n120595), .B1(n120707), .B2(n120589), 
        .ZN(n7257) );
  OAI22_X1 U87765 ( .A1(n98685), .A2(n120595), .B1(n120710), .B2(n120589), 
        .ZN(n7258) );
  OAI22_X1 U87766 ( .A1(n98684), .A2(n120595), .B1(n120713), .B2(n120589), 
        .ZN(n7259) );
  OAI22_X1 U87767 ( .A1(n98683), .A2(n120595), .B1(n120716), .B2(n120589), 
        .ZN(n7260) );
  OAI22_X1 U87768 ( .A1(n98682), .A2(n120595), .B1(n120719), .B2(n120589), 
        .ZN(n7261) );
  OAI22_X1 U87769 ( .A1(n98681), .A2(n120595), .B1(n120722), .B2(n120589), 
        .ZN(n7262) );
  OAI22_X1 U87770 ( .A1(n98680), .A2(n120595), .B1(n120725), .B2(n120589), 
        .ZN(n7263) );
  OAI22_X1 U87771 ( .A1(n98679), .A2(n120595), .B1(n120728), .B2(n120589), 
        .ZN(n7264) );
  OAI22_X1 U87772 ( .A1(n98678), .A2(n120595), .B1(n120731), .B2(n120589), 
        .ZN(n7265) );
  OAI22_X1 U87773 ( .A1(n98677), .A2(n120596), .B1(n120734), .B2(n120589), 
        .ZN(n7266) );
  OAI22_X1 U87774 ( .A1(n98676), .A2(n120596), .B1(n120737), .B2(n120590), 
        .ZN(n7267) );
  OAI22_X1 U87775 ( .A1(n98675), .A2(n120596), .B1(n120740), .B2(n120590), 
        .ZN(n7268) );
  OAI22_X1 U87776 ( .A1(n98674), .A2(n120596), .B1(n120743), .B2(n120590), 
        .ZN(n7269) );
  OAI22_X1 U87777 ( .A1(n98673), .A2(n120596), .B1(n120746), .B2(n120590), 
        .ZN(n7270) );
  OAI22_X1 U87778 ( .A1(n98672), .A2(n120596), .B1(n120749), .B2(n120590), 
        .ZN(n7271) );
  OAI22_X1 U87779 ( .A1(n98671), .A2(n120596), .B1(n120752), .B2(n120590), 
        .ZN(n7272) );
  OAI22_X1 U87780 ( .A1(n98670), .A2(n120596), .B1(n120755), .B2(n120590), 
        .ZN(n7273) );
  OAI22_X1 U87781 ( .A1(n98669), .A2(n120596), .B1(n120758), .B2(n120590), 
        .ZN(n7274) );
  OAI22_X1 U87782 ( .A1(n98668), .A2(n120596), .B1(n120761), .B2(n120590), 
        .ZN(n7275) );
  OAI22_X1 U87783 ( .A1(n98667), .A2(n120596), .B1(n120764), .B2(n120590), 
        .ZN(n7276) );
  OAI22_X1 U87784 ( .A1(n98666), .A2(n120596), .B1(n120767), .B2(n120590), 
        .ZN(n7277) );
  OAI22_X1 U87785 ( .A1(n98665), .A2(n120597), .B1(n120770), .B2(n120590), 
        .ZN(n7278) );
  OAI22_X1 U87786 ( .A1(n98664), .A2(n120597), .B1(n120773), .B2(n120591), 
        .ZN(n7279) );
  OAI22_X1 U87787 ( .A1(n98663), .A2(n120597), .B1(n120776), .B2(n120591), 
        .ZN(n7280) );
  OAI22_X1 U87788 ( .A1(n98662), .A2(n120597), .B1(n120779), .B2(n120591), 
        .ZN(n7281) );
  OAI22_X1 U87789 ( .A1(n98661), .A2(n120597), .B1(n120782), .B2(n120591), 
        .ZN(n7282) );
  OAI22_X1 U87790 ( .A1(n98660), .A2(n120597), .B1(n120785), .B2(n120591), 
        .ZN(n7283) );
  OAI22_X1 U87791 ( .A1(n98659), .A2(n120597), .B1(n120788), .B2(n120591), 
        .ZN(n7284) );
  OAI22_X1 U87792 ( .A1(n98658), .A2(n120597), .B1(n120791), .B2(n120591), 
        .ZN(n7285) );
  OAI22_X1 U87793 ( .A1(n98657), .A2(n120597), .B1(n120794), .B2(n120591), 
        .ZN(n7286) );
  OAI22_X1 U87794 ( .A1(n98656), .A2(n120597), .B1(n120797), .B2(n120591), 
        .ZN(n7287) );
  OAI22_X1 U87795 ( .A1(n98655), .A2(n120597), .B1(n120800), .B2(n120591), 
        .ZN(n7288) );
  OAI22_X1 U87796 ( .A1(n98654), .A2(n120597), .B1(n120803), .B2(n120591), 
        .ZN(n7289) );
  OAI22_X1 U87797 ( .A1(n98653), .A2(n120598), .B1(n120806), .B2(n120591), 
        .ZN(n7290) );
  OAI22_X1 U87798 ( .A1(n98645), .A2(n120605), .B1(n120629), .B2(n120599), 
        .ZN(n7295) );
  OAI22_X1 U87799 ( .A1(n98644), .A2(n120605), .B1(n120632), .B2(n120599), 
        .ZN(n7296) );
  OAI22_X1 U87800 ( .A1(n98643), .A2(n120605), .B1(n120635), .B2(n120599), 
        .ZN(n7297) );
  OAI22_X1 U87801 ( .A1(n98642), .A2(n120605), .B1(n120638), .B2(n120599), 
        .ZN(n7298) );
  OAI22_X1 U87802 ( .A1(n98641), .A2(n120605), .B1(n120641), .B2(n120599), 
        .ZN(n7299) );
  OAI22_X1 U87803 ( .A1(n98640), .A2(n120605), .B1(n120644), .B2(n120599), 
        .ZN(n7300) );
  OAI22_X1 U87804 ( .A1(n98639), .A2(n120605), .B1(n120647), .B2(n120599), 
        .ZN(n7301) );
  OAI22_X1 U87805 ( .A1(n98638), .A2(n120605), .B1(n120650), .B2(n120599), 
        .ZN(n7302) );
  OAI22_X1 U87806 ( .A1(n98637), .A2(n120605), .B1(n120653), .B2(n120599), 
        .ZN(n7303) );
  OAI22_X1 U87807 ( .A1(n98636), .A2(n120605), .B1(n120656), .B2(n120599), 
        .ZN(n7304) );
  OAI22_X1 U87808 ( .A1(n98635), .A2(n120605), .B1(n120659), .B2(n120599), 
        .ZN(n7305) );
  OAI22_X1 U87809 ( .A1(n98634), .A2(n120606), .B1(n120662), .B2(n120599), 
        .ZN(n7306) );
  OAI22_X1 U87810 ( .A1(n98633), .A2(n120606), .B1(n120665), .B2(n120600), 
        .ZN(n7307) );
  OAI22_X1 U87811 ( .A1(n98632), .A2(n120606), .B1(n120668), .B2(n120600), 
        .ZN(n7308) );
  OAI22_X1 U87812 ( .A1(n98631), .A2(n120606), .B1(n120671), .B2(n120600), 
        .ZN(n7309) );
  OAI22_X1 U87813 ( .A1(n98630), .A2(n120606), .B1(n120674), .B2(n120600), 
        .ZN(n7310) );
  OAI22_X1 U87814 ( .A1(n98629), .A2(n120606), .B1(n120677), .B2(n120600), 
        .ZN(n7311) );
  OAI22_X1 U87815 ( .A1(n98628), .A2(n120606), .B1(n120680), .B2(n120600), 
        .ZN(n7312) );
  OAI22_X1 U87816 ( .A1(n98627), .A2(n120606), .B1(n120683), .B2(n120600), 
        .ZN(n7313) );
  OAI22_X1 U87817 ( .A1(n98626), .A2(n120606), .B1(n120686), .B2(n120600), 
        .ZN(n7314) );
  OAI22_X1 U87818 ( .A1(n98625), .A2(n120606), .B1(n120689), .B2(n120600), 
        .ZN(n7315) );
  OAI22_X1 U87819 ( .A1(n98624), .A2(n120606), .B1(n120692), .B2(n120600), 
        .ZN(n7316) );
  OAI22_X1 U87820 ( .A1(n98623), .A2(n120606), .B1(n120695), .B2(n120600), 
        .ZN(n7317) );
  OAI22_X1 U87821 ( .A1(n98622), .A2(n120607), .B1(n120698), .B2(n120600), 
        .ZN(n7318) );
  OAI22_X1 U87822 ( .A1(n98621), .A2(n120607), .B1(n120701), .B2(n120601), 
        .ZN(n7319) );
  OAI22_X1 U87823 ( .A1(n98620), .A2(n120607), .B1(n120704), .B2(n120601), 
        .ZN(n7320) );
  OAI22_X1 U87824 ( .A1(n98619), .A2(n120607), .B1(n120707), .B2(n120601), 
        .ZN(n7321) );
  OAI22_X1 U87825 ( .A1(n98618), .A2(n120607), .B1(n120710), .B2(n120601), 
        .ZN(n7322) );
  OAI22_X1 U87826 ( .A1(n98617), .A2(n120607), .B1(n120713), .B2(n120601), 
        .ZN(n7323) );
  OAI22_X1 U87827 ( .A1(n98616), .A2(n120607), .B1(n120716), .B2(n120601), 
        .ZN(n7324) );
  OAI22_X1 U87828 ( .A1(n98615), .A2(n120607), .B1(n120719), .B2(n120601), 
        .ZN(n7325) );
  OAI22_X1 U87829 ( .A1(n98614), .A2(n120607), .B1(n120722), .B2(n120601), 
        .ZN(n7326) );
  OAI22_X1 U87830 ( .A1(n98613), .A2(n120607), .B1(n120725), .B2(n120601), 
        .ZN(n7327) );
  OAI22_X1 U87831 ( .A1(n98612), .A2(n120607), .B1(n120728), .B2(n120601), 
        .ZN(n7328) );
  OAI22_X1 U87832 ( .A1(n98611), .A2(n120607), .B1(n120731), .B2(n120601), 
        .ZN(n7329) );
  OAI22_X1 U87833 ( .A1(n98610), .A2(n120608), .B1(n120734), .B2(n120601), 
        .ZN(n7330) );
  OAI22_X1 U87834 ( .A1(n98609), .A2(n120608), .B1(n120737), .B2(n120602), 
        .ZN(n7331) );
  OAI22_X1 U87835 ( .A1(n98608), .A2(n120608), .B1(n120740), .B2(n120602), 
        .ZN(n7332) );
  OAI22_X1 U87836 ( .A1(n98607), .A2(n120608), .B1(n120743), .B2(n120602), 
        .ZN(n7333) );
  OAI22_X1 U87837 ( .A1(n98606), .A2(n120608), .B1(n120746), .B2(n120602), 
        .ZN(n7334) );
  OAI22_X1 U87838 ( .A1(n98605), .A2(n120608), .B1(n120749), .B2(n120602), 
        .ZN(n7335) );
  OAI22_X1 U87839 ( .A1(n98604), .A2(n120608), .B1(n120752), .B2(n120602), 
        .ZN(n7336) );
  OAI22_X1 U87840 ( .A1(n98603), .A2(n120608), .B1(n120755), .B2(n120602), 
        .ZN(n7337) );
  OAI22_X1 U87841 ( .A1(n98602), .A2(n120608), .B1(n120758), .B2(n120602), 
        .ZN(n7338) );
  OAI22_X1 U87842 ( .A1(n98601), .A2(n120608), .B1(n120761), .B2(n120602), 
        .ZN(n7339) );
  OAI22_X1 U87843 ( .A1(n98600), .A2(n120608), .B1(n120764), .B2(n120602), 
        .ZN(n7340) );
  OAI22_X1 U87844 ( .A1(n98599), .A2(n120608), .B1(n120767), .B2(n120602), 
        .ZN(n7341) );
  OAI22_X1 U87845 ( .A1(n98598), .A2(n120609), .B1(n120770), .B2(n120602), 
        .ZN(n7342) );
  OAI22_X1 U87846 ( .A1(n98597), .A2(n120609), .B1(n120773), .B2(n120603), 
        .ZN(n7343) );
  OAI22_X1 U87847 ( .A1(n98596), .A2(n120609), .B1(n120776), .B2(n120603), 
        .ZN(n7344) );
  OAI22_X1 U87848 ( .A1(n98595), .A2(n120609), .B1(n120779), .B2(n120603), 
        .ZN(n7345) );
  OAI22_X1 U87849 ( .A1(n98594), .A2(n120609), .B1(n120782), .B2(n120603), 
        .ZN(n7346) );
  OAI22_X1 U87850 ( .A1(n98593), .A2(n120609), .B1(n120785), .B2(n120603), 
        .ZN(n7347) );
  OAI22_X1 U87851 ( .A1(n98592), .A2(n120609), .B1(n120788), .B2(n120603), 
        .ZN(n7348) );
  OAI22_X1 U87852 ( .A1(n98591), .A2(n120609), .B1(n120791), .B2(n120603), 
        .ZN(n7349) );
  OAI22_X1 U87853 ( .A1(n98590), .A2(n120609), .B1(n120794), .B2(n120603), 
        .ZN(n7350) );
  OAI22_X1 U87854 ( .A1(n98589), .A2(n120609), .B1(n120797), .B2(n120603), 
        .ZN(n7351) );
  OAI22_X1 U87855 ( .A1(n98588), .A2(n120609), .B1(n120800), .B2(n120603), 
        .ZN(n7352) );
  OAI22_X1 U87856 ( .A1(n98587), .A2(n120609), .B1(n120803), .B2(n120603), 
        .ZN(n7353) );
  OAI22_X1 U87857 ( .A1(n98586), .A2(n120610), .B1(n120806), .B2(n120603), 
        .ZN(n7354) );
  OAI22_X1 U87858 ( .A1(n99644), .A2(n120360), .B1(n120630), .B2(n120354), 
        .ZN(n6015) );
  OAI22_X1 U87859 ( .A1(n99643), .A2(n120360), .B1(n120633), .B2(n120354), 
        .ZN(n6016) );
  OAI22_X1 U87860 ( .A1(n99642), .A2(n120360), .B1(n120636), .B2(n120354), 
        .ZN(n6017) );
  OAI22_X1 U87861 ( .A1(n99641), .A2(n120360), .B1(n120639), .B2(n120354), 
        .ZN(n6018) );
  OAI22_X1 U87862 ( .A1(n99640), .A2(n120360), .B1(n120642), .B2(n120354), 
        .ZN(n6019) );
  OAI22_X1 U87863 ( .A1(n99639), .A2(n120360), .B1(n120645), .B2(n120354), 
        .ZN(n6020) );
  OAI22_X1 U87864 ( .A1(n99638), .A2(n120360), .B1(n120648), .B2(n120354), 
        .ZN(n6021) );
  OAI22_X1 U87865 ( .A1(n99637), .A2(n120360), .B1(n120651), .B2(n120354), 
        .ZN(n6022) );
  OAI22_X1 U87866 ( .A1(n99636), .A2(n120360), .B1(n120654), .B2(n120354), 
        .ZN(n6023) );
  OAI22_X1 U87867 ( .A1(n99635), .A2(n120360), .B1(n120657), .B2(n120354), 
        .ZN(n6024) );
  OAI22_X1 U87868 ( .A1(n99634), .A2(n120360), .B1(n120660), .B2(n120354), 
        .ZN(n6025) );
  OAI22_X1 U87869 ( .A1(n99633), .A2(n120361), .B1(n120663), .B2(n120354), 
        .ZN(n6026) );
  OAI22_X1 U87870 ( .A1(n99632), .A2(n120361), .B1(n120666), .B2(n120355), 
        .ZN(n6027) );
  OAI22_X1 U87871 ( .A1(n99631), .A2(n120361), .B1(n120669), .B2(n120355), 
        .ZN(n6028) );
  OAI22_X1 U87872 ( .A1(n99630), .A2(n120361), .B1(n120672), .B2(n120355), 
        .ZN(n6029) );
  OAI22_X1 U87873 ( .A1(n99629), .A2(n120361), .B1(n120675), .B2(n120355), 
        .ZN(n6030) );
  OAI22_X1 U87874 ( .A1(n99628), .A2(n120361), .B1(n120678), .B2(n120355), 
        .ZN(n6031) );
  OAI22_X1 U87875 ( .A1(n99627), .A2(n120361), .B1(n120681), .B2(n120355), 
        .ZN(n6032) );
  OAI22_X1 U87876 ( .A1(n99626), .A2(n120361), .B1(n120684), .B2(n120355), 
        .ZN(n6033) );
  OAI22_X1 U87877 ( .A1(n99625), .A2(n120361), .B1(n120687), .B2(n120355), 
        .ZN(n6034) );
  OAI22_X1 U87878 ( .A1(n99624), .A2(n120361), .B1(n120690), .B2(n120355), 
        .ZN(n6035) );
  OAI22_X1 U87879 ( .A1(n99623), .A2(n120361), .B1(n120693), .B2(n120355), 
        .ZN(n6036) );
  OAI22_X1 U87880 ( .A1(n99622), .A2(n120361), .B1(n120696), .B2(n120355), 
        .ZN(n6037) );
  OAI22_X1 U87881 ( .A1(n99621), .A2(n120362), .B1(n120699), .B2(n120355), 
        .ZN(n6038) );
  OAI22_X1 U87882 ( .A1(n99620), .A2(n120362), .B1(n120702), .B2(n120356), 
        .ZN(n6039) );
  OAI22_X1 U87883 ( .A1(n99619), .A2(n120362), .B1(n120705), .B2(n120356), 
        .ZN(n6040) );
  OAI22_X1 U87884 ( .A1(n99618), .A2(n120362), .B1(n120708), .B2(n120356), 
        .ZN(n6041) );
  OAI22_X1 U87885 ( .A1(n99617), .A2(n120362), .B1(n120711), .B2(n120356), 
        .ZN(n6042) );
  OAI22_X1 U87886 ( .A1(n99616), .A2(n120362), .B1(n120714), .B2(n120356), 
        .ZN(n6043) );
  OAI22_X1 U87887 ( .A1(n99615), .A2(n120362), .B1(n120717), .B2(n120356), 
        .ZN(n6044) );
  OAI22_X1 U87888 ( .A1(n99614), .A2(n120362), .B1(n120720), .B2(n120356), 
        .ZN(n6045) );
  OAI22_X1 U87889 ( .A1(n99613), .A2(n120362), .B1(n120723), .B2(n120356), 
        .ZN(n6046) );
  OAI22_X1 U87890 ( .A1(n99612), .A2(n120362), .B1(n120726), .B2(n120356), 
        .ZN(n6047) );
  OAI22_X1 U87891 ( .A1(n99611), .A2(n120362), .B1(n120729), .B2(n120356), 
        .ZN(n6048) );
  OAI22_X1 U87892 ( .A1(n99610), .A2(n120362), .B1(n120732), .B2(n120356), 
        .ZN(n6049) );
  OAI22_X1 U87893 ( .A1(n99609), .A2(n120363), .B1(n120735), .B2(n120356), 
        .ZN(n6050) );
  OAI22_X1 U87894 ( .A1(n99608), .A2(n120363), .B1(n120738), .B2(n120357), 
        .ZN(n6051) );
  OAI22_X1 U87895 ( .A1(n99607), .A2(n120363), .B1(n120741), .B2(n120357), 
        .ZN(n6052) );
  OAI22_X1 U87896 ( .A1(n99606), .A2(n120363), .B1(n120744), .B2(n120357), 
        .ZN(n6053) );
  OAI22_X1 U87897 ( .A1(n99605), .A2(n120363), .B1(n120747), .B2(n120357), 
        .ZN(n6054) );
  OAI22_X1 U87898 ( .A1(n99604), .A2(n120363), .B1(n120750), .B2(n120357), 
        .ZN(n6055) );
  OAI22_X1 U87899 ( .A1(n99603), .A2(n120363), .B1(n120753), .B2(n120357), 
        .ZN(n6056) );
  OAI22_X1 U87900 ( .A1(n99602), .A2(n120363), .B1(n120756), .B2(n120357), 
        .ZN(n6057) );
  OAI22_X1 U87901 ( .A1(n99601), .A2(n120363), .B1(n120759), .B2(n120357), 
        .ZN(n6058) );
  OAI22_X1 U87902 ( .A1(n99600), .A2(n120363), .B1(n120762), .B2(n120357), 
        .ZN(n6059) );
  OAI22_X1 U87903 ( .A1(n99599), .A2(n120363), .B1(n120765), .B2(n120357), 
        .ZN(n6060) );
  OAI22_X1 U87904 ( .A1(n99598), .A2(n120363), .B1(n120768), .B2(n120357), 
        .ZN(n6061) );
  OAI22_X1 U87905 ( .A1(n99597), .A2(n120364), .B1(n120771), .B2(n120357), 
        .ZN(n6062) );
  OAI22_X1 U87906 ( .A1(n99596), .A2(n120364), .B1(n120774), .B2(n120358), 
        .ZN(n6063) );
  OAI22_X1 U87907 ( .A1(n99595), .A2(n120364), .B1(n120777), .B2(n120358), 
        .ZN(n6064) );
  OAI22_X1 U87908 ( .A1(n99594), .A2(n120364), .B1(n120780), .B2(n120358), 
        .ZN(n6065) );
  OAI22_X1 U87909 ( .A1(n99593), .A2(n120364), .B1(n120783), .B2(n120358), 
        .ZN(n6066) );
  OAI22_X1 U87910 ( .A1(n99592), .A2(n120364), .B1(n120786), .B2(n120358), 
        .ZN(n6067) );
  OAI22_X1 U87911 ( .A1(n99591), .A2(n120364), .B1(n120789), .B2(n120358), 
        .ZN(n6068) );
  OAI22_X1 U87912 ( .A1(n99590), .A2(n120364), .B1(n120792), .B2(n120358), 
        .ZN(n6069) );
  OAI22_X1 U87913 ( .A1(n99589), .A2(n120364), .B1(n120795), .B2(n120358), 
        .ZN(n6070) );
  OAI22_X1 U87914 ( .A1(n99588), .A2(n120364), .B1(n120798), .B2(n120358), 
        .ZN(n6071) );
  OAI22_X1 U87915 ( .A1(n99587), .A2(n120364), .B1(n120801), .B2(n120358), 
        .ZN(n6072) );
  OAI22_X1 U87916 ( .A1(n99586), .A2(n120364), .B1(n120804), .B2(n120358), 
        .ZN(n6073) );
  OAI22_X1 U87917 ( .A1(n99585), .A2(n120365), .B1(n120807), .B2(n120358), 
        .ZN(n6074) );
  OAI22_X1 U87918 ( .A1(n120337), .A2(n114370), .B1(n120630), .B2(n120329), 
        .ZN(n5887) );
  OAI22_X1 U87919 ( .A1(n120337), .A2(n114369), .B1(n120633), .B2(n120329), 
        .ZN(n5888) );
  OAI22_X1 U87920 ( .A1(n120337), .A2(n114368), .B1(n120636), .B2(n120329), 
        .ZN(n5889) );
  OAI22_X1 U87921 ( .A1(n120337), .A2(n114367), .B1(n120639), .B2(n120329), 
        .ZN(n5890) );
  OAI22_X1 U87922 ( .A1(n120337), .A2(n114366), .B1(n120642), .B2(n120329), 
        .ZN(n5891) );
  OAI22_X1 U87923 ( .A1(n120337), .A2(n114365), .B1(n120645), .B2(n120329), 
        .ZN(n5892) );
  OAI22_X1 U87924 ( .A1(n120337), .A2(n114364), .B1(n120648), .B2(n120329), 
        .ZN(n5893) );
  OAI22_X1 U87925 ( .A1(n120337), .A2(n114363), .B1(n120651), .B2(n120329), 
        .ZN(n5894) );
  OAI22_X1 U87926 ( .A1(n120337), .A2(n114362), .B1(n120654), .B2(n120329), 
        .ZN(n5895) );
  OAI22_X1 U87927 ( .A1(n120337), .A2(n114361), .B1(n120657), .B2(n120329), 
        .ZN(n5896) );
  OAI22_X1 U87928 ( .A1(n120337), .A2(n114360), .B1(n120660), .B2(n120329), 
        .ZN(n5897) );
  OAI22_X1 U87929 ( .A1(n120337), .A2(n114359), .B1(n120663), .B2(n120329), 
        .ZN(n5898) );
  OAI22_X1 U87930 ( .A1(n120338), .A2(n114358), .B1(n120666), .B2(n120330), 
        .ZN(n5899) );
  OAI22_X1 U87931 ( .A1(n120338), .A2(n114357), .B1(n120669), .B2(n120330), 
        .ZN(n5900) );
  OAI22_X1 U87932 ( .A1(n120338), .A2(n114356), .B1(n120672), .B2(n120330), 
        .ZN(n5901) );
  OAI22_X1 U87933 ( .A1(n120338), .A2(n114355), .B1(n120675), .B2(n120330), 
        .ZN(n5902) );
  OAI22_X1 U87934 ( .A1(n120338), .A2(n114354), .B1(n120678), .B2(n120330), 
        .ZN(n5903) );
  OAI22_X1 U87935 ( .A1(n120338), .A2(n114353), .B1(n120681), .B2(n120330), 
        .ZN(n5904) );
  OAI22_X1 U87936 ( .A1(n120338), .A2(n114352), .B1(n120684), .B2(n120330), 
        .ZN(n5905) );
  OAI22_X1 U87937 ( .A1(n120338), .A2(n114351), .B1(n120687), .B2(n120330), 
        .ZN(n5906) );
  OAI22_X1 U87938 ( .A1(n120338), .A2(n114350), .B1(n120690), .B2(n120330), 
        .ZN(n5907) );
  OAI22_X1 U87939 ( .A1(n120338), .A2(n114349), .B1(n120693), .B2(n120330), 
        .ZN(n5908) );
  OAI22_X1 U87940 ( .A1(n120338), .A2(n114348), .B1(n120696), .B2(n120330), 
        .ZN(n5909) );
  OAI22_X1 U87941 ( .A1(n120338), .A2(n114347), .B1(n120699), .B2(n120330), 
        .ZN(n5910) );
  OAI22_X1 U87942 ( .A1(n120338), .A2(n114346), .B1(n120702), .B2(n120331), 
        .ZN(n5911) );
  OAI22_X1 U87943 ( .A1(n120339), .A2(n114345), .B1(n120705), .B2(n120331), 
        .ZN(n5912) );
  OAI22_X1 U87944 ( .A1(n120339), .A2(n114344), .B1(n120708), .B2(n120331), 
        .ZN(n5913) );
  OAI22_X1 U87945 ( .A1(n120339), .A2(n114343), .B1(n120711), .B2(n120331), 
        .ZN(n5914) );
  OAI22_X1 U87946 ( .A1(n120339), .A2(n114342), .B1(n120714), .B2(n120331), 
        .ZN(n5915) );
  OAI22_X1 U87947 ( .A1(n120339), .A2(n114341), .B1(n120717), .B2(n120331), 
        .ZN(n5916) );
  OAI22_X1 U87948 ( .A1(n120339), .A2(n114340), .B1(n120720), .B2(n120331), 
        .ZN(n5917) );
  OAI22_X1 U87949 ( .A1(n120339), .A2(n114339), .B1(n120723), .B2(n120331), 
        .ZN(n5918) );
  OAI22_X1 U87950 ( .A1(n120339), .A2(n114338), .B1(n120726), .B2(n120331), 
        .ZN(n5919) );
  OAI22_X1 U87951 ( .A1(n120339), .A2(n114337), .B1(n120729), .B2(n120331), 
        .ZN(n5920) );
  OAI22_X1 U87952 ( .A1(n120339), .A2(n114336), .B1(n120732), .B2(n120331), 
        .ZN(n5921) );
  OAI22_X1 U87953 ( .A1(n120339), .A2(n114335), .B1(n120735), .B2(n120331), 
        .ZN(n5922) );
  OAI22_X1 U87954 ( .A1(n120339), .A2(n114334), .B1(n120738), .B2(n120332), 
        .ZN(n5923) );
  OAI22_X1 U87955 ( .A1(n120339), .A2(n114333), .B1(n120741), .B2(n120332), 
        .ZN(n5924) );
  OAI22_X1 U87956 ( .A1(n120340), .A2(n114332), .B1(n120744), .B2(n120332), 
        .ZN(n5925) );
  OAI22_X1 U87957 ( .A1(n120340), .A2(n114331), .B1(n120747), .B2(n120332), 
        .ZN(n5926) );
  OAI22_X1 U87958 ( .A1(n120340), .A2(n114330), .B1(n120750), .B2(n120332), 
        .ZN(n5927) );
  OAI22_X1 U87959 ( .A1(n120340), .A2(n114329), .B1(n120753), .B2(n120332), 
        .ZN(n5928) );
  OAI22_X1 U87960 ( .A1(n120340), .A2(n114328), .B1(n120756), .B2(n120332), 
        .ZN(n5929) );
  OAI22_X1 U87961 ( .A1(n120340), .A2(n114327), .B1(n120759), .B2(n120332), 
        .ZN(n5930) );
  OAI22_X1 U87962 ( .A1(n120340), .A2(n114326), .B1(n120762), .B2(n120332), 
        .ZN(n5931) );
  OAI22_X1 U87963 ( .A1(n120340), .A2(n114325), .B1(n120765), .B2(n120332), 
        .ZN(n5932) );
  OAI22_X1 U87964 ( .A1(n120340), .A2(n114324), .B1(n120768), .B2(n120332), 
        .ZN(n5933) );
  OAI22_X1 U87965 ( .A1(n120340), .A2(n114323), .B1(n120771), .B2(n120332), 
        .ZN(n5934) );
  OAI22_X1 U87966 ( .A1(n120340), .A2(n114322), .B1(n120774), .B2(n120333), 
        .ZN(n5935) );
  OAI22_X1 U87967 ( .A1(n120340), .A2(n114321), .B1(n120777), .B2(n120333), 
        .ZN(n5936) );
  OAI22_X1 U87968 ( .A1(n120340), .A2(n114320), .B1(n120780), .B2(n120333), 
        .ZN(n5937) );
  OAI22_X1 U87969 ( .A1(n120341), .A2(n114319), .B1(n120783), .B2(n120333), 
        .ZN(n5938) );
  OAI22_X1 U87970 ( .A1(n120341), .A2(n114318), .B1(n120786), .B2(n120333), 
        .ZN(n5939) );
  OAI22_X1 U87971 ( .A1(n120341), .A2(n114317), .B1(n120789), .B2(n120333), 
        .ZN(n5940) );
  OAI22_X1 U87972 ( .A1(n120341), .A2(n114316), .B1(n120792), .B2(n120333), 
        .ZN(n5941) );
  OAI22_X1 U87973 ( .A1(n120341), .A2(n114315), .B1(n120795), .B2(n120333), 
        .ZN(n5942) );
  OAI22_X1 U87974 ( .A1(n120341), .A2(n114314), .B1(n120798), .B2(n120333), 
        .ZN(n5943) );
  OAI22_X1 U87975 ( .A1(n120341), .A2(n114313), .B1(n120801), .B2(n120333), 
        .ZN(n5944) );
  OAI22_X1 U87976 ( .A1(n120341), .A2(n114312), .B1(n120804), .B2(n120333), 
        .ZN(n5945) );
  OAI22_X1 U87977 ( .A1(n120341), .A2(n114311), .B1(n120807), .B2(n120333), 
        .ZN(n5946) );
  OAI22_X1 U87978 ( .A1(n99510), .A2(n120397), .B1(n120630), .B2(n120391), 
        .ZN(n6207) );
  OAI22_X1 U87979 ( .A1(n99509), .A2(n120397), .B1(n120633), .B2(n120391), 
        .ZN(n6208) );
  OAI22_X1 U87980 ( .A1(n99508), .A2(n120397), .B1(n120636), .B2(n120391), 
        .ZN(n6209) );
  OAI22_X1 U87981 ( .A1(n99507), .A2(n120397), .B1(n120639), .B2(n120391), 
        .ZN(n6210) );
  OAI22_X1 U87982 ( .A1(n99506), .A2(n120397), .B1(n120642), .B2(n120391), 
        .ZN(n6211) );
  OAI22_X1 U87983 ( .A1(n99505), .A2(n120397), .B1(n120645), .B2(n120391), 
        .ZN(n6212) );
  OAI22_X1 U87984 ( .A1(n99504), .A2(n120397), .B1(n120648), .B2(n120391), 
        .ZN(n6213) );
  OAI22_X1 U87985 ( .A1(n99503), .A2(n120397), .B1(n120651), .B2(n120391), 
        .ZN(n6214) );
  OAI22_X1 U87986 ( .A1(n99502), .A2(n120397), .B1(n120654), .B2(n120391), 
        .ZN(n6215) );
  OAI22_X1 U87987 ( .A1(n99501), .A2(n120397), .B1(n120657), .B2(n120391), 
        .ZN(n6216) );
  OAI22_X1 U87988 ( .A1(n99500), .A2(n120397), .B1(n120660), .B2(n120391), 
        .ZN(n6217) );
  OAI22_X1 U87989 ( .A1(n99499), .A2(n120398), .B1(n120663), .B2(n120391), 
        .ZN(n6218) );
  OAI22_X1 U87990 ( .A1(n99498), .A2(n120398), .B1(n120666), .B2(n120392), 
        .ZN(n6219) );
  OAI22_X1 U87991 ( .A1(n99497), .A2(n120398), .B1(n120669), .B2(n120392), 
        .ZN(n6220) );
  OAI22_X1 U87992 ( .A1(n99496), .A2(n120398), .B1(n120672), .B2(n120392), 
        .ZN(n6221) );
  OAI22_X1 U87993 ( .A1(n99495), .A2(n120398), .B1(n120675), .B2(n120392), 
        .ZN(n6222) );
  OAI22_X1 U87994 ( .A1(n99494), .A2(n120398), .B1(n120678), .B2(n120392), 
        .ZN(n6223) );
  OAI22_X1 U87995 ( .A1(n99493), .A2(n120398), .B1(n120681), .B2(n120392), 
        .ZN(n6224) );
  OAI22_X1 U87996 ( .A1(n99492), .A2(n120398), .B1(n120684), .B2(n120392), 
        .ZN(n6225) );
  OAI22_X1 U87997 ( .A1(n99491), .A2(n120398), .B1(n120687), .B2(n120392), 
        .ZN(n6226) );
  OAI22_X1 U87998 ( .A1(n99490), .A2(n120398), .B1(n120690), .B2(n120392), 
        .ZN(n6227) );
  OAI22_X1 U87999 ( .A1(n99489), .A2(n120398), .B1(n120693), .B2(n120392), 
        .ZN(n6228) );
  OAI22_X1 U88000 ( .A1(n99488), .A2(n120398), .B1(n120696), .B2(n120392), 
        .ZN(n6229) );
  OAI22_X1 U88001 ( .A1(n99487), .A2(n120399), .B1(n120699), .B2(n120392), 
        .ZN(n6230) );
  OAI22_X1 U88002 ( .A1(n99486), .A2(n120399), .B1(n120702), .B2(n120393), 
        .ZN(n6231) );
  OAI22_X1 U88003 ( .A1(n99485), .A2(n120399), .B1(n120705), .B2(n120393), 
        .ZN(n6232) );
  OAI22_X1 U88004 ( .A1(n99484), .A2(n120399), .B1(n120708), .B2(n120393), 
        .ZN(n6233) );
  OAI22_X1 U88005 ( .A1(n99483), .A2(n120399), .B1(n120711), .B2(n120393), 
        .ZN(n6234) );
  OAI22_X1 U88006 ( .A1(n99482), .A2(n120399), .B1(n120714), .B2(n120393), 
        .ZN(n6235) );
  OAI22_X1 U88007 ( .A1(n99481), .A2(n120399), .B1(n120717), .B2(n120393), 
        .ZN(n6236) );
  OAI22_X1 U88008 ( .A1(n99480), .A2(n120399), .B1(n120720), .B2(n120393), 
        .ZN(n6237) );
  OAI22_X1 U88009 ( .A1(n99479), .A2(n120399), .B1(n120723), .B2(n120393), 
        .ZN(n6238) );
  OAI22_X1 U88010 ( .A1(n99478), .A2(n120399), .B1(n120726), .B2(n120393), 
        .ZN(n6239) );
  OAI22_X1 U88011 ( .A1(n99477), .A2(n120399), .B1(n120729), .B2(n120393), 
        .ZN(n6240) );
  OAI22_X1 U88012 ( .A1(n99476), .A2(n120399), .B1(n120732), .B2(n120393), 
        .ZN(n6241) );
  OAI22_X1 U88013 ( .A1(n99475), .A2(n120400), .B1(n120735), .B2(n120393), 
        .ZN(n6242) );
  OAI22_X1 U88014 ( .A1(n99474), .A2(n120400), .B1(n120738), .B2(n120394), 
        .ZN(n6243) );
  OAI22_X1 U88015 ( .A1(n99473), .A2(n120400), .B1(n120741), .B2(n120394), 
        .ZN(n6244) );
  OAI22_X1 U88016 ( .A1(n99472), .A2(n120400), .B1(n120744), .B2(n120394), 
        .ZN(n6245) );
  OAI22_X1 U88017 ( .A1(n99471), .A2(n120400), .B1(n120747), .B2(n120394), 
        .ZN(n6246) );
  OAI22_X1 U88018 ( .A1(n99470), .A2(n120400), .B1(n120750), .B2(n120394), 
        .ZN(n6247) );
  OAI22_X1 U88019 ( .A1(n99469), .A2(n120400), .B1(n120753), .B2(n120394), 
        .ZN(n6248) );
  OAI22_X1 U88020 ( .A1(n99468), .A2(n120400), .B1(n120756), .B2(n120394), 
        .ZN(n6249) );
  OAI22_X1 U88021 ( .A1(n99467), .A2(n120400), .B1(n120759), .B2(n120394), 
        .ZN(n6250) );
  OAI22_X1 U88022 ( .A1(n99466), .A2(n120400), .B1(n120762), .B2(n120394), 
        .ZN(n6251) );
  OAI22_X1 U88023 ( .A1(n99465), .A2(n120400), .B1(n120765), .B2(n120394), 
        .ZN(n6252) );
  OAI22_X1 U88024 ( .A1(n99464), .A2(n120400), .B1(n120768), .B2(n120394), 
        .ZN(n6253) );
  OAI22_X1 U88025 ( .A1(n99463), .A2(n120401), .B1(n120771), .B2(n120394), 
        .ZN(n6254) );
  OAI22_X1 U88026 ( .A1(n99462), .A2(n120401), .B1(n120774), .B2(n120395), 
        .ZN(n6255) );
  OAI22_X1 U88027 ( .A1(n99461), .A2(n120401), .B1(n120777), .B2(n120395), 
        .ZN(n6256) );
  OAI22_X1 U88028 ( .A1(n99460), .A2(n120401), .B1(n120780), .B2(n120395), 
        .ZN(n6257) );
  OAI22_X1 U88029 ( .A1(n99459), .A2(n120401), .B1(n120783), .B2(n120395), 
        .ZN(n6258) );
  OAI22_X1 U88030 ( .A1(n99458), .A2(n120401), .B1(n120786), .B2(n120395), 
        .ZN(n6259) );
  OAI22_X1 U88031 ( .A1(n99457), .A2(n120401), .B1(n120789), .B2(n120395), 
        .ZN(n6260) );
  OAI22_X1 U88032 ( .A1(n99456), .A2(n120401), .B1(n120792), .B2(n120395), 
        .ZN(n6261) );
  OAI22_X1 U88033 ( .A1(n99455), .A2(n120401), .B1(n120795), .B2(n120395), 
        .ZN(n6262) );
  OAI22_X1 U88034 ( .A1(n99454), .A2(n120401), .B1(n120798), .B2(n120395), 
        .ZN(n6263) );
  OAI22_X1 U88035 ( .A1(n99453), .A2(n120401), .B1(n120801), .B2(n120395), 
        .ZN(n6264) );
  OAI22_X1 U88036 ( .A1(n99452), .A2(n120401), .B1(n120804), .B2(n120395), 
        .ZN(n6265) );
  OAI22_X1 U88037 ( .A1(n99451), .A2(n120402), .B1(n120807), .B2(n120395), 
        .ZN(n6266) );
  OAI22_X1 U88038 ( .A1(n90557), .A2(n120388), .B1(n120687), .B2(n120380), 
        .ZN(n6162) );
  OAI22_X1 U88039 ( .A1(n90556), .A2(n120388), .B1(n120690), .B2(n120380), 
        .ZN(n6163) );
  OAI22_X1 U88040 ( .A1(n90555), .A2(n120388), .B1(n120693), .B2(n120380), 
        .ZN(n6164) );
  OAI22_X1 U88041 ( .A1(n90554), .A2(n120388), .B1(n120696), .B2(n120380), 
        .ZN(n6165) );
  OAI22_X1 U88042 ( .A1(n90553), .A2(n120388), .B1(n120699), .B2(n120380), 
        .ZN(n6166) );
  OAI22_X1 U88043 ( .A1(n90552), .A2(n120388), .B1(n120702), .B2(n120381), 
        .ZN(n6167) );
  OAI22_X1 U88044 ( .A1(n90551), .A2(n120388), .B1(n120705), .B2(n120381), 
        .ZN(n6168) );
  OAI22_X1 U88045 ( .A1(n90550), .A2(n120388), .B1(n120708), .B2(n120381), 
        .ZN(n6169) );
  OAI22_X1 U88046 ( .A1(n90549), .A2(n120388), .B1(n120711), .B2(n120381), 
        .ZN(n6170) );
  OAI22_X1 U88047 ( .A1(n90548), .A2(n120388), .B1(n120714), .B2(n120381), 
        .ZN(n6171) );
  OAI22_X1 U88048 ( .A1(n90547), .A2(n120387), .B1(n120717), .B2(n120381), 
        .ZN(n6172) );
  OAI22_X1 U88049 ( .A1(n90546), .A2(n120387), .B1(n120720), .B2(n120381), 
        .ZN(n6173) );
  OAI22_X1 U88050 ( .A1(n90545), .A2(n120387), .B1(n120723), .B2(n120381), 
        .ZN(n6174) );
  OAI22_X1 U88051 ( .A1(n90544), .A2(n120387), .B1(n120726), .B2(n120381), 
        .ZN(n6175) );
  OAI22_X1 U88052 ( .A1(n90543), .A2(n120387), .B1(n120729), .B2(n120381), 
        .ZN(n6176) );
  OAI22_X1 U88053 ( .A1(n90542), .A2(n120387), .B1(n120732), .B2(n120381), 
        .ZN(n6177) );
  OAI22_X1 U88054 ( .A1(n90541), .A2(n120387), .B1(n120735), .B2(n120381), 
        .ZN(n6178) );
  OAI22_X1 U88055 ( .A1(n90540), .A2(n120387), .B1(n120738), .B2(n120382), 
        .ZN(n6179) );
  OAI22_X1 U88056 ( .A1(n90539), .A2(n120387), .B1(n120741), .B2(n120382), 
        .ZN(n6180) );
  OAI22_X1 U88057 ( .A1(n90538), .A2(n120387), .B1(n120744), .B2(n120382), 
        .ZN(n6181) );
  OAI22_X1 U88058 ( .A1(n90537), .A2(n120387), .B1(n120747), .B2(n120382), 
        .ZN(n6182) );
  OAI22_X1 U88059 ( .A1(n90536), .A2(n120386), .B1(n120750), .B2(n120382), 
        .ZN(n6183) );
  OAI22_X1 U88060 ( .A1(n90535), .A2(n120386), .B1(n120753), .B2(n120382), 
        .ZN(n6184) );
  OAI22_X1 U88061 ( .A1(n90534), .A2(n120386), .B1(n120756), .B2(n120382), 
        .ZN(n6185) );
  OAI22_X1 U88062 ( .A1(n90533), .A2(n120386), .B1(n120759), .B2(n120382), 
        .ZN(n6186) );
  OAI22_X1 U88063 ( .A1(n90532), .A2(n120386), .B1(n120762), .B2(n120382), 
        .ZN(n6187) );
  OAI22_X1 U88064 ( .A1(n90531), .A2(n120386), .B1(n120765), .B2(n120382), 
        .ZN(n6188) );
  OAI22_X1 U88065 ( .A1(n90530), .A2(n120386), .B1(n120768), .B2(n120382), 
        .ZN(n6189) );
  OAI22_X1 U88066 ( .A1(n90529), .A2(n120386), .B1(n120771), .B2(n120382), 
        .ZN(n6190) );
  OAI22_X1 U88067 ( .A1(n90528), .A2(n120386), .B1(n120774), .B2(n120383), 
        .ZN(n6191) );
  OAI22_X1 U88068 ( .A1(n90527), .A2(n120386), .B1(n120777), .B2(n120383), 
        .ZN(n6192) );
  OAI22_X1 U88069 ( .A1(n90526), .A2(n120386), .B1(n120780), .B2(n120383), 
        .ZN(n6193) );
  OAI22_X1 U88070 ( .A1(n90525), .A2(n120386), .B1(n120783), .B2(n120383), 
        .ZN(n6194) );
  OAI22_X1 U88071 ( .A1(n90524), .A2(n120385), .B1(n120786), .B2(n120383), 
        .ZN(n6195) );
  OAI22_X1 U88072 ( .A1(n90523), .A2(n120385), .B1(n120789), .B2(n120383), 
        .ZN(n6196) );
  OAI22_X1 U88073 ( .A1(n90522), .A2(n120385), .B1(n120792), .B2(n120383), 
        .ZN(n6197) );
  OAI22_X1 U88074 ( .A1(n90521), .A2(n120385), .B1(n120795), .B2(n120383), 
        .ZN(n6198) );
  OAI22_X1 U88075 ( .A1(n90520), .A2(n120385), .B1(n120798), .B2(n120383), 
        .ZN(n6199) );
  OAI22_X1 U88076 ( .A1(n90519), .A2(n120385), .B1(n120801), .B2(n120383), 
        .ZN(n6200) );
  OAI22_X1 U88077 ( .A1(n90518), .A2(n120385), .B1(n120804), .B2(n120383), 
        .ZN(n6201) );
  OAI22_X1 U88078 ( .A1(n90517), .A2(n120385), .B1(n120807), .B2(n120383), 
        .ZN(n6202) );
  OAI22_X1 U88079 ( .A1(n90370), .A2(n120434), .B1(n120630), .B2(n120428), 
        .ZN(n6399) );
  OAI22_X1 U88080 ( .A1(n90369), .A2(n120434), .B1(n120633), .B2(n120428), 
        .ZN(n6400) );
  OAI22_X1 U88081 ( .A1(n90368), .A2(n120434), .B1(n120636), .B2(n120428), 
        .ZN(n6401) );
  OAI22_X1 U88082 ( .A1(n90367), .A2(n120434), .B1(n120639), .B2(n120428), 
        .ZN(n6402) );
  OAI22_X1 U88083 ( .A1(n90366), .A2(n120434), .B1(n120642), .B2(n120428), 
        .ZN(n6403) );
  OAI22_X1 U88084 ( .A1(n90365), .A2(n120434), .B1(n120645), .B2(n120428), 
        .ZN(n6404) );
  OAI22_X1 U88085 ( .A1(n90364), .A2(n120434), .B1(n120648), .B2(n120428), 
        .ZN(n6405) );
  OAI22_X1 U88086 ( .A1(n90363), .A2(n120434), .B1(n120651), .B2(n120428), 
        .ZN(n6406) );
  OAI22_X1 U88087 ( .A1(n90362), .A2(n120434), .B1(n120654), .B2(n120428), 
        .ZN(n6407) );
  OAI22_X1 U88088 ( .A1(n90361), .A2(n120434), .B1(n120657), .B2(n120428), 
        .ZN(n6408) );
  OAI22_X1 U88089 ( .A1(n90360), .A2(n120434), .B1(n120660), .B2(n120428), 
        .ZN(n6409) );
  OAI22_X1 U88090 ( .A1(n90359), .A2(n120435), .B1(n120663), .B2(n120428), 
        .ZN(n6410) );
  OAI22_X1 U88091 ( .A1(n90358), .A2(n120435), .B1(n120666), .B2(n120429), 
        .ZN(n6411) );
  OAI22_X1 U88092 ( .A1(n90357), .A2(n120435), .B1(n120669), .B2(n120429), 
        .ZN(n6412) );
  OAI22_X1 U88093 ( .A1(n90356), .A2(n120435), .B1(n120672), .B2(n120429), 
        .ZN(n6413) );
  OAI22_X1 U88094 ( .A1(n90355), .A2(n120435), .B1(n120675), .B2(n120429), 
        .ZN(n6414) );
  OAI22_X1 U88095 ( .A1(n90354), .A2(n120435), .B1(n120678), .B2(n120429), 
        .ZN(n6415) );
  OAI22_X1 U88096 ( .A1(n90353), .A2(n120435), .B1(n120681), .B2(n120429), 
        .ZN(n6416) );
  OAI22_X1 U88097 ( .A1(n90352), .A2(n120435), .B1(n120684), .B2(n120429), 
        .ZN(n6417) );
  OAI22_X1 U88098 ( .A1(n90351), .A2(n120435), .B1(n120687), .B2(n120429), 
        .ZN(n6418) );
  OAI22_X1 U88099 ( .A1(n90350), .A2(n120435), .B1(n120690), .B2(n120429), 
        .ZN(n6419) );
  OAI22_X1 U88100 ( .A1(n90349), .A2(n120435), .B1(n120693), .B2(n120429), 
        .ZN(n6420) );
  OAI22_X1 U88101 ( .A1(n90348), .A2(n120435), .B1(n120696), .B2(n120429), 
        .ZN(n6421) );
  OAI22_X1 U88102 ( .A1(n90347), .A2(n120436), .B1(n120699), .B2(n120429), 
        .ZN(n6422) );
  OAI22_X1 U88103 ( .A1(n90346), .A2(n120436), .B1(n120702), .B2(n120430), 
        .ZN(n6423) );
  OAI22_X1 U88104 ( .A1(n90345), .A2(n120436), .B1(n120705), .B2(n120430), 
        .ZN(n6424) );
  OAI22_X1 U88105 ( .A1(n90344), .A2(n120436), .B1(n120708), .B2(n120430), 
        .ZN(n6425) );
  OAI22_X1 U88106 ( .A1(n90343), .A2(n120436), .B1(n120711), .B2(n120430), 
        .ZN(n6426) );
  OAI22_X1 U88107 ( .A1(n90342), .A2(n120436), .B1(n120714), .B2(n120430), 
        .ZN(n6427) );
  OAI22_X1 U88108 ( .A1(n90341), .A2(n120436), .B1(n120717), .B2(n120430), 
        .ZN(n6428) );
  OAI22_X1 U88109 ( .A1(n90340), .A2(n120436), .B1(n120720), .B2(n120430), 
        .ZN(n6429) );
  OAI22_X1 U88110 ( .A1(n90339), .A2(n120436), .B1(n120723), .B2(n120430), 
        .ZN(n6430) );
  OAI22_X1 U88111 ( .A1(n90338), .A2(n120436), .B1(n120726), .B2(n120430), 
        .ZN(n6431) );
  OAI22_X1 U88112 ( .A1(n90337), .A2(n120436), .B1(n120729), .B2(n120430), 
        .ZN(n6432) );
  OAI22_X1 U88113 ( .A1(n90336), .A2(n120436), .B1(n120732), .B2(n120430), 
        .ZN(n6433) );
  OAI22_X1 U88114 ( .A1(n90335), .A2(n120437), .B1(n120735), .B2(n120430), 
        .ZN(n6434) );
  OAI22_X1 U88115 ( .A1(n90334), .A2(n120437), .B1(n120738), .B2(n120431), 
        .ZN(n6435) );
  OAI22_X1 U88116 ( .A1(n90333), .A2(n120437), .B1(n120741), .B2(n120431), 
        .ZN(n6436) );
  OAI22_X1 U88117 ( .A1(n90332), .A2(n120437), .B1(n120744), .B2(n120431), 
        .ZN(n6437) );
  OAI22_X1 U88118 ( .A1(n90331), .A2(n120437), .B1(n120747), .B2(n120431), 
        .ZN(n6438) );
  OAI22_X1 U88119 ( .A1(n90330), .A2(n120437), .B1(n120750), .B2(n120431), 
        .ZN(n6439) );
  OAI22_X1 U88120 ( .A1(n90329), .A2(n120437), .B1(n120753), .B2(n120431), 
        .ZN(n6440) );
  OAI22_X1 U88121 ( .A1(n90328), .A2(n120437), .B1(n120756), .B2(n120431), 
        .ZN(n6441) );
  OAI22_X1 U88122 ( .A1(n90327), .A2(n120437), .B1(n120759), .B2(n120431), 
        .ZN(n6442) );
  OAI22_X1 U88123 ( .A1(n90326), .A2(n120437), .B1(n120762), .B2(n120431), 
        .ZN(n6443) );
  OAI22_X1 U88124 ( .A1(n90325), .A2(n120437), .B1(n120765), .B2(n120431), 
        .ZN(n6444) );
  OAI22_X1 U88125 ( .A1(n90324), .A2(n120437), .B1(n120768), .B2(n120431), 
        .ZN(n6445) );
  OAI22_X1 U88126 ( .A1(n90323), .A2(n120438), .B1(n120771), .B2(n120431), 
        .ZN(n6446) );
  OAI22_X1 U88127 ( .A1(n90322), .A2(n120438), .B1(n120774), .B2(n120432), 
        .ZN(n6447) );
  OAI22_X1 U88128 ( .A1(n90321), .A2(n120438), .B1(n120777), .B2(n120432), 
        .ZN(n6448) );
  OAI22_X1 U88129 ( .A1(n90320), .A2(n120438), .B1(n120780), .B2(n120432), 
        .ZN(n6449) );
  OAI22_X1 U88130 ( .A1(n90319), .A2(n120438), .B1(n120783), .B2(n120432), 
        .ZN(n6450) );
  OAI22_X1 U88131 ( .A1(n90318), .A2(n120438), .B1(n120786), .B2(n120432), 
        .ZN(n6451) );
  OAI22_X1 U88132 ( .A1(n90317), .A2(n120438), .B1(n120789), .B2(n120432), 
        .ZN(n6452) );
  OAI22_X1 U88133 ( .A1(n90316), .A2(n120438), .B1(n120792), .B2(n120432), 
        .ZN(n6453) );
  OAI22_X1 U88134 ( .A1(n90315), .A2(n120438), .B1(n120795), .B2(n120432), 
        .ZN(n6454) );
  OAI22_X1 U88135 ( .A1(n90314), .A2(n120438), .B1(n120798), .B2(n120432), 
        .ZN(n6455) );
  OAI22_X1 U88136 ( .A1(n90313), .A2(n120438), .B1(n120801), .B2(n120432), 
        .ZN(n6456) );
  OAI22_X1 U88137 ( .A1(n90312), .A2(n120438), .B1(n120804), .B2(n120432), 
        .ZN(n6457) );
  OAI22_X1 U88138 ( .A1(n90311), .A2(n120439), .B1(n120807), .B2(n120432), 
        .ZN(n6458) );
  OAI22_X1 U88139 ( .A1(n90437), .A2(n120422), .B1(n120630), .B2(n120416), 
        .ZN(n6335) );
  OAI22_X1 U88140 ( .A1(n90436), .A2(n120422), .B1(n120633), .B2(n120416), 
        .ZN(n6336) );
  OAI22_X1 U88141 ( .A1(n90435), .A2(n120422), .B1(n120636), .B2(n120416), 
        .ZN(n6337) );
  OAI22_X1 U88142 ( .A1(n90434), .A2(n120422), .B1(n120639), .B2(n120416), 
        .ZN(n6338) );
  OAI22_X1 U88143 ( .A1(n90433), .A2(n120422), .B1(n120642), .B2(n120416), 
        .ZN(n6339) );
  OAI22_X1 U88144 ( .A1(n90432), .A2(n120422), .B1(n120645), .B2(n120416), 
        .ZN(n6340) );
  OAI22_X1 U88145 ( .A1(n90431), .A2(n120422), .B1(n120648), .B2(n120416), 
        .ZN(n6341) );
  OAI22_X1 U88146 ( .A1(n90430), .A2(n120422), .B1(n120651), .B2(n120416), 
        .ZN(n6342) );
  OAI22_X1 U88147 ( .A1(n90429), .A2(n120422), .B1(n120654), .B2(n120416), 
        .ZN(n6343) );
  OAI22_X1 U88148 ( .A1(n90428), .A2(n120422), .B1(n120657), .B2(n120416), 
        .ZN(n6344) );
  OAI22_X1 U88149 ( .A1(n90427), .A2(n120422), .B1(n120660), .B2(n120416), 
        .ZN(n6345) );
  OAI22_X1 U88150 ( .A1(n90426), .A2(n120423), .B1(n120663), .B2(n120416), 
        .ZN(n6346) );
  OAI22_X1 U88151 ( .A1(n90425), .A2(n120423), .B1(n120666), .B2(n120417), 
        .ZN(n6347) );
  OAI22_X1 U88152 ( .A1(n90424), .A2(n120423), .B1(n120669), .B2(n120417), 
        .ZN(n6348) );
  OAI22_X1 U88153 ( .A1(n90423), .A2(n120423), .B1(n120672), .B2(n120417), 
        .ZN(n6349) );
  OAI22_X1 U88154 ( .A1(n90422), .A2(n120423), .B1(n120675), .B2(n120417), 
        .ZN(n6350) );
  OAI22_X1 U88155 ( .A1(n90421), .A2(n120423), .B1(n120678), .B2(n120417), 
        .ZN(n6351) );
  OAI22_X1 U88156 ( .A1(n90420), .A2(n120423), .B1(n120681), .B2(n120417), 
        .ZN(n6352) );
  OAI22_X1 U88157 ( .A1(n90419), .A2(n120423), .B1(n120684), .B2(n120417), 
        .ZN(n6353) );
  OAI22_X1 U88158 ( .A1(n90418), .A2(n120423), .B1(n120687), .B2(n120417), 
        .ZN(n6354) );
  OAI22_X1 U88159 ( .A1(n90417), .A2(n120423), .B1(n120690), .B2(n120417), 
        .ZN(n6355) );
  OAI22_X1 U88160 ( .A1(n90416), .A2(n120423), .B1(n120693), .B2(n120417), 
        .ZN(n6356) );
  OAI22_X1 U88161 ( .A1(n90415), .A2(n120423), .B1(n120696), .B2(n120417), 
        .ZN(n6357) );
  OAI22_X1 U88162 ( .A1(n90414), .A2(n120424), .B1(n120699), .B2(n120417), 
        .ZN(n6358) );
  OAI22_X1 U88163 ( .A1(n90413), .A2(n120424), .B1(n120702), .B2(n120418), 
        .ZN(n6359) );
  OAI22_X1 U88164 ( .A1(n90412), .A2(n120424), .B1(n120705), .B2(n120418), 
        .ZN(n6360) );
  OAI22_X1 U88165 ( .A1(n90411), .A2(n120424), .B1(n120708), .B2(n120418), 
        .ZN(n6361) );
  OAI22_X1 U88166 ( .A1(n90410), .A2(n120424), .B1(n120711), .B2(n120418), 
        .ZN(n6362) );
  OAI22_X1 U88167 ( .A1(n90409), .A2(n120424), .B1(n120714), .B2(n120418), 
        .ZN(n6363) );
  OAI22_X1 U88168 ( .A1(n90408), .A2(n120424), .B1(n120717), .B2(n120418), 
        .ZN(n6364) );
  OAI22_X1 U88169 ( .A1(n90407), .A2(n120424), .B1(n120720), .B2(n120418), 
        .ZN(n6365) );
  OAI22_X1 U88170 ( .A1(n90406), .A2(n120424), .B1(n120723), .B2(n120418), 
        .ZN(n6366) );
  OAI22_X1 U88171 ( .A1(n90405), .A2(n120424), .B1(n120726), .B2(n120418), 
        .ZN(n6367) );
  OAI22_X1 U88172 ( .A1(n90404), .A2(n120424), .B1(n120729), .B2(n120418), 
        .ZN(n6368) );
  OAI22_X1 U88173 ( .A1(n90403), .A2(n120424), .B1(n120732), .B2(n120418), 
        .ZN(n6369) );
  OAI22_X1 U88174 ( .A1(n90402), .A2(n120425), .B1(n120735), .B2(n120418), 
        .ZN(n6370) );
  OAI22_X1 U88175 ( .A1(n90401), .A2(n120425), .B1(n120738), .B2(n120419), 
        .ZN(n6371) );
  OAI22_X1 U88176 ( .A1(n90400), .A2(n120425), .B1(n120741), .B2(n120419), 
        .ZN(n6372) );
  OAI22_X1 U88177 ( .A1(n90399), .A2(n120425), .B1(n120744), .B2(n120419), 
        .ZN(n6373) );
  OAI22_X1 U88178 ( .A1(n90398), .A2(n120425), .B1(n120747), .B2(n120419), 
        .ZN(n6374) );
  OAI22_X1 U88179 ( .A1(n90397), .A2(n120425), .B1(n120750), .B2(n120419), 
        .ZN(n6375) );
  OAI22_X1 U88180 ( .A1(n90396), .A2(n120425), .B1(n120753), .B2(n120419), 
        .ZN(n6376) );
  OAI22_X1 U88181 ( .A1(n90395), .A2(n120425), .B1(n120756), .B2(n120419), 
        .ZN(n6377) );
  OAI22_X1 U88182 ( .A1(n90394), .A2(n120425), .B1(n120759), .B2(n120419), 
        .ZN(n6378) );
  OAI22_X1 U88183 ( .A1(n90393), .A2(n120425), .B1(n120762), .B2(n120419), 
        .ZN(n6379) );
  OAI22_X1 U88184 ( .A1(n90392), .A2(n120425), .B1(n120765), .B2(n120419), 
        .ZN(n6380) );
  OAI22_X1 U88185 ( .A1(n90391), .A2(n120425), .B1(n120768), .B2(n120419), 
        .ZN(n6381) );
  OAI22_X1 U88186 ( .A1(n90390), .A2(n120426), .B1(n120771), .B2(n120419), 
        .ZN(n6382) );
  OAI22_X1 U88187 ( .A1(n90389), .A2(n120426), .B1(n120774), .B2(n120420), 
        .ZN(n6383) );
  OAI22_X1 U88188 ( .A1(n90388), .A2(n120426), .B1(n120777), .B2(n120420), 
        .ZN(n6384) );
  OAI22_X1 U88189 ( .A1(n90387), .A2(n120426), .B1(n120780), .B2(n120420), 
        .ZN(n6385) );
  OAI22_X1 U88190 ( .A1(n90386), .A2(n120426), .B1(n120783), .B2(n120420), 
        .ZN(n6386) );
  OAI22_X1 U88191 ( .A1(n90385), .A2(n120426), .B1(n120786), .B2(n120420), 
        .ZN(n6387) );
  OAI22_X1 U88192 ( .A1(n90384), .A2(n120426), .B1(n120789), .B2(n120420), 
        .ZN(n6388) );
  OAI22_X1 U88193 ( .A1(n90383), .A2(n120426), .B1(n120792), .B2(n120420), 
        .ZN(n6389) );
  OAI22_X1 U88194 ( .A1(n90382), .A2(n120426), .B1(n120795), .B2(n120420), 
        .ZN(n6390) );
  OAI22_X1 U88195 ( .A1(n90381), .A2(n120426), .B1(n120798), .B2(n120420), 
        .ZN(n6391) );
  OAI22_X1 U88196 ( .A1(n90380), .A2(n120426), .B1(n120801), .B2(n120420), 
        .ZN(n6392) );
  OAI22_X1 U88197 ( .A1(n90379), .A2(n120426), .B1(n120804), .B2(n120420), 
        .ZN(n6393) );
  OAI22_X1 U88198 ( .A1(n90378), .A2(n120427), .B1(n120807), .B2(n120420), 
        .ZN(n6394) );
  OAI22_X1 U88199 ( .A1(n90775), .A2(n120348), .B1(n120630), .B2(n120342), 
        .ZN(n5951) );
  OAI22_X1 U88200 ( .A1(n90774), .A2(n120348), .B1(n120633), .B2(n120342), 
        .ZN(n5952) );
  OAI22_X1 U88201 ( .A1(n90773), .A2(n120348), .B1(n120636), .B2(n120342), 
        .ZN(n5953) );
  OAI22_X1 U88202 ( .A1(n90772), .A2(n120348), .B1(n120639), .B2(n120342), 
        .ZN(n5954) );
  OAI22_X1 U88203 ( .A1(n90771), .A2(n120348), .B1(n120642), .B2(n120342), 
        .ZN(n5955) );
  OAI22_X1 U88204 ( .A1(n90770), .A2(n120348), .B1(n120645), .B2(n120342), 
        .ZN(n5956) );
  OAI22_X1 U88205 ( .A1(n90769), .A2(n120348), .B1(n120648), .B2(n120342), 
        .ZN(n5957) );
  OAI22_X1 U88206 ( .A1(n90768), .A2(n120348), .B1(n120651), .B2(n120342), 
        .ZN(n5958) );
  OAI22_X1 U88207 ( .A1(n90767), .A2(n120348), .B1(n120654), .B2(n120342), 
        .ZN(n5959) );
  OAI22_X1 U88208 ( .A1(n90766), .A2(n120348), .B1(n120657), .B2(n120342), 
        .ZN(n5960) );
  OAI22_X1 U88209 ( .A1(n90765), .A2(n120348), .B1(n120660), .B2(n120342), 
        .ZN(n5961) );
  OAI22_X1 U88210 ( .A1(n90764), .A2(n120349), .B1(n120663), .B2(n120342), 
        .ZN(n5962) );
  OAI22_X1 U88211 ( .A1(n90763), .A2(n120349), .B1(n120666), .B2(n120343), 
        .ZN(n5963) );
  OAI22_X1 U88212 ( .A1(n90762), .A2(n120349), .B1(n120669), .B2(n120343), 
        .ZN(n5964) );
  OAI22_X1 U88213 ( .A1(n90761), .A2(n120349), .B1(n120672), .B2(n120343), 
        .ZN(n5965) );
  OAI22_X1 U88214 ( .A1(n90760), .A2(n120349), .B1(n120675), .B2(n120343), 
        .ZN(n5966) );
  OAI22_X1 U88215 ( .A1(n90759), .A2(n120349), .B1(n120678), .B2(n120343), 
        .ZN(n5967) );
  OAI22_X1 U88216 ( .A1(n90758), .A2(n120349), .B1(n120681), .B2(n120343), 
        .ZN(n5968) );
  OAI22_X1 U88217 ( .A1(n90757), .A2(n120349), .B1(n120684), .B2(n120343), 
        .ZN(n5969) );
  OAI22_X1 U88218 ( .A1(n90756), .A2(n120349), .B1(n120687), .B2(n120343), 
        .ZN(n5970) );
  OAI22_X1 U88219 ( .A1(n90755), .A2(n120349), .B1(n120690), .B2(n120343), 
        .ZN(n5971) );
  OAI22_X1 U88220 ( .A1(n90754), .A2(n120349), .B1(n120693), .B2(n120343), 
        .ZN(n5972) );
  OAI22_X1 U88221 ( .A1(n90753), .A2(n120349), .B1(n120696), .B2(n120343), 
        .ZN(n5973) );
  OAI22_X1 U88222 ( .A1(n90752), .A2(n120350), .B1(n120699), .B2(n120343), 
        .ZN(n5974) );
  OAI22_X1 U88223 ( .A1(n90751), .A2(n120350), .B1(n120702), .B2(n120344), 
        .ZN(n5975) );
  OAI22_X1 U88224 ( .A1(n90750), .A2(n120350), .B1(n120705), .B2(n120344), 
        .ZN(n5976) );
  OAI22_X1 U88225 ( .A1(n90749), .A2(n120350), .B1(n120708), .B2(n120344), 
        .ZN(n5977) );
  OAI22_X1 U88226 ( .A1(n90748), .A2(n120350), .B1(n120711), .B2(n120344), 
        .ZN(n5978) );
  OAI22_X1 U88227 ( .A1(n90747), .A2(n120350), .B1(n120714), .B2(n120344), 
        .ZN(n5979) );
  OAI22_X1 U88228 ( .A1(n90746), .A2(n120350), .B1(n120717), .B2(n120344), 
        .ZN(n5980) );
  OAI22_X1 U88229 ( .A1(n90745), .A2(n120350), .B1(n120720), .B2(n120344), 
        .ZN(n5981) );
  OAI22_X1 U88230 ( .A1(n90744), .A2(n120350), .B1(n120723), .B2(n120344), 
        .ZN(n5982) );
  OAI22_X1 U88231 ( .A1(n90743), .A2(n120350), .B1(n120726), .B2(n120344), 
        .ZN(n5983) );
  OAI22_X1 U88232 ( .A1(n90742), .A2(n120350), .B1(n120729), .B2(n120344), 
        .ZN(n5984) );
  OAI22_X1 U88233 ( .A1(n90741), .A2(n120350), .B1(n120732), .B2(n120344), 
        .ZN(n5985) );
  OAI22_X1 U88234 ( .A1(n90740), .A2(n120351), .B1(n120735), .B2(n120344), 
        .ZN(n5986) );
  OAI22_X1 U88235 ( .A1(n90739), .A2(n120351), .B1(n120738), .B2(n120345), 
        .ZN(n5987) );
  OAI22_X1 U88236 ( .A1(n90738), .A2(n120351), .B1(n120741), .B2(n120345), 
        .ZN(n5988) );
  OAI22_X1 U88237 ( .A1(n90737), .A2(n120351), .B1(n120744), .B2(n120345), 
        .ZN(n5989) );
  OAI22_X1 U88238 ( .A1(n90736), .A2(n120351), .B1(n120747), .B2(n120345), 
        .ZN(n5990) );
  OAI22_X1 U88239 ( .A1(n90735), .A2(n120351), .B1(n120750), .B2(n120345), 
        .ZN(n5991) );
  OAI22_X1 U88240 ( .A1(n90734), .A2(n120351), .B1(n120753), .B2(n120345), 
        .ZN(n5992) );
  OAI22_X1 U88241 ( .A1(n90733), .A2(n120351), .B1(n120756), .B2(n120345), 
        .ZN(n5993) );
  OAI22_X1 U88242 ( .A1(n90732), .A2(n120351), .B1(n120759), .B2(n120345), 
        .ZN(n5994) );
  OAI22_X1 U88243 ( .A1(n90731), .A2(n120351), .B1(n120762), .B2(n120345), 
        .ZN(n5995) );
  OAI22_X1 U88244 ( .A1(n90730), .A2(n120351), .B1(n120765), .B2(n120345), 
        .ZN(n5996) );
  OAI22_X1 U88245 ( .A1(n90729), .A2(n120351), .B1(n120768), .B2(n120345), 
        .ZN(n5997) );
  OAI22_X1 U88246 ( .A1(n90728), .A2(n120352), .B1(n120771), .B2(n120345), 
        .ZN(n5998) );
  OAI22_X1 U88247 ( .A1(n90727), .A2(n120352), .B1(n120774), .B2(n120346), 
        .ZN(n5999) );
  OAI22_X1 U88248 ( .A1(n90726), .A2(n120352), .B1(n120777), .B2(n120346), 
        .ZN(n6000) );
  OAI22_X1 U88249 ( .A1(n90725), .A2(n120352), .B1(n120780), .B2(n120346), 
        .ZN(n6001) );
  OAI22_X1 U88250 ( .A1(n90724), .A2(n120352), .B1(n120783), .B2(n120346), 
        .ZN(n6002) );
  OAI22_X1 U88251 ( .A1(n90723), .A2(n120352), .B1(n120786), .B2(n120346), 
        .ZN(n6003) );
  OAI22_X1 U88252 ( .A1(n90722), .A2(n120352), .B1(n120789), .B2(n120346), 
        .ZN(n6004) );
  OAI22_X1 U88253 ( .A1(n90721), .A2(n120352), .B1(n120792), .B2(n120346), 
        .ZN(n6005) );
  OAI22_X1 U88254 ( .A1(n90720), .A2(n120352), .B1(n120795), .B2(n120346), 
        .ZN(n6006) );
  OAI22_X1 U88255 ( .A1(n90719), .A2(n120352), .B1(n120798), .B2(n120346), 
        .ZN(n6007) );
  OAI22_X1 U88256 ( .A1(n90718), .A2(n120352), .B1(n120801), .B2(n120346), 
        .ZN(n6008) );
  OAI22_X1 U88257 ( .A1(n90717), .A2(n120352), .B1(n120804), .B2(n120346), 
        .ZN(n6009) );
  OAI22_X1 U88258 ( .A1(n90716), .A2(n120353), .B1(n120807), .B2(n120346), 
        .ZN(n6010) );
  OAI22_X1 U88259 ( .A1(n90095), .A2(n120531), .B1(n120629), .B2(n120525), 
        .ZN(n6911) );
  OAI22_X1 U88260 ( .A1(n90094), .A2(n120531), .B1(n120632), .B2(n120525), 
        .ZN(n6912) );
  OAI22_X1 U88261 ( .A1(n90093), .A2(n120531), .B1(n120635), .B2(n120525), 
        .ZN(n6913) );
  OAI22_X1 U88262 ( .A1(n90092), .A2(n120531), .B1(n120638), .B2(n120525), 
        .ZN(n6914) );
  OAI22_X1 U88263 ( .A1(n90091), .A2(n120531), .B1(n120641), .B2(n120525), 
        .ZN(n6915) );
  OAI22_X1 U88264 ( .A1(n90090), .A2(n120531), .B1(n120644), .B2(n120525), 
        .ZN(n6916) );
  OAI22_X1 U88265 ( .A1(n90089), .A2(n120531), .B1(n120647), .B2(n120525), 
        .ZN(n6917) );
  OAI22_X1 U88266 ( .A1(n90088), .A2(n120531), .B1(n120650), .B2(n120525), 
        .ZN(n6918) );
  OAI22_X1 U88267 ( .A1(n90087), .A2(n120531), .B1(n120653), .B2(n120525), 
        .ZN(n6919) );
  OAI22_X1 U88268 ( .A1(n90086), .A2(n120531), .B1(n120656), .B2(n120525), 
        .ZN(n6920) );
  OAI22_X1 U88269 ( .A1(n90085), .A2(n120531), .B1(n120659), .B2(n120525), 
        .ZN(n6921) );
  OAI22_X1 U88270 ( .A1(n90084), .A2(n120532), .B1(n120662), .B2(n120525), 
        .ZN(n6922) );
  OAI22_X1 U88271 ( .A1(n90083), .A2(n120532), .B1(n120665), .B2(n120526), 
        .ZN(n6923) );
  OAI22_X1 U88272 ( .A1(n90082), .A2(n120532), .B1(n120668), .B2(n120526), 
        .ZN(n6924) );
  OAI22_X1 U88273 ( .A1(n90081), .A2(n120532), .B1(n120671), .B2(n120526), 
        .ZN(n6925) );
  OAI22_X1 U88274 ( .A1(n90080), .A2(n120532), .B1(n120674), .B2(n120526), 
        .ZN(n6926) );
  OAI22_X1 U88275 ( .A1(n90079), .A2(n120532), .B1(n120677), .B2(n120526), 
        .ZN(n6927) );
  OAI22_X1 U88276 ( .A1(n90078), .A2(n120532), .B1(n120680), .B2(n120526), 
        .ZN(n6928) );
  OAI22_X1 U88277 ( .A1(n90077), .A2(n120532), .B1(n120683), .B2(n120526), 
        .ZN(n6929) );
  OAI22_X1 U88278 ( .A1(n90076), .A2(n120532), .B1(n120686), .B2(n120526), 
        .ZN(n6930) );
  OAI22_X1 U88279 ( .A1(n90075), .A2(n120532), .B1(n120689), .B2(n120526), 
        .ZN(n6931) );
  OAI22_X1 U88280 ( .A1(n90074), .A2(n120532), .B1(n120692), .B2(n120526), 
        .ZN(n6932) );
  OAI22_X1 U88281 ( .A1(n90073), .A2(n120532), .B1(n120695), .B2(n120526), 
        .ZN(n6933) );
  OAI22_X1 U88282 ( .A1(n90072), .A2(n120533), .B1(n120698), .B2(n120526), 
        .ZN(n6934) );
  OAI22_X1 U88283 ( .A1(n90071), .A2(n120533), .B1(n120701), .B2(n120527), 
        .ZN(n6935) );
  OAI22_X1 U88284 ( .A1(n90070), .A2(n120533), .B1(n120704), .B2(n120527), 
        .ZN(n6936) );
  OAI22_X1 U88285 ( .A1(n90069), .A2(n120533), .B1(n120707), .B2(n120527), 
        .ZN(n6937) );
  OAI22_X1 U88286 ( .A1(n90068), .A2(n120533), .B1(n120710), .B2(n120527), 
        .ZN(n6938) );
  OAI22_X1 U88287 ( .A1(n90067), .A2(n120533), .B1(n120713), .B2(n120527), 
        .ZN(n6939) );
  OAI22_X1 U88288 ( .A1(n90066), .A2(n120533), .B1(n120716), .B2(n120527), 
        .ZN(n6940) );
  OAI22_X1 U88289 ( .A1(n90065), .A2(n120533), .B1(n120719), .B2(n120527), 
        .ZN(n6941) );
  OAI22_X1 U88290 ( .A1(n90064), .A2(n120533), .B1(n120722), .B2(n120527), 
        .ZN(n6942) );
  OAI22_X1 U88291 ( .A1(n90063), .A2(n120533), .B1(n120725), .B2(n120527), 
        .ZN(n6943) );
  OAI22_X1 U88292 ( .A1(n90062), .A2(n120533), .B1(n120728), .B2(n120527), 
        .ZN(n6944) );
  OAI22_X1 U88293 ( .A1(n90061), .A2(n120533), .B1(n120731), .B2(n120527), 
        .ZN(n6945) );
  OAI22_X1 U88294 ( .A1(n90060), .A2(n120534), .B1(n120734), .B2(n120527), 
        .ZN(n6946) );
  OAI22_X1 U88295 ( .A1(n90059), .A2(n120534), .B1(n120737), .B2(n120528), 
        .ZN(n6947) );
  OAI22_X1 U88296 ( .A1(n90058), .A2(n120534), .B1(n120740), .B2(n120528), 
        .ZN(n6948) );
  OAI22_X1 U88297 ( .A1(n90057), .A2(n120534), .B1(n120743), .B2(n120528), 
        .ZN(n6949) );
  OAI22_X1 U88298 ( .A1(n90056), .A2(n120534), .B1(n120746), .B2(n120528), 
        .ZN(n6950) );
  OAI22_X1 U88299 ( .A1(n90055), .A2(n120534), .B1(n120749), .B2(n120528), 
        .ZN(n6951) );
  OAI22_X1 U88300 ( .A1(n90054), .A2(n120534), .B1(n120752), .B2(n120528), 
        .ZN(n6952) );
  OAI22_X1 U88301 ( .A1(n90053), .A2(n120534), .B1(n120755), .B2(n120528), 
        .ZN(n6953) );
  OAI22_X1 U88302 ( .A1(n90052), .A2(n120534), .B1(n120758), .B2(n120528), 
        .ZN(n6954) );
  OAI22_X1 U88303 ( .A1(n90051), .A2(n120534), .B1(n120761), .B2(n120528), 
        .ZN(n6955) );
  OAI22_X1 U88304 ( .A1(n90050), .A2(n120534), .B1(n120764), .B2(n120528), 
        .ZN(n6956) );
  OAI22_X1 U88305 ( .A1(n90049), .A2(n120534), .B1(n120767), .B2(n120528), 
        .ZN(n6957) );
  OAI22_X1 U88306 ( .A1(n90048), .A2(n120535), .B1(n120770), .B2(n120528), 
        .ZN(n6958) );
  OAI22_X1 U88307 ( .A1(n90047), .A2(n120535), .B1(n120773), .B2(n120529), 
        .ZN(n6959) );
  OAI22_X1 U88308 ( .A1(n90046), .A2(n120535), .B1(n120776), .B2(n120529), 
        .ZN(n6960) );
  OAI22_X1 U88309 ( .A1(n90045), .A2(n120535), .B1(n120779), .B2(n120529), 
        .ZN(n6961) );
  OAI22_X1 U88310 ( .A1(n90044), .A2(n120535), .B1(n120782), .B2(n120529), 
        .ZN(n6962) );
  OAI22_X1 U88311 ( .A1(n90043), .A2(n120535), .B1(n120785), .B2(n120529), 
        .ZN(n6963) );
  OAI22_X1 U88312 ( .A1(n90042), .A2(n120535), .B1(n120788), .B2(n120529), 
        .ZN(n6964) );
  OAI22_X1 U88313 ( .A1(n90041), .A2(n120535), .B1(n120791), .B2(n120529), 
        .ZN(n6965) );
  OAI22_X1 U88314 ( .A1(n90040), .A2(n120535), .B1(n120794), .B2(n120529), 
        .ZN(n6966) );
  OAI22_X1 U88315 ( .A1(n90039), .A2(n120535), .B1(n120797), .B2(n120529), 
        .ZN(n6967) );
  OAI22_X1 U88316 ( .A1(n90038), .A2(n120535), .B1(n120800), .B2(n120529), 
        .ZN(n6968) );
  OAI22_X1 U88317 ( .A1(n90037), .A2(n120535), .B1(n120803), .B2(n120529), 
        .ZN(n6969) );
  OAI22_X1 U88318 ( .A1(n90036), .A2(n120536), .B1(n120806), .B2(n120529), 
        .ZN(n6970) );
  INV_X1 U88319 ( .A(ADD_RD2[3]), .ZN(n117958) );
  INV_X1 U88320 ( .A(ADD_RD1[4]), .ZN(n116471) );
  INV_X1 U88321 ( .A(ADD_RD2[0]), .ZN(n117967) );
  INV_X1 U88322 ( .A(ADD_RD1[3]), .ZN(n116470) );
  INV_X1 U88323 ( .A(ADD_RD2[4]), .ZN(n117970) );
  INV_X1 U88324 ( .A(ADD_RD1[0]), .ZN(n116469) );
  NAND4_X1 U88325 ( .A1(n117693), .A2(n117694), .A3(n117695), .A4(n117696), 
        .ZN(n5322) );
  AOI221_X1 U88326 ( .B1(n119886), .B2(n118798), .C1(n119880), .C2(n109990), 
        .A(n117713), .ZN(n117694) );
  AOI221_X1 U88327 ( .B1(n119862), .B2(n95440), .C1(n119856), .C2(n118396), 
        .A(n117714), .ZN(n117693) );
  NOR4_X1 U88328 ( .A1(n117709), .A2(n117710), .A3(n117711), .A4(n117712), 
        .ZN(n117695) );
  NAND4_X1 U88329 ( .A1(n117671), .A2(n117672), .A3(n117673), .A4(n117674), 
        .ZN(n5323) );
  AOI221_X1 U88330 ( .B1(n119887), .B2(n118799), .C1(n119881), .C2(n109991), 
        .A(n117691), .ZN(n117672) );
  AOI221_X1 U88331 ( .B1(n119863), .B2(n95441), .C1(n119857), .C2(n118397), 
        .A(n117692), .ZN(n117671) );
  NOR4_X1 U88332 ( .A1(n117687), .A2(n117688), .A3(n117689), .A4(n117690), 
        .ZN(n117673) );
  NAND4_X1 U88333 ( .A1(n117649), .A2(n117650), .A3(n117651), .A4(n117652), 
        .ZN(n5324) );
  AOI221_X1 U88334 ( .B1(n119887), .B2(n118800), .C1(n119881), .C2(n109992), 
        .A(n117669), .ZN(n117650) );
  AOI221_X1 U88335 ( .B1(n119863), .B2(n95442), .C1(n119857), .C2(n118398), 
        .A(n117670), .ZN(n117649) );
  NOR4_X1 U88336 ( .A1(n117665), .A2(n117666), .A3(n117667), .A4(n117668), 
        .ZN(n117651) );
  NAND4_X1 U88337 ( .A1(n117627), .A2(n117628), .A3(n117629), .A4(n117630), 
        .ZN(n5325) );
  AOI221_X1 U88338 ( .B1(n119887), .B2(n118801), .C1(n119881), .C2(n109993), 
        .A(n117647), .ZN(n117628) );
  AOI221_X1 U88339 ( .B1(n119863), .B2(n95443), .C1(n119857), .C2(n118399), 
        .A(n117648), .ZN(n117627) );
  NOR4_X1 U88340 ( .A1(n117643), .A2(n117644), .A3(n117645), .A4(n117646), 
        .ZN(n117629) );
  NAND4_X1 U88341 ( .A1(n117605), .A2(n117606), .A3(n117607), .A4(n117608), 
        .ZN(n5326) );
  AOI221_X1 U88342 ( .B1(n119887), .B2(n118802), .C1(n119881), .C2(n109994), 
        .A(n117625), .ZN(n117606) );
  AOI221_X1 U88343 ( .B1(n119863), .B2(n95444), .C1(n119857), .C2(n118400), 
        .A(n117626), .ZN(n117605) );
  NOR4_X1 U88344 ( .A1(n117621), .A2(n117622), .A3(n117623), .A4(n117624), 
        .ZN(n117607) );
  NAND4_X1 U88345 ( .A1(n117583), .A2(n117584), .A3(n117585), .A4(n117586), 
        .ZN(n5327) );
  AOI221_X1 U88346 ( .B1(n119887), .B2(n118803), .C1(n119881), .C2(n109995), 
        .A(n117603), .ZN(n117584) );
  AOI221_X1 U88347 ( .B1(n119863), .B2(n95445), .C1(n119857), .C2(n118401), 
        .A(n117604), .ZN(n117583) );
  NOR4_X1 U88348 ( .A1(n117599), .A2(n117600), .A3(n117601), .A4(n117602), 
        .ZN(n117585) );
  NAND4_X1 U88349 ( .A1(n117561), .A2(n117562), .A3(n117563), .A4(n117564), 
        .ZN(n5328) );
  AOI221_X1 U88350 ( .B1(n119887), .B2(n118804), .C1(n119881), .C2(n109996), 
        .A(n117581), .ZN(n117562) );
  AOI221_X1 U88351 ( .B1(n119863), .B2(n95446), .C1(n119857), .C2(n118402), 
        .A(n117582), .ZN(n117561) );
  NOR4_X1 U88352 ( .A1(n117577), .A2(n117578), .A3(n117579), .A4(n117580), 
        .ZN(n117563) );
  NAND4_X1 U88353 ( .A1(n117539), .A2(n117540), .A3(n117541), .A4(n117542), 
        .ZN(n5329) );
  AOI221_X1 U88354 ( .B1(n119887), .B2(n118805), .C1(n119881), .C2(n109997), 
        .A(n117559), .ZN(n117540) );
  AOI221_X1 U88355 ( .B1(n119863), .B2(n95447), .C1(n119857), .C2(n118403), 
        .A(n117560), .ZN(n117539) );
  NOR4_X1 U88356 ( .A1(n117555), .A2(n117556), .A3(n117557), .A4(n117558), 
        .ZN(n117541) );
  NAND4_X1 U88357 ( .A1(n117516), .A2(n117517), .A3(n117518), .A4(n117519), 
        .ZN(n5330) );
  AOI221_X1 U88358 ( .B1(n119887), .B2(n118505), .C1(n119881), .C2(n118817), 
        .A(n117537), .ZN(n117517) );
  AOI221_X1 U88359 ( .B1(n119863), .B2(n95448), .C1(n119857), .C2(n118404), 
        .A(n117538), .ZN(n117516) );
  NOR4_X1 U88360 ( .A1(n117532), .A2(n117533), .A3(n117534), .A4(n117535), 
        .ZN(n117518) );
  NAND4_X1 U88361 ( .A1(n117493), .A2(n117494), .A3(n117495), .A4(n117496), 
        .ZN(n5331) );
  AOI221_X1 U88362 ( .B1(n119887), .B2(n118506), .C1(n119881), .C2(n118818), 
        .A(n117514), .ZN(n117494) );
  AOI221_X1 U88363 ( .B1(n119863), .B2(n95449), .C1(n119857), .C2(n118405), 
        .A(n117515), .ZN(n117493) );
  NOR4_X1 U88364 ( .A1(n117509), .A2(n117510), .A3(n117511), .A4(n117512), 
        .ZN(n117495) );
  NAND4_X1 U88365 ( .A1(n117470), .A2(n117471), .A3(n117472), .A4(n117473), 
        .ZN(n5332) );
  AOI221_X1 U88366 ( .B1(n119887), .B2(n118507), .C1(n119881), .C2(n118819), 
        .A(n117491), .ZN(n117471) );
  AOI221_X1 U88367 ( .B1(n119863), .B2(n95450), .C1(n119857), .C2(n118406), 
        .A(n117492), .ZN(n117470) );
  NOR4_X1 U88368 ( .A1(n117486), .A2(n117487), .A3(n117488), .A4(n117489), 
        .ZN(n117472) );
  NAND4_X1 U88369 ( .A1(n117447), .A2(n117448), .A3(n117449), .A4(n117450), 
        .ZN(n5333) );
  AOI221_X1 U88370 ( .B1(n119887), .B2(n118508), .C1(n119881), .C2(n118820), 
        .A(n117468), .ZN(n117448) );
  AOI221_X1 U88371 ( .B1(n119863), .B2(n95451), .C1(n119857), .C2(n118407), 
        .A(n117469), .ZN(n117447) );
  NOR4_X1 U88372 ( .A1(n117463), .A2(n117464), .A3(n117465), .A4(n117466), 
        .ZN(n117449) );
  NAND4_X1 U88373 ( .A1(n117424), .A2(n117425), .A3(n117426), .A4(n117427), 
        .ZN(n5334) );
  AOI221_X1 U88374 ( .B1(n119887), .B2(n118509), .C1(n119881), .C2(n118821), 
        .A(n117445), .ZN(n117425) );
  AOI221_X1 U88375 ( .B1(n119863), .B2(n95452), .C1(n119857), .C2(n118408), 
        .A(n117446), .ZN(n117424) );
  NOR4_X1 U88376 ( .A1(n117440), .A2(n117441), .A3(n117442), .A4(n117443), 
        .ZN(n117426) );
  NAND4_X1 U88377 ( .A1(n117401), .A2(n117402), .A3(n117403), .A4(n117404), 
        .ZN(n5335) );
  AOI221_X1 U88378 ( .B1(n119888), .B2(n118510), .C1(n119882), .C2(n118822), 
        .A(n117422), .ZN(n117402) );
  AOI221_X1 U88379 ( .B1(n119864), .B2(n95453), .C1(n119858), .C2(n118409), 
        .A(n117423), .ZN(n117401) );
  NOR4_X1 U88380 ( .A1(n117417), .A2(n117418), .A3(n117419), .A4(n117420), 
        .ZN(n117403) );
  NAND4_X1 U88381 ( .A1(n117378), .A2(n117379), .A3(n117380), .A4(n117381), 
        .ZN(n5336) );
  AOI221_X1 U88382 ( .B1(n119888), .B2(n118511), .C1(n119882), .C2(n118823), 
        .A(n117399), .ZN(n117379) );
  AOI221_X1 U88383 ( .B1(n119864), .B2(n95454), .C1(n119858), .C2(n118410), 
        .A(n117400), .ZN(n117378) );
  NOR4_X1 U88384 ( .A1(n117394), .A2(n117395), .A3(n117396), .A4(n117397), 
        .ZN(n117380) );
  NAND4_X1 U88385 ( .A1(n117355), .A2(n117356), .A3(n117357), .A4(n117358), 
        .ZN(n5337) );
  AOI221_X1 U88386 ( .B1(n119888), .B2(n118512), .C1(n119882), .C2(n118824), 
        .A(n117376), .ZN(n117356) );
  AOI221_X1 U88387 ( .B1(n119864), .B2(n95455), .C1(n119858), .C2(n118411), 
        .A(n117377), .ZN(n117355) );
  NOR4_X1 U88388 ( .A1(n117371), .A2(n117372), .A3(n117373), .A4(n117374), 
        .ZN(n117357) );
  NAND4_X1 U88389 ( .A1(n117332), .A2(n117333), .A3(n117334), .A4(n117335), 
        .ZN(n5338) );
  AOI221_X1 U88390 ( .B1(n119888), .B2(n118513), .C1(n119882), .C2(n118825), 
        .A(n117353), .ZN(n117333) );
  AOI221_X1 U88391 ( .B1(n119864), .B2(n95456), .C1(n119858), .C2(n118412), 
        .A(n117354), .ZN(n117332) );
  NOR4_X1 U88392 ( .A1(n117348), .A2(n117349), .A3(n117350), .A4(n117351), 
        .ZN(n117334) );
  NAND4_X1 U88393 ( .A1(n117309), .A2(n117310), .A3(n117311), .A4(n117312), 
        .ZN(n5339) );
  AOI221_X1 U88394 ( .B1(n119888), .B2(n118514), .C1(n119882), .C2(n118826), 
        .A(n117330), .ZN(n117310) );
  AOI221_X1 U88395 ( .B1(n119864), .B2(n95457), .C1(n119858), .C2(n118413), 
        .A(n117331), .ZN(n117309) );
  NOR4_X1 U88396 ( .A1(n117325), .A2(n117326), .A3(n117327), .A4(n117328), 
        .ZN(n117311) );
  NAND4_X1 U88397 ( .A1(n117286), .A2(n117287), .A3(n117288), .A4(n117289), 
        .ZN(n5340) );
  AOI221_X1 U88398 ( .B1(n119888), .B2(n118515), .C1(n119882), .C2(n118827), 
        .A(n117307), .ZN(n117287) );
  AOI221_X1 U88399 ( .B1(n119864), .B2(n95458), .C1(n119858), .C2(n118414), 
        .A(n117308), .ZN(n117286) );
  NOR4_X1 U88400 ( .A1(n117302), .A2(n117303), .A3(n117304), .A4(n117305), 
        .ZN(n117288) );
  NAND4_X1 U88401 ( .A1(n117263), .A2(n117264), .A3(n117265), .A4(n117266), 
        .ZN(n5341) );
  AOI221_X1 U88402 ( .B1(n119888), .B2(n118516), .C1(n119882), .C2(n118828), 
        .A(n117284), .ZN(n117264) );
  AOI221_X1 U88403 ( .B1(n119864), .B2(n95459), .C1(n119858), .C2(n118415), 
        .A(n117285), .ZN(n117263) );
  NOR4_X1 U88404 ( .A1(n117279), .A2(n117280), .A3(n117281), .A4(n117282), 
        .ZN(n117265) );
  NAND4_X1 U88405 ( .A1(n117240), .A2(n117241), .A3(n117242), .A4(n117243), 
        .ZN(n5342) );
  AOI221_X1 U88406 ( .B1(n119888), .B2(n118517), .C1(n119882), .C2(n118829), 
        .A(n117261), .ZN(n117241) );
  AOI221_X1 U88407 ( .B1(n119864), .B2(n95460), .C1(n119858), .C2(n118416), 
        .A(n117262), .ZN(n117240) );
  NOR4_X1 U88408 ( .A1(n117256), .A2(n117257), .A3(n117258), .A4(n117259), 
        .ZN(n117242) );
  NAND4_X1 U88409 ( .A1(n117217), .A2(n117218), .A3(n117219), .A4(n117220), 
        .ZN(n5343) );
  AOI221_X1 U88410 ( .B1(n119888), .B2(n118518), .C1(n119882), .C2(n118830), 
        .A(n117238), .ZN(n117218) );
  AOI221_X1 U88411 ( .B1(n119864), .B2(n95461), .C1(n119858), .C2(n118417), 
        .A(n117239), .ZN(n117217) );
  NOR4_X1 U88412 ( .A1(n117233), .A2(n117234), .A3(n117235), .A4(n117236), 
        .ZN(n117219) );
  NAND4_X1 U88413 ( .A1(n117194), .A2(n117195), .A3(n117196), .A4(n117197), 
        .ZN(n5344) );
  AOI221_X1 U88414 ( .B1(n119888), .B2(n118519), .C1(n119882), .C2(n118831), 
        .A(n117215), .ZN(n117195) );
  AOI221_X1 U88415 ( .B1(n119864), .B2(n95462), .C1(n119858), .C2(n118418), 
        .A(n117216), .ZN(n117194) );
  NOR4_X1 U88416 ( .A1(n117210), .A2(n117211), .A3(n117212), .A4(n117213), 
        .ZN(n117196) );
  NAND4_X1 U88417 ( .A1(n117171), .A2(n117172), .A3(n117173), .A4(n117174), 
        .ZN(n5345) );
  AOI221_X1 U88418 ( .B1(n119888), .B2(n118520), .C1(n119882), .C2(n118832), 
        .A(n117192), .ZN(n117172) );
  AOI221_X1 U88419 ( .B1(n119864), .B2(n95463), .C1(n119858), .C2(n118419), 
        .A(n117193), .ZN(n117171) );
  NOR4_X1 U88420 ( .A1(n117187), .A2(n117188), .A3(n117189), .A4(n117190), 
        .ZN(n117173) );
  NAND4_X1 U88421 ( .A1(n117148), .A2(n117149), .A3(n117150), .A4(n117151), 
        .ZN(n5346) );
  AOI221_X1 U88422 ( .B1(n119888), .B2(n118521), .C1(n119882), .C2(n118833), 
        .A(n117169), .ZN(n117149) );
  AOI221_X1 U88423 ( .B1(n119864), .B2(n95464), .C1(n119858), .C2(n118420), 
        .A(n117170), .ZN(n117148) );
  NOR4_X1 U88424 ( .A1(n117164), .A2(n117165), .A3(n117166), .A4(n117167), 
        .ZN(n117150) );
  NAND4_X1 U88425 ( .A1(n117125), .A2(n117126), .A3(n117127), .A4(n117128), 
        .ZN(n5347) );
  AOI221_X1 U88426 ( .B1(n119889), .B2(n118522), .C1(n119883), .C2(n118834), 
        .A(n117146), .ZN(n117126) );
  AOI221_X1 U88427 ( .B1(n119865), .B2(n95465), .C1(n119859), .C2(n118421), 
        .A(n117147), .ZN(n117125) );
  NOR4_X1 U88428 ( .A1(n117141), .A2(n117142), .A3(n117143), .A4(n117144), 
        .ZN(n117127) );
  NAND4_X1 U88429 ( .A1(n117102), .A2(n117103), .A3(n117104), .A4(n117105), 
        .ZN(n5348) );
  AOI221_X1 U88430 ( .B1(n119889), .B2(n118523), .C1(n119883), .C2(n118835), 
        .A(n117123), .ZN(n117103) );
  AOI221_X1 U88431 ( .B1(n119865), .B2(n95466), .C1(n119859), .C2(n118422), 
        .A(n117124), .ZN(n117102) );
  NOR4_X1 U88432 ( .A1(n117118), .A2(n117119), .A3(n117120), .A4(n117121), 
        .ZN(n117104) );
  NAND4_X1 U88433 ( .A1(n117079), .A2(n117080), .A3(n117081), .A4(n117082), 
        .ZN(n5349) );
  AOI221_X1 U88434 ( .B1(n119889), .B2(n118524), .C1(n119883), .C2(n118836), 
        .A(n117100), .ZN(n117080) );
  AOI221_X1 U88435 ( .B1(n119865), .B2(n95467), .C1(n119859), .C2(n118423), 
        .A(n117101), .ZN(n117079) );
  NOR4_X1 U88436 ( .A1(n117095), .A2(n117096), .A3(n117097), .A4(n117098), 
        .ZN(n117081) );
  NAND4_X1 U88437 ( .A1(n117056), .A2(n117057), .A3(n117058), .A4(n117059), 
        .ZN(n5350) );
  AOI221_X1 U88438 ( .B1(n119889), .B2(n118525), .C1(n119883), .C2(n118837), 
        .A(n117077), .ZN(n117057) );
  AOI221_X1 U88439 ( .B1(n119865), .B2(n95468), .C1(n119859), .C2(n118424), 
        .A(n117078), .ZN(n117056) );
  NOR4_X1 U88440 ( .A1(n117072), .A2(n117073), .A3(n117074), .A4(n117075), 
        .ZN(n117058) );
  NAND4_X1 U88441 ( .A1(n117033), .A2(n117034), .A3(n117035), .A4(n117036), 
        .ZN(n5351) );
  AOI221_X1 U88442 ( .B1(n119889), .B2(n118526), .C1(n119883), .C2(n118838), 
        .A(n117054), .ZN(n117034) );
  AOI221_X1 U88443 ( .B1(n119865), .B2(n95469), .C1(n119859), .C2(n118425), 
        .A(n117055), .ZN(n117033) );
  NOR4_X1 U88444 ( .A1(n117049), .A2(n117050), .A3(n117051), .A4(n117052), 
        .ZN(n117035) );
  NAND4_X1 U88445 ( .A1(n117010), .A2(n117011), .A3(n117012), .A4(n117013), 
        .ZN(n5352) );
  AOI221_X1 U88446 ( .B1(n119889), .B2(n118527), .C1(n119883), .C2(n118839), 
        .A(n117031), .ZN(n117011) );
  AOI221_X1 U88447 ( .B1(n119865), .B2(n95470), .C1(n119859), .C2(n118426), 
        .A(n117032), .ZN(n117010) );
  NOR4_X1 U88448 ( .A1(n117026), .A2(n117027), .A3(n117028), .A4(n117029), 
        .ZN(n117012) );
  NAND4_X1 U88449 ( .A1(n116987), .A2(n116988), .A3(n116989), .A4(n116990), 
        .ZN(n5353) );
  AOI221_X1 U88450 ( .B1(n119889), .B2(n118528), .C1(n119883), .C2(n118840), 
        .A(n117008), .ZN(n116988) );
  AOI221_X1 U88451 ( .B1(n119865), .B2(n95471), .C1(n119859), .C2(n118427), 
        .A(n117009), .ZN(n116987) );
  NOR4_X1 U88452 ( .A1(n117003), .A2(n117004), .A3(n117005), .A4(n117006), 
        .ZN(n116989) );
  NAND4_X1 U88453 ( .A1(n116964), .A2(n116965), .A3(n116966), .A4(n116967), 
        .ZN(n5354) );
  AOI221_X1 U88454 ( .B1(n119889), .B2(n118529), .C1(n119883), .C2(n118841), 
        .A(n116985), .ZN(n116965) );
  AOI221_X1 U88455 ( .B1(n119865), .B2(n95472), .C1(n119859), .C2(n118428), 
        .A(n116986), .ZN(n116964) );
  NOR4_X1 U88456 ( .A1(n116980), .A2(n116981), .A3(n116982), .A4(n116983), 
        .ZN(n116966) );
  NAND4_X1 U88457 ( .A1(n116941), .A2(n116942), .A3(n116943), .A4(n116944), 
        .ZN(n5355) );
  AOI221_X1 U88458 ( .B1(n119889), .B2(n118530), .C1(n119883), .C2(n118842), 
        .A(n116962), .ZN(n116942) );
  AOI221_X1 U88459 ( .B1(n119865), .B2(n95473), .C1(n119859), .C2(n118429), 
        .A(n116963), .ZN(n116941) );
  NOR4_X1 U88460 ( .A1(n116957), .A2(n116958), .A3(n116959), .A4(n116960), 
        .ZN(n116943) );
  NAND4_X1 U88461 ( .A1(n116918), .A2(n116919), .A3(n116920), .A4(n116921), 
        .ZN(n5356) );
  AOI221_X1 U88462 ( .B1(n119889), .B2(n118531), .C1(n119883), .C2(n118843), 
        .A(n116939), .ZN(n116919) );
  AOI221_X1 U88463 ( .B1(n119865), .B2(n95474), .C1(n119859), .C2(n118430), 
        .A(n116940), .ZN(n116918) );
  NOR4_X1 U88464 ( .A1(n116934), .A2(n116935), .A3(n116936), .A4(n116937), 
        .ZN(n116920) );
  NAND4_X1 U88465 ( .A1(n116895), .A2(n116896), .A3(n116897), .A4(n116898), 
        .ZN(n5357) );
  AOI221_X1 U88466 ( .B1(n119889), .B2(n118532), .C1(n119883), .C2(n118844), 
        .A(n116916), .ZN(n116896) );
  AOI221_X1 U88467 ( .B1(n119865), .B2(n95475), .C1(n119859), .C2(n118431), 
        .A(n116917), .ZN(n116895) );
  NOR4_X1 U88468 ( .A1(n116911), .A2(n116912), .A3(n116913), .A4(n116914), 
        .ZN(n116897) );
  NAND4_X1 U88469 ( .A1(n116872), .A2(n116873), .A3(n116874), .A4(n116875), 
        .ZN(n5358) );
  AOI221_X1 U88470 ( .B1(n119889), .B2(n118533), .C1(n119883), .C2(n118845), 
        .A(n116893), .ZN(n116873) );
  AOI221_X1 U88471 ( .B1(n119865), .B2(n95476), .C1(n119859), .C2(n118432), 
        .A(n116894), .ZN(n116872) );
  NOR4_X1 U88472 ( .A1(n116888), .A2(n116889), .A3(n116890), .A4(n116891), 
        .ZN(n116874) );
  NAND4_X1 U88473 ( .A1(n116849), .A2(n116850), .A3(n116851), .A4(n116852), 
        .ZN(n5359) );
  AOI221_X1 U88474 ( .B1(n119890), .B2(n118534), .C1(n119884), .C2(n118846), 
        .A(n116870), .ZN(n116850) );
  AOI221_X1 U88475 ( .B1(n119866), .B2(n95477), .C1(n119860), .C2(n118433), 
        .A(n116871), .ZN(n116849) );
  NOR4_X1 U88476 ( .A1(n116865), .A2(n116866), .A3(n116867), .A4(n116868), 
        .ZN(n116851) );
  NAND4_X1 U88477 ( .A1(n116826), .A2(n116827), .A3(n116828), .A4(n116829), 
        .ZN(n5360) );
  AOI221_X1 U88478 ( .B1(n119890), .B2(n118535), .C1(n119884), .C2(n118847), 
        .A(n116847), .ZN(n116827) );
  AOI221_X1 U88479 ( .B1(n119866), .B2(n95478), .C1(n119860), .C2(n118434), 
        .A(n116848), .ZN(n116826) );
  NOR4_X1 U88480 ( .A1(n116842), .A2(n116843), .A3(n116844), .A4(n116845), 
        .ZN(n116828) );
  NAND4_X1 U88481 ( .A1(n116803), .A2(n116804), .A3(n116805), .A4(n116806), 
        .ZN(n5361) );
  AOI221_X1 U88482 ( .B1(n119890), .B2(n118536), .C1(n119884), .C2(n118848), 
        .A(n116824), .ZN(n116804) );
  AOI221_X1 U88483 ( .B1(n119866), .B2(n95479), .C1(n119860), .C2(n118435), 
        .A(n116825), .ZN(n116803) );
  NOR4_X1 U88484 ( .A1(n116819), .A2(n116820), .A3(n116821), .A4(n116822), 
        .ZN(n116805) );
  NAND4_X1 U88485 ( .A1(n116780), .A2(n116781), .A3(n116782), .A4(n116783), 
        .ZN(n5362) );
  AOI221_X1 U88486 ( .B1(n119890), .B2(n118537), .C1(n119884), .C2(n118849), 
        .A(n116801), .ZN(n116781) );
  AOI221_X1 U88487 ( .B1(n119866), .B2(n95480), .C1(n119860), .C2(n118436), 
        .A(n116802), .ZN(n116780) );
  NOR4_X1 U88488 ( .A1(n116796), .A2(n116797), .A3(n116798), .A4(n116799), 
        .ZN(n116782) );
  NAND4_X1 U88489 ( .A1(n116757), .A2(n116758), .A3(n116759), .A4(n116760), 
        .ZN(n5363) );
  AOI221_X1 U88490 ( .B1(n119890), .B2(n118538), .C1(n119884), .C2(n118850), 
        .A(n116778), .ZN(n116758) );
  AOI221_X1 U88491 ( .B1(n119866), .B2(n95481), .C1(n119860), .C2(n118437), 
        .A(n116779), .ZN(n116757) );
  NOR4_X1 U88492 ( .A1(n116773), .A2(n116774), .A3(n116775), .A4(n116776), 
        .ZN(n116759) );
  NAND4_X1 U88493 ( .A1(n116734), .A2(n116735), .A3(n116736), .A4(n116737), 
        .ZN(n5364) );
  AOI221_X1 U88494 ( .B1(n119890), .B2(n118539), .C1(n119884), .C2(n118851), 
        .A(n116755), .ZN(n116735) );
  AOI221_X1 U88495 ( .B1(n119866), .B2(n95482), .C1(n119860), .C2(n118438), 
        .A(n116756), .ZN(n116734) );
  NOR4_X1 U88496 ( .A1(n116750), .A2(n116751), .A3(n116752), .A4(n116753), 
        .ZN(n116736) );
  NAND4_X1 U88497 ( .A1(n116711), .A2(n116712), .A3(n116713), .A4(n116714), 
        .ZN(n5365) );
  AOI221_X1 U88498 ( .B1(n119890), .B2(n118540), .C1(n119884), .C2(n118852), 
        .A(n116732), .ZN(n116712) );
  AOI221_X1 U88499 ( .B1(n119866), .B2(n95483), .C1(n119860), .C2(n118439), 
        .A(n116733), .ZN(n116711) );
  NOR4_X1 U88500 ( .A1(n116727), .A2(n116728), .A3(n116729), .A4(n116730), 
        .ZN(n116713) );
  NAND4_X1 U88501 ( .A1(n116688), .A2(n116689), .A3(n116690), .A4(n116691), 
        .ZN(n5366) );
  AOI221_X1 U88502 ( .B1(n119890), .B2(n118541), .C1(n119884), .C2(n118853), 
        .A(n116709), .ZN(n116689) );
  AOI221_X1 U88503 ( .B1(n119866), .B2(n95484), .C1(n119860), .C2(n118440), 
        .A(n116710), .ZN(n116688) );
  NOR4_X1 U88504 ( .A1(n116704), .A2(n116705), .A3(n116706), .A4(n116707), 
        .ZN(n116690) );
  NAND4_X1 U88505 ( .A1(n116665), .A2(n116666), .A3(n116667), .A4(n116668), 
        .ZN(n5367) );
  AOI221_X1 U88506 ( .B1(n119890), .B2(n118542), .C1(n119884), .C2(n118854), 
        .A(n116686), .ZN(n116666) );
  AOI221_X1 U88507 ( .B1(n119866), .B2(n95485), .C1(n119860), .C2(n118441), 
        .A(n116687), .ZN(n116665) );
  NOR4_X1 U88508 ( .A1(n116681), .A2(n116682), .A3(n116683), .A4(n116684), 
        .ZN(n116667) );
  NAND4_X1 U88509 ( .A1(n116642), .A2(n116643), .A3(n116644), .A4(n116645), 
        .ZN(n5368) );
  AOI221_X1 U88510 ( .B1(n119890), .B2(n118543), .C1(n119884), .C2(n118855), 
        .A(n116663), .ZN(n116643) );
  AOI221_X1 U88511 ( .B1(n119866), .B2(n95486), .C1(n119860), .C2(n118442), 
        .A(n116664), .ZN(n116642) );
  NOR4_X1 U88512 ( .A1(n116658), .A2(n116659), .A3(n116660), .A4(n116661), 
        .ZN(n116644) );
  NAND4_X1 U88513 ( .A1(n116619), .A2(n116620), .A3(n116621), .A4(n116622), 
        .ZN(n5369) );
  AOI221_X1 U88514 ( .B1(n119890), .B2(n118544), .C1(n119884), .C2(n118856), 
        .A(n116640), .ZN(n116620) );
  AOI221_X1 U88515 ( .B1(n119866), .B2(n95487), .C1(n119860), .C2(n118443), 
        .A(n116641), .ZN(n116619) );
  NOR4_X1 U88516 ( .A1(n116635), .A2(n116636), .A3(n116637), .A4(n116638), 
        .ZN(n116621) );
  NAND4_X1 U88517 ( .A1(n116596), .A2(n116597), .A3(n116598), .A4(n116599), 
        .ZN(n5370) );
  AOI221_X1 U88518 ( .B1(n119890), .B2(n118545), .C1(n119884), .C2(n118857), 
        .A(n116617), .ZN(n116597) );
  AOI221_X1 U88519 ( .B1(n119866), .B2(n95488), .C1(n119860), .C2(n118444), 
        .A(n116618), .ZN(n116596) );
  NOR4_X1 U88520 ( .A1(n116612), .A2(n116613), .A3(n116614), .A4(n116615), 
        .ZN(n116598) );
  NAND4_X1 U88521 ( .A1(n114757), .A2(n114758), .A3(n114759), .A4(n114760), 
        .ZN(n5495) );
  AOI221_X1 U88522 ( .B1(n120065), .B2(n119174), .C1(n120059), .C2(n117985), 
        .A(n114781), .ZN(n114757) );
  NOR4_X1 U88523 ( .A1(n114761), .A2(n114762), .A3(n114763), .A4(n114764), 
        .ZN(n114760) );
  NOR4_X1 U88524 ( .A1(n114773), .A2(n114774), .A3(n114775), .A4(n114776), 
        .ZN(n114759) );
  NAND4_X1 U88525 ( .A1(n114731), .A2(n114732), .A3(n114733), .A4(n114734), 
        .ZN(n5497) );
  AOI221_X1 U88526 ( .B1(n120065), .B2(n119175), .C1(n120059), .C2(n117986), 
        .A(n114755), .ZN(n114731) );
  NOR4_X1 U88527 ( .A1(n114735), .A2(n114736), .A3(n114737), .A4(n114738), 
        .ZN(n114734) );
  NOR4_X1 U88528 ( .A1(n114747), .A2(n114748), .A3(n114749), .A4(n114750), 
        .ZN(n114733) );
  NAND4_X1 U88529 ( .A1(n114705), .A2(n114706), .A3(n114707), .A4(n114708), 
        .ZN(n5499) );
  AOI221_X1 U88530 ( .B1(n120065), .B2(n119176), .C1(n120059), .C2(n117987), 
        .A(n114729), .ZN(n114705) );
  NOR4_X1 U88531 ( .A1(n114709), .A2(n114710), .A3(n114711), .A4(n114712), 
        .ZN(n114708) );
  NOR4_X1 U88532 ( .A1(n114721), .A2(n114722), .A3(n114723), .A4(n114724), 
        .ZN(n114707) );
  NAND4_X1 U88533 ( .A1(n114646), .A2(n114647), .A3(n114648), .A4(n114649), 
        .ZN(n5501) );
  AOI221_X1 U88534 ( .B1(n120065), .B2(n119177), .C1(n120059), .C2(n117988), 
        .A(n114701), .ZN(n114646) );
  NOR4_X1 U88535 ( .A1(n114650), .A2(n114651), .A3(n114652), .A4(n114653), 
        .ZN(n114649) );
  NOR4_X1 U88536 ( .A1(n114678), .A2(n114679), .A3(n114680), .A4(n114681), 
        .ZN(n114648) );
  NAND4_X1 U88537 ( .A1(n116575), .A2(n116576), .A3(n116577), .A4(n116578), 
        .ZN(n5371) );
  NOR4_X1 U88538 ( .A1(n116589), .A2(n116590), .A3(n116591), .A4(n116592), 
        .ZN(n116577) );
  AOI221_X1 U88539 ( .B1(n119891), .B2(n109895), .C1(n119885), .C2(n118858), 
        .A(n116594), .ZN(n116576) );
  NOR4_X1 U88540 ( .A1(n116579), .A2(n116580), .A3(n116581), .A4(n116582), 
        .ZN(n116578) );
  NAND4_X1 U88541 ( .A1(n116554), .A2(n116555), .A3(n116556), .A4(n116557), 
        .ZN(n5372) );
  NOR4_X1 U88542 ( .A1(n116568), .A2(n116569), .A3(n116570), .A4(n116571), 
        .ZN(n116556) );
  AOI221_X1 U88543 ( .B1(n119891), .B2(n109896), .C1(n119885), .C2(n118859), 
        .A(n116573), .ZN(n116555) );
  NOR4_X1 U88544 ( .A1(n116558), .A2(n116559), .A3(n116560), .A4(n116561), 
        .ZN(n116557) );
  NAND4_X1 U88545 ( .A1(n116533), .A2(n116534), .A3(n116535), .A4(n116536), 
        .ZN(n5373) );
  NOR4_X1 U88546 ( .A1(n116547), .A2(n116548), .A3(n116549), .A4(n116550), 
        .ZN(n116535) );
  AOI221_X1 U88547 ( .B1(n119891), .B2(n109897), .C1(n119885), .C2(n118860), 
        .A(n116552), .ZN(n116534) );
  NOR4_X1 U88548 ( .A1(n116537), .A2(n116538), .A3(n116539), .A4(n116540), 
        .ZN(n116536) );
  NAND4_X1 U88549 ( .A1(n116479), .A2(n116480), .A3(n116481), .A4(n116482), 
        .ZN(n5374) );
  NOR4_X1 U88550 ( .A1(n116509), .A2(n116510), .A3(n116511), .A4(n116512), 
        .ZN(n116481) );
  AOI221_X1 U88551 ( .B1(n119891), .B2(n109898), .C1(n119885), .C2(n118861), 
        .A(n116525), .ZN(n116480) );
  NOR4_X1 U88552 ( .A1(n116483), .A2(n116484), .A3(n116485), .A4(n116486), 
        .ZN(n116482) );
  NAND4_X1 U88553 ( .A1(n115147), .A2(n115148), .A3(n115149), .A4(n115150), 
        .ZN(n5467) );
  AOI221_X1 U88554 ( .B1(n120063), .B2(n119178), .C1(n120057), .C2(n118431), 
        .A(n115173), .ZN(n115147) );
  AOI221_X1 U88555 ( .B1(n120087), .B2(n118986), .C1(n120081), .C2(n118550), 
        .A(n115171), .ZN(n115148) );
  NOR4_X1 U88556 ( .A1(n115165), .A2(n115166), .A3(n115167), .A4(n115168), 
        .ZN(n115149) );
  NAND4_X1 U88557 ( .A1(n115119), .A2(n115120), .A3(n115121), .A4(n115122), 
        .ZN(n5469) );
  AOI221_X1 U88558 ( .B1(n120063), .B2(n119179), .C1(n120057), .C2(n118432), 
        .A(n115145), .ZN(n115119) );
  AOI221_X1 U88559 ( .B1(n120087), .B2(n118987), .C1(n120081), .C2(n118551), 
        .A(n115143), .ZN(n115120) );
  NOR4_X1 U88560 ( .A1(n115137), .A2(n115138), .A3(n115139), .A4(n115140), 
        .ZN(n115121) );
  NAND4_X1 U88561 ( .A1(n115091), .A2(n115092), .A3(n115093), .A4(n115094), 
        .ZN(n5471) );
  AOI221_X1 U88562 ( .B1(n120064), .B2(n119180), .C1(n120058), .C2(n118433), 
        .A(n115117), .ZN(n115091) );
  AOI221_X1 U88563 ( .B1(n120088), .B2(n118988), .C1(n120082), .C2(n118552), 
        .A(n115115), .ZN(n115092) );
  NOR4_X1 U88564 ( .A1(n115109), .A2(n115110), .A3(n115111), .A4(n115112), 
        .ZN(n115093) );
  NAND4_X1 U88565 ( .A1(n115063), .A2(n115064), .A3(n115065), .A4(n115066), 
        .ZN(n5473) );
  AOI221_X1 U88566 ( .B1(n120064), .B2(n119181), .C1(n120058), .C2(n118434), 
        .A(n115089), .ZN(n115063) );
  AOI221_X1 U88567 ( .B1(n120088), .B2(n118989), .C1(n120082), .C2(n118553), 
        .A(n115087), .ZN(n115064) );
  NOR4_X1 U88568 ( .A1(n115081), .A2(n115082), .A3(n115083), .A4(n115084), 
        .ZN(n115065) );
  NAND4_X1 U88569 ( .A1(n115035), .A2(n115036), .A3(n115037), .A4(n115038), 
        .ZN(n5475) );
  AOI221_X1 U88570 ( .B1(n120064), .B2(n119182), .C1(n120058), .C2(n118435), 
        .A(n115061), .ZN(n115035) );
  AOI221_X1 U88571 ( .B1(n120088), .B2(n118990), .C1(n120082), .C2(n118554), 
        .A(n115059), .ZN(n115036) );
  NOR4_X1 U88572 ( .A1(n115053), .A2(n115054), .A3(n115055), .A4(n115056), 
        .ZN(n115037) );
  NAND4_X1 U88573 ( .A1(n115007), .A2(n115008), .A3(n115009), .A4(n115010), 
        .ZN(n5477) );
  AOI221_X1 U88574 ( .B1(n120064), .B2(n119183), .C1(n120058), .C2(n118436), 
        .A(n115033), .ZN(n115007) );
  AOI221_X1 U88575 ( .B1(n120088), .B2(n118991), .C1(n120082), .C2(n118555), 
        .A(n115031), .ZN(n115008) );
  NOR4_X1 U88576 ( .A1(n115025), .A2(n115026), .A3(n115027), .A4(n115028), 
        .ZN(n115009) );
  NAND4_X1 U88577 ( .A1(n114979), .A2(n114980), .A3(n114981), .A4(n114982), 
        .ZN(n5479) );
  AOI221_X1 U88578 ( .B1(n120064), .B2(n119184), .C1(n120058), .C2(n118437), 
        .A(n115005), .ZN(n114979) );
  AOI221_X1 U88579 ( .B1(n120088), .B2(n118992), .C1(n120082), .C2(n118556), 
        .A(n115003), .ZN(n114980) );
  NOR4_X1 U88580 ( .A1(n114997), .A2(n114998), .A3(n114999), .A4(n115000), 
        .ZN(n114981) );
  NAND4_X1 U88581 ( .A1(n114951), .A2(n114952), .A3(n114953), .A4(n114954), 
        .ZN(n5481) );
  AOI221_X1 U88582 ( .B1(n120064), .B2(n119185), .C1(n120058), .C2(n118438), 
        .A(n114977), .ZN(n114951) );
  AOI221_X1 U88583 ( .B1(n120088), .B2(n118993), .C1(n120082), .C2(n118557), 
        .A(n114975), .ZN(n114952) );
  NOR4_X1 U88584 ( .A1(n114969), .A2(n114970), .A3(n114971), .A4(n114972), 
        .ZN(n114953) );
  NAND4_X1 U88585 ( .A1(n114923), .A2(n114924), .A3(n114925), .A4(n114926), 
        .ZN(n5483) );
  AOI221_X1 U88586 ( .B1(n120064), .B2(n119186), .C1(n120058), .C2(n118439), 
        .A(n114949), .ZN(n114923) );
  AOI221_X1 U88587 ( .B1(n120088), .B2(n118994), .C1(n120082), .C2(n118558), 
        .A(n114947), .ZN(n114924) );
  NOR4_X1 U88588 ( .A1(n114941), .A2(n114942), .A3(n114943), .A4(n114944), 
        .ZN(n114925) );
  NAND4_X1 U88589 ( .A1(n114895), .A2(n114896), .A3(n114897), .A4(n114898), 
        .ZN(n5485) );
  AOI221_X1 U88590 ( .B1(n120064), .B2(n119187), .C1(n120058), .C2(n118440), 
        .A(n114921), .ZN(n114895) );
  AOI221_X1 U88591 ( .B1(n120088), .B2(n118995), .C1(n120082), .C2(n118559), 
        .A(n114919), .ZN(n114896) );
  NOR4_X1 U88592 ( .A1(n114913), .A2(n114914), .A3(n114915), .A4(n114916), 
        .ZN(n114897) );
  NAND4_X1 U88593 ( .A1(n114867), .A2(n114868), .A3(n114869), .A4(n114870), 
        .ZN(n5487) );
  AOI221_X1 U88594 ( .B1(n120064), .B2(n119188), .C1(n120058), .C2(n118441), 
        .A(n114893), .ZN(n114867) );
  AOI221_X1 U88595 ( .B1(n120088), .B2(n118996), .C1(n120082), .C2(n118560), 
        .A(n114891), .ZN(n114868) );
  NOR4_X1 U88596 ( .A1(n114885), .A2(n114886), .A3(n114887), .A4(n114888), 
        .ZN(n114869) );
  NAND4_X1 U88597 ( .A1(n114839), .A2(n114840), .A3(n114841), .A4(n114842), 
        .ZN(n5489) );
  AOI221_X1 U88598 ( .B1(n120064), .B2(n119189), .C1(n120058), .C2(n118442), 
        .A(n114865), .ZN(n114839) );
  AOI221_X1 U88599 ( .B1(n120088), .B2(n118997), .C1(n120082), .C2(n118561), 
        .A(n114863), .ZN(n114840) );
  NOR4_X1 U88600 ( .A1(n114857), .A2(n114858), .A3(n114859), .A4(n114860), 
        .ZN(n114841) );
  NAND4_X1 U88601 ( .A1(n114811), .A2(n114812), .A3(n114813), .A4(n114814), 
        .ZN(n5491) );
  AOI221_X1 U88602 ( .B1(n120064), .B2(n119190), .C1(n120058), .C2(n118443), 
        .A(n114837), .ZN(n114811) );
  AOI221_X1 U88603 ( .B1(n120088), .B2(n118998), .C1(n120082), .C2(n118562), 
        .A(n114835), .ZN(n114812) );
  NOR4_X1 U88604 ( .A1(n114829), .A2(n114830), .A3(n114831), .A4(n114832), 
        .ZN(n114813) );
  NAND4_X1 U88605 ( .A1(n114783), .A2(n114784), .A3(n114785), .A4(n114786), 
        .ZN(n5493) );
  AOI221_X1 U88606 ( .B1(n120064), .B2(n119191), .C1(n120058), .C2(n118444), 
        .A(n114809), .ZN(n114783) );
  AOI221_X1 U88607 ( .B1(n120088), .B2(n118999), .C1(n120082), .C2(n118563), 
        .A(n114807), .ZN(n114784) );
  NOR4_X1 U88608 ( .A1(n114801), .A2(n114802), .A3(n114803), .A4(n114804), 
        .ZN(n114785) );
  NAND4_X1 U88609 ( .A1(n116435), .A2(n116436), .A3(n116437), .A4(n116438), 
        .ZN(n5375) );
  AOI221_X1 U88610 ( .B1(n120060), .B2(n119192), .C1(n120054), .C2(n118385), 
        .A(n116477), .ZN(n116435) );
  AOI221_X1 U88611 ( .B1(n120084), .B2(n119000), .C1(n120078), .C2(n118564), 
        .A(n116474), .ZN(n116436) );
  NOR4_X1 U88612 ( .A1(n116465), .A2(n116466), .A3(n116467), .A4(n116468), 
        .ZN(n116437) );
  NAND4_X1 U88613 ( .A1(n116407), .A2(n116408), .A3(n116409), .A4(n116410), 
        .ZN(n5377) );
  AOI221_X1 U88614 ( .B1(n120060), .B2(n119193), .C1(n120054), .C2(n118386), 
        .A(n116433), .ZN(n116407) );
  AOI221_X1 U88615 ( .B1(n120084), .B2(n119001), .C1(n120078), .C2(n118565), 
        .A(n116431), .ZN(n116408) );
  NOR4_X1 U88616 ( .A1(n116425), .A2(n116426), .A3(n116427), .A4(n116428), 
        .ZN(n116409) );
  NAND4_X1 U88617 ( .A1(n116379), .A2(n116380), .A3(n116381), .A4(n116382), 
        .ZN(n5379) );
  AOI221_X1 U88618 ( .B1(n120060), .B2(n119194), .C1(n120054), .C2(n118387), 
        .A(n116405), .ZN(n116379) );
  AOI221_X1 U88619 ( .B1(n120084), .B2(n119002), .C1(n120078), .C2(n118566), 
        .A(n116403), .ZN(n116380) );
  NOR4_X1 U88620 ( .A1(n116397), .A2(n116398), .A3(n116399), .A4(n116400), 
        .ZN(n116381) );
  NAND4_X1 U88621 ( .A1(n116351), .A2(n116352), .A3(n116353), .A4(n116354), 
        .ZN(n5381) );
  AOI221_X1 U88622 ( .B1(n120060), .B2(n119195), .C1(n120054), .C2(n118388), 
        .A(n116377), .ZN(n116351) );
  AOI221_X1 U88623 ( .B1(n120084), .B2(n119003), .C1(n120078), .C2(n118567), 
        .A(n116375), .ZN(n116352) );
  NOR4_X1 U88624 ( .A1(n116369), .A2(n116370), .A3(n116371), .A4(n116372), 
        .ZN(n116353) );
  NAND4_X1 U88625 ( .A1(n117781), .A2(n117782), .A3(n117783), .A4(n117784), 
        .ZN(n5318) );
  AOI221_X1 U88626 ( .B1(n119886), .B2(n118806), .C1(n119880), .C2(n109986), 
        .A(n117801), .ZN(n117782) );
  AOI221_X1 U88627 ( .B1(n119862), .B2(n95436), .C1(n119856), .C2(n118392), 
        .A(n117802), .ZN(n117781) );
  NOR4_X1 U88628 ( .A1(n117797), .A2(n117798), .A3(n117799), .A4(n117800), 
        .ZN(n117783) );
  NAND4_X1 U88629 ( .A1(n117759), .A2(n117760), .A3(n117761), .A4(n117762), 
        .ZN(n5319) );
  AOI221_X1 U88630 ( .B1(n119886), .B2(n118807), .C1(n119880), .C2(n109987), 
        .A(n117779), .ZN(n117760) );
  AOI221_X1 U88631 ( .B1(n119862), .B2(n95437), .C1(n119856), .C2(n118393), 
        .A(n117780), .ZN(n117759) );
  NOR4_X1 U88632 ( .A1(n117775), .A2(n117776), .A3(n117777), .A4(n117778), 
        .ZN(n117761) );
  NAND4_X1 U88633 ( .A1(n117737), .A2(n117738), .A3(n117739), .A4(n117740), 
        .ZN(n5320) );
  AOI221_X1 U88634 ( .B1(n119886), .B2(n118808), .C1(n119880), .C2(n109988), 
        .A(n117757), .ZN(n117738) );
  AOI221_X1 U88635 ( .B1(n119862), .B2(n95438), .C1(n119856), .C2(n118394), 
        .A(n117758), .ZN(n117737) );
  NOR4_X1 U88636 ( .A1(n117753), .A2(n117754), .A3(n117755), .A4(n117756), 
        .ZN(n117739) );
  NAND4_X1 U88637 ( .A1(n117715), .A2(n117716), .A3(n117717), .A4(n117718), 
        .ZN(n5321) );
  AOI221_X1 U88638 ( .B1(n119886), .B2(n118809), .C1(n119880), .C2(n109989), 
        .A(n117735), .ZN(n117716) );
  AOI221_X1 U88639 ( .B1(n119862), .B2(n95439), .C1(n119856), .C2(n118395), 
        .A(n117736), .ZN(n117715) );
  NOR4_X1 U88640 ( .A1(n117731), .A2(n117732), .A3(n117733), .A4(n117734), 
        .ZN(n117717) );
  NAND4_X1 U88641 ( .A1(n117935), .A2(n117936), .A3(n117937), .A4(n117938), 
        .ZN(n5311) );
  AOI221_X1 U88642 ( .B1(n119886), .B2(n118810), .C1(n119880), .C2(n109979), 
        .A(n117969), .ZN(n117936) );
  AOI221_X1 U88643 ( .B1(n119862), .B2(n95429), .C1(n119856), .C2(n118385), 
        .A(n117972), .ZN(n117935) );
  NOR4_X1 U88644 ( .A1(n117963), .A2(n117964), .A3(n117965), .A4(n117966), 
        .ZN(n117937) );
  NAND4_X1 U88645 ( .A1(n117913), .A2(n117914), .A3(n117915), .A4(n117916), 
        .ZN(n5312) );
  AOI221_X1 U88646 ( .B1(n119886), .B2(n118811), .C1(n119880), .C2(n109980), 
        .A(n117933), .ZN(n117914) );
  AOI221_X1 U88647 ( .B1(n119862), .B2(n95430), .C1(n119856), .C2(n118386), 
        .A(n117934), .ZN(n117913) );
  NOR4_X1 U88648 ( .A1(n117929), .A2(n117930), .A3(n117931), .A4(n117932), 
        .ZN(n117915) );
  NAND4_X1 U88649 ( .A1(n117891), .A2(n117892), .A3(n117893), .A4(n117894), 
        .ZN(n5313) );
  AOI221_X1 U88650 ( .B1(n119886), .B2(n118812), .C1(n119880), .C2(n109981), 
        .A(n117911), .ZN(n117892) );
  AOI221_X1 U88651 ( .B1(n119862), .B2(n95431), .C1(n119856), .C2(n118387), 
        .A(n117912), .ZN(n117891) );
  NOR4_X1 U88652 ( .A1(n117907), .A2(n117908), .A3(n117909), .A4(n117910), 
        .ZN(n117893) );
  NAND4_X1 U88653 ( .A1(n117869), .A2(n117870), .A3(n117871), .A4(n117872), 
        .ZN(n5314) );
  AOI221_X1 U88654 ( .B1(n119886), .B2(n118813), .C1(n119880), .C2(n109982), 
        .A(n117889), .ZN(n117870) );
  AOI221_X1 U88655 ( .B1(n119862), .B2(n95432), .C1(n119856), .C2(n118388), 
        .A(n117890), .ZN(n117869) );
  NOR4_X1 U88656 ( .A1(n117885), .A2(n117886), .A3(n117887), .A4(n117888), 
        .ZN(n117871) );
  NAND4_X1 U88657 ( .A1(n117847), .A2(n117848), .A3(n117849), .A4(n117850), 
        .ZN(n5315) );
  AOI221_X1 U88658 ( .B1(n119886), .B2(n118814), .C1(n119880), .C2(n109983), 
        .A(n117867), .ZN(n117848) );
  AOI221_X1 U88659 ( .B1(n119862), .B2(n95433), .C1(n119856), .C2(n118389), 
        .A(n117868), .ZN(n117847) );
  NOR4_X1 U88660 ( .A1(n117863), .A2(n117864), .A3(n117865), .A4(n117866), 
        .ZN(n117849) );
  NAND4_X1 U88661 ( .A1(n117825), .A2(n117826), .A3(n117827), .A4(n117828), 
        .ZN(n5316) );
  AOI221_X1 U88662 ( .B1(n119886), .B2(n118815), .C1(n119880), .C2(n109984), 
        .A(n117845), .ZN(n117826) );
  AOI221_X1 U88663 ( .B1(n119862), .B2(n95434), .C1(n119856), .C2(n118390), 
        .A(n117846), .ZN(n117825) );
  NOR4_X1 U88664 ( .A1(n117841), .A2(n117842), .A3(n117843), .A4(n117844), 
        .ZN(n117827) );
  NAND4_X1 U88665 ( .A1(n117803), .A2(n117804), .A3(n117805), .A4(n117806), 
        .ZN(n5317) );
  AOI221_X1 U88666 ( .B1(n119886), .B2(n118816), .C1(n119880), .C2(n109985), 
        .A(n117823), .ZN(n117804) );
  AOI221_X1 U88667 ( .B1(n119862), .B2(n95435), .C1(n119856), .C2(n118391), 
        .A(n117824), .ZN(n117803) );
  NOR4_X1 U88668 ( .A1(n117819), .A2(n117820), .A3(n117821), .A4(n117822), 
        .ZN(n117805) );
  NAND4_X1 U88669 ( .A1(n116323), .A2(n116324), .A3(n116325), .A4(n116326), 
        .ZN(n5383) );
  AOI221_X1 U88670 ( .B1(n120060), .B2(n119196), .C1(n120054), .C2(n118389), 
        .A(n116349), .ZN(n116323) );
  AOI221_X1 U88671 ( .B1(n120084), .B2(n119004), .C1(n120078), .C2(n118568), 
        .A(n116347), .ZN(n116324) );
  NOR4_X1 U88672 ( .A1(n116341), .A2(n116342), .A3(n116343), .A4(n116344), 
        .ZN(n116325) );
  NAND4_X1 U88673 ( .A1(n116295), .A2(n116296), .A3(n116297), .A4(n116298), 
        .ZN(n5385) );
  AOI221_X1 U88674 ( .B1(n120060), .B2(n119197), .C1(n120054), .C2(n118390), 
        .A(n116321), .ZN(n116295) );
  AOI221_X1 U88675 ( .B1(n120084), .B2(n119005), .C1(n120078), .C2(n118569), 
        .A(n116319), .ZN(n116296) );
  NOR4_X1 U88676 ( .A1(n116313), .A2(n116314), .A3(n116315), .A4(n116316), 
        .ZN(n116297) );
  NAND4_X1 U88677 ( .A1(n116267), .A2(n116268), .A3(n116269), .A4(n116270), 
        .ZN(n5387) );
  AOI221_X1 U88678 ( .B1(n120060), .B2(n119198), .C1(n120054), .C2(n118391), 
        .A(n116293), .ZN(n116267) );
  AOI221_X1 U88679 ( .B1(n120084), .B2(n119006), .C1(n120078), .C2(n118570), 
        .A(n116291), .ZN(n116268) );
  NOR4_X1 U88680 ( .A1(n116285), .A2(n116286), .A3(n116287), .A4(n116288), 
        .ZN(n116269) );
  NAND4_X1 U88681 ( .A1(n116239), .A2(n116240), .A3(n116241), .A4(n116242), 
        .ZN(n5389) );
  AOI221_X1 U88682 ( .B1(n120060), .B2(n119199), .C1(n120054), .C2(n118392), 
        .A(n116265), .ZN(n116239) );
  AOI221_X1 U88683 ( .B1(n120084), .B2(n119007), .C1(n120078), .C2(n118571), 
        .A(n116263), .ZN(n116240) );
  NOR4_X1 U88684 ( .A1(n116257), .A2(n116258), .A3(n116259), .A4(n116260), 
        .ZN(n116241) );
  NAND4_X1 U88685 ( .A1(n116211), .A2(n116212), .A3(n116213), .A4(n116214), 
        .ZN(n5391) );
  AOI221_X1 U88686 ( .B1(n120060), .B2(n119200), .C1(n120054), .C2(n118393), 
        .A(n116237), .ZN(n116211) );
  AOI221_X1 U88687 ( .B1(n120084), .B2(n119008), .C1(n120078), .C2(n118572), 
        .A(n116235), .ZN(n116212) );
  NOR4_X1 U88688 ( .A1(n116229), .A2(n116230), .A3(n116231), .A4(n116232), 
        .ZN(n116213) );
  NAND4_X1 U88689 ( .A1(n116183), .A2(n116184), .A3(n116185), .A4(n116186), 
        .ZN(n5393) );
  AOI221_X1 U88690 ( .B1(n120060), .B2(n119201), .C1(n120054), .C2(n118394), 
        .A(n116209), .ZN(n116183) );
  AOI221_X1 U88691 ( .B1(n120084), .B2(n119009), .C1(n120078), .C2(n118573), 
        .A(n116207), .ZN(n116184) );
  NOR4_X1 U88692 ( .A1(n116201), .A2(n116202), .A3(n116203), .A4(n116204), 
        .ZN(n116185) );
  NAND4_X1 U88693 ( .A1(n116155), .A2(n116156), .A3(n116157), .A4(n116158), 
        .ZN(n5395) );
  AOI221_X1 U88694 ( .B1(n120060), .B2(n119202), .C1(n120054), .C2(n118395), 
        .A(n116181), .ZN(n116155) );
  AOI221_X1 U88695 ( .B1(n120084), .B2(n119010), .C1(n120078), .C2(n118574), 
        .A(n116179), .ZN(n116156) );
  NOR4_X1 U88696 ( .A1(n116173), .A2(n116174), .A3(n116175), .A4(n116176), 
        .ZN(n116157) );
  NAND4_X1 U88697 ( .A1(n116127), .A2(n116128), .A3(n116129), .A4(n116130), 
        .ZN(n5397) );
  AOI221_X1 U88698 ( .B1(n120060), .B2(n119203), .C1(n120054), .C2(n118396), 
        .A(n116153), .ZN(n116127) );
  AOI221_X1 U88699 ( .B1(n120084), .B2(n119011), .C1(n120078), .C2(n118575), 
        .A(n116151), .ZN(n116128) );
  NOR4_X1 U88700 ( .A1(n116145), .A2(n116146), .A3(n116147), .A4(n116148), 
        .ZN(n116129) );
  NAND4_X1 U88701 ( .A1(n116099), .A2(n116100), .A3(n116101), .A4(n116102), 
        .ZN(n5399) );
  AOI221_X1 U88702 ( .B1(n120061), .B2(n119204), .C1(n120055), .C2(n118397), 
        .A(n116125), .ZN(n116099) );
  AOI221_X1 U88703 ( .B1(n120085), .B2(n119012), .C1(n120079), .C2(n118576), 
        .A(n116123), .ZN(n116100) );
  NOR4_X1 U88704 ( .A1(n116117), .A2(n116118), .A3(n116119), .A4(n116120), 
        .ZN(n116101) );
  NAND4_X1 U88705 ( .A1(n116071), .A2(n116072), .A3(n116073), .A4(n116074), 
        .ZN(n5401) );
  AOI221_X1 U88706 ( .B1(n120061), .B2(n119205), .C1(n120055), .C2(n118398), 
        .A(n116097), .ZN(n116071) );
  AOI221_X1 U88707 ( .B1(n120085), .B2(n119013), .C1(n120079), .C2(n118577), 
        .A(n116095), .ZN(n116072) );
  NOR4_X1 U88708 ( .A1(n116089), .A2(n116090), .A3(n116091), .A4(n116092), 
        .ZN(n116073) );
  NAND4_X1 U88709 ( .A1(n116043), .A2(n116044), .A3(n116045), .A4(n116046), 
        .ZN(n5403) );
  AOI221_X1 U88710 ( .B1(n120061), .B2(n119206), .C1(n120055), .C2(n118399), 
        .A(n116069), .ZN(n116043) );
  AOI221_X1 U88711 ( .B1(n120085), .B2(n119014), .C1(n120079), .C2(n118578), 
        .A(n116067), .ZN(n116044) );
  NOR4_X1 U88712 ( .A1(n116061), .A2(n116062), .A3(n116063), .A4(n116064), 
        .ZN(n116045) );
  NAND4_X1 U88713 ( .A1(n116015), .A2(n116016), .A3(n116017), .A4(n116018), 
        .ZN(n5405) );
  AOI221_X1 U88714 ( .B1(n120061), .B2(n119207), .C1(n120055), .C2(n118400), 
        .A(n116041), .ZN(n116015) );
  AOI221_X1 U88715 ( .B1(n120085), .B2(n119015), .C1(n120079), .C2(n118579), 
        .A(n116039), .ZN(n116016) );
  NOR4_X1 U88716 ( .A1(n116033), .A2(n116034), .A3(n116035), .A4(n116036), 
        .ZN(n116017) );
  NAND4_X1 U88717 ( .A1(n115987), .A2(n115988), .A3(n115989), .A4(n115990), 
        .ZN(n5407) );
  AOI221_X1 U88718 ( .B1(n120061), .B2(n119208), .C1(n120055), .C2(n118401), 
        .A(n116013), .ZN(n115987) );
  AOI221_X1 U88719 ( .B1(n120085), .B2(n119016), .C1(n120079), .C2(n118580), 
        .A(n116011), .ZN(n115988) );
  NOR4_X1 U88720 ( .A1(n116005), .A2(n116006), .A3(n116007), .A4(n116008), 
        .ZN(n115989) );
  NAND4_X1 U88721 ( .A1(n115959), .A2(n115960), .A3(n115961), .A4(n115962), 
        .ZN(n5409) );
  AOI221_X1 U88722 ( .B1(n120061), .B2(n119209), .C1(n120055), .C2(n118402), 
        .A(n115985), .ZN(n115959) );
  AOI221_X1 U88723 ( .B1(n120085), .B2(n119017), .C1(n120079), .C2(n118581), 
        .A(n115983), .ZN(n115960) );
  NOR4_X1 U88724 ( .A1(n115977), .A2(n115978), .A3(n115979), .A4(n115980), 
        .ZN(n115961) );
  NAND4_X1 U88725 ( .A1(n115931), .A2(n115932), .A3(n115933), .A4(n115934), 
        .ZN(n5411) );
  AOI221_X1 U88726 ( .B1(n120061), .B2(n119210), .C1(n120055), .C2(n118403), 
        .A(n115957), .ZN(n115931) );
  AOI221_X1 U88727 ( .B1(n120085), .B2(n119018), .C1(n120079), .C2(n118582), 
        .A(n115955), .ZN(n115932) );
  NOR4_X1 U88728 ( .A1(n115949), .A2(n115950), .A3(n115951), .A4(n115952), 
        .ZN(n115933) );
  NAND4_X1 U88729 ( .A1(n115903), .A2(n115904), .A3(n115905), .A4(n115906), 
        .ZN(n5413) );
  AOI221_X1 U88730 ( .B1(n120061), .B2(n119211), .C1(n120055), .C2(n118404), 
        .A(n115929), .ZN(n115903) );
  AOI221_X1 U88731 ( .B1(n120085), .B2(n119019), .C1(n120079), .C2(n118583), 
        .A(n115927), .ZN(n115904) );
  NOR4_X1 U88732 ( .A1(n115921), .A2(n115922), .A3(n115923), .A4(n115924), 
        .ZN(n115905) );
  NAND4_X1 U88733 ( .A1(n115875), .A2(n115876), .A3(n115877), .A4(n115878), 
        .ZN(n5415) );
  AOI221_X1 U88734 ( .B1(n120061), .B2(n119212), .C1(n120055), .C2(n118405), 
        .A(n115901), .ZN(n115875) );
  AOI221_X1 U88735 ( .B1(n120085), .B2(n119020), .C1(n120079), .C2(n118584), 
        .A(n115899), .ZN(n115876) );
  NOR4_X1 U88736 ( .A1(n115893), .A2(n115894), .A3(n115895), .A4(n115896), 
        .ZN(n115877) );
  NAND4_X1 U88737 ( .A1(n115847), .A2(n115848), .A3(n115849), .A4(n115850), 
        .ZN(n5417) );
  AOI221_X1 U88738 ( .B1(n120061), .B2(n119213), .C1(n120055), .C2(n118406), 
        .A(n115873), .ZN(n115847) );
  AOI221_X1 U88739 ( .B1(n120085), .B2(n119021), .C1(n120079), .C2(n118585), 
        .A(n115871), .ZN(n115848) );
  NOR4_X1 U88740 ( .A1(n115865), .A2(n115866), .A3(n115867), .A4(n115868), 
        .ZN(n115849) );
  NAND4_X1 U88741 ( .A1(n115819), .A2(n115820), .A3(n115821), .A4(n115822), 
        .ZN(n5419) );
  AOI221_X1 U88742 ( .B1(n120061), .B2(n119214), .C1(n120055), .C2(n118407), 
        .A(n115845), .ZN(n115819) );
  AOI221_X1 U88743 ( .B1(n120085), .B2(n119022), .C1(n120079), .C2(n118586), 
        .A(n115843), .ZN(n115820) );
  NOR4_X1 U88744 ( .A1(n115837), .A2(n115838), .A3(n115839), .A4(n115840), 
        .ZN(n115821) );
  NAND4_X1 U88745 ( .A1(n115791), .A2(n115792), .A3(n115793), .A4(n115794), 
        .ZN(n5421) );
  AOI221_X1 U88746 ( .B1(n120061), .B2(n119215), .C1(n120055), .C2(n118408), 
        .A(n115817), .ZN(n115791) );
  AOI221_X1 U88747 ( .B1(n120085), .B2(n119023), .C1(n120079), .C2(n118587), 
        .A(n115815), .ZN(n115792) );
  NOR4_X1 U88748 ( .A1(n115809), .A2(n115810), .A3(n115811), .A4(n115812), 
        .ZN(n115793) );
  NAND4_X1 U88749 ( .A1(n115763), .A2(n115764), .A3(n115765), .A4(n115766), 
        .ZN(n5423) );
  AOI221_X1 U88750 ( .B1(n120062), .B2(n119216), .C1(n120056), .C2(n118409), 
        .A(n115789), .ZN(n115763) );
  AOI221_X1 U88751 ( .B1(n120086), .B2(n119024), .C1(n120080), .C2(n118588), 
        .A(n115787), .ZN(n115764) );
  NOR4_X1 U88752 ( .A1(n115781), .A2(n115782), .A3(n115783), .A4(n115784), 
        .ZN(n115765) );
  NAND4_X1 U88753 ( .A1(n115735), .A2(n115736), .A3(n115737), .A4(n115738), 
        .ZN(n5425) );
  AOI221_X1 U88754 ( .B1(n120062), .B2(n119217), .C1(n120056), .C2(n118410), 
        .A(n115761), .ZN(n115735) );
  AOI221_X1 U88755 ( .B1(n120086), .B2(n119025), .C1(n120080), .C2(n118589), 
        .A(n115759), .ZN(n115736) );
  NOR4_X1 U88756 ( .A1(n115753), .A2(n115754), .A3(n115755), .A4(n115756), 
        .ZN(n115737) );
  NAND4_X1 U88757 ( .A1(n115707), .A2(n115708), .A3(n115709), .A4(n115710), 
        .ZN(n5427) );
  AOI221_X1 U88758 ( .B1(n120062), .B2(n119218), .C1(n120056), .C2(n118411), 
        .A(n115733), .ZN(n115707) );
  AOI221_X1 U88759 ( .B1(n120086), .B2(n119026), .C1(n120080), .C2(n118590), 
        .A(n115731), .ZN(n115708) );
  NOR4_X1 U88760 ( .A1(n115725), .A2(n115726), .A3(n115727), .A4(n115728), 
        .ZN(n115709) );
  NAND4_X1 U88761 ( .A1(n115679), .A2(n115680), .A3(n115681), .A4(n115682), 
        .ZN(n5429) );
  AOI221_X1 U88762 ( .B1(n120062), .B2(n119219), .C1(n120056), .C2(n118412), 
        .A(n115705), .ZN(n115679) );
  AOI221_X1 U88763 ( .B1(n120086), .B2(n119027), .C1(n120080), .C2(n118591), 
        .A(n115703), .ZN(n115680) );
  NOR4_X1 U88764 ( .A1(n115697), .A2(n115698), .A3(n115699), .A4(n115700), 
        .ZN(n115681) );
  NAND4_X1 U88765 ( .A1(n115651), .A2(n115652), .A3(n115653), .A4(n115654), 
        .ZN(n5431) );
  AOI221_X1 U88766 ( .B1(n120062), .B2(n119220), .C1(n120056), .C2(n118413), 
        .A(n115677), .ZN(n115651) );
  AOI221_X1 U88767 ( .B1(n120086), .B2(n119028), .C1(n120080), .C2(n118592), 
        .A(n115675), .ZN(n115652) );
  NOR4_X1 U88768 ( .A1(n115669), .A2(n115670), .A3(n115671), .A4(n115672), 
        .ZN(n115653) );
  NAND4_X1 U88769 ( .A1(n115623), .A2(n115624), .A3(n115625), .A4(n115626), 
        .ZN(n5433) );
  AOI221_X1 U88770 ( .B1(n120062), .B2(n119221), .C1(n120056), .C2(n118414), 
        .A(n115649), .ZN(n115623) );
  AOI221_X1 U88771 ( .B1(n120086), .B2(n119029), .C1(n120080), .C2(n118593), 
        .A(n115647), .ZN(n115624) );
  NOR4_X1 U88772 ( .A1(n115641), .A2(n115642), .A3(n115643), .A4(n115644), 
        .ZN(n115625) );
  NAND4_X1 U88773 ( .A1(n115595), .A2(n115596), .A3(n115597), .A4(n115598), 
        .ZN(n5435) );
  AOI221_X1 U88774 ( .B1(n120062), .B2(n119222), .C1(n120056), .C2(n118415), 
        .A(n115621), .ZN(n115595) );
  AOI221_X1 U88775 ( .B1(n120086), .B2(n119030), .C1(n120080), .C2(n118594), 
        .A(n115619), .ZN(n115596) );
  NOR4_X1 U88776 ( .A1(n115613), .A2(n115614), .A3(n115615), .A4(n115616), 
        .ZN(n115597) );
  NAND4_X1 U88777 ( .A1(n115567), .A2(n115568), .A3(n115569), .A4(n115570), 
        .ZN(n5437) );
  AOI221_X1 U88778 ( .B1(n120062), .B2(n119223), .C1(n120056), .C2(n118416), 
        .A(n115593), .ZN(n115567) );
  AOI221_X1 U88779 ( .B1(n120086), .B2(n119031), .C1(n120080), .C2(n118595), 
        .A(n115591), .ZN(n115568) );
  NOR4_X1 U88780 ( .A1(n115585), .A2(n115586), .A3(n115587), .A4(n115588), 
        .ZN(n115569) );
  NAND4_X1 U88781 ( .A1(n115539), .A2(n115540), .A3(n115541), .A4(n115542), 
        .ZN(n5439) );
  AOI221_X1 U88782 ( .B1(n120062), .B2(n119224), .C1(n120056), .C2(n118417), 
        .A(n115565), .ZN(n115539) );
  AOI221_X1 U88783 ( .B1(n120086), .B2(n119032), .C1(n120080), .C2(n118596), 
        .A(n115563), .ZN(n115540) );
  NOR4_X1 U88784 ( .A1(n115557), .A2(n115558), .A3(n115559), .A4(n115560), 
        .ZN(n115541) );
  NAND4_X1 U88785 ( .A1(n115511), .A2(n115512), .A3(n115513), .A4(n115514), 
        .ZN(n5441) );
  AOI221_X1 U88786 ( .B1(n120062), .B2(n119225), .C1(n120056), .C2(n118418), 
        .A(n115537), .ZN(n115511) );
  AOI221_X1 U88787 ( .B1(n120086), .B2(n119033), .C1(n120080), .C2(n118597), 
        .A(n115535), .ZN(n115512) );
  NOR4_X1 U88788 ( .A1(n115529), .A2(n115530), .A3(n115531), .A4(n115532), 
        .ZN(n115513) );
  NAND4_X1 U88789 ( .A1(n115483), .A2(n115484), .A3(n115485), .A4(n115486), 
        .ZN(n5443) );
  AOI221_X1 U88790 ( .B1(n120062), .B2(n119226), .C1(n120056), .C2(n118419), 
        .A(n115509), .ZN(n115483) );
  AOI221_X1 U88791 ( .B1(n120086), .B2(n119034), .C1(n120080), .C2(n118598), 
        .A(n115507), .ZN(n115484) );
  NOR4_X1 U88792 ( .A1(n115501), .A2(n115502), .A3(n115503), .A4(n115504), 
        .ZN(n115485) );
  NAND4_X1 U88793 ( .A1(n115455), .A2(n115456), .A3(n115457), .A4(n115458), 
        .ZN(n5445) );
  AOI221_X1 U88794 ( .B1(n120062), .B2(n119227), .C1(n120056), .C2(n118420), 
        .A(n115481), .ZN(n115455) );
  AOI221_X1 U88795 ( .B1(n120086), .B2(n119035), .C1(n120080), .C2(n118599), 
        .A(n115479), .ZN(n115456) );
  NOR4_X1 U88796 ( .A1(n115473), .A2(n115474), .A3(n115475), .A4(n115476), 
        .ZN(n115457) );
  NAND4_X1 U88797 ( .A1(n115427), .A2(n115428), .A3(n115429), .A4(n115430), 
        .ZN(n5447) );
  AOI221_X1 U88798 ( .B1(n120063), .B2(n119228), .C1(n120057), .C2(n118421), 
        .A(n115453), .ZN(n115427) );
  AOI221_X1 U88799 ( .B1(n120087), .B2(n119036), .C1(n120081), .C2(n118600), 
        .A(n115451), .ZN(n115428) );
  NOR4_X1 U88800 ( .A1(n115445), .A2(n115446), .A3(n115447), .A4(n115448), 
        .ZN(n115429) );
  NAND4_X1 U88801 ( .A1(n115399), .A2(n115400), .A3(n115401), .A4(n115402), 
        .ZN(n5449) );
  AOI221_X1 U88802 ( .B1(n120063), .B2(n119229), .C1(n120057), .C2(n118422), 
        .A(n115425), .ZN(n115399) );
  AOI221_X1 U88803 ( .B1(n120087), .B2(n119037), .C1(n120081), .C2(n118601), 
        .A(n115423), .ZN(n115400) );
  NOR4_X1 U88804 ( .A1(n115417), .A2(n115418), .A3(n115419), .A4(n115420), 
        .ZN(n115401) );
  NAND4_X1 U88805 ( .A1(n115371), .A2(n115372), .A3(n115373), .A4(n115374), 
        .ZN(n5451) );
  AOI221_X1 U88806 ( .B1(n120063), .B2(n119230), .C1(n120057), .C2(n118423), 
        .A(n115397), .ZN(n115371) );
  AOI221_X1 U88807 ( .B1(n120087), .B2(n119038), .C1(n120081), .C2(n118602), 
        .A(n115395), .ZN(n115372) );
  NOR4_X1 U88808 ( .A1(n115389), .A2(n115390), .A3(n115391), .A4(n115392), 
        .ZN(n115373) );
  NAND4_X1 U88809 ( .A1(n115343), .A2(n115344), .A3(n115345), .A4(n115346), 
        .ZN(n5453) );
  AOI221_X1 U88810 ( .B1(n120063), .B2(n119231), .C1(n120057), .C2(n118424), 
        .A(n115369), .ZN(n115343) );
  AOI221_X1 U88811 ( .B1(n120087), .B2(n119039), .C1(n120081), .C2(n118603), 
        .A(n115367), .ZN(n115344) );
  NOR4_X1 U88812 ( .A1(n115361), .A2(n115362), .A3(n115363), .A4(n115364), 
        .ZN(n115345) );
  NAND4_X1 U88813 ( .A1(n115315), .A2(n115316), .A3(n115317), .A4(n115318), 
        .ZN(n5455) );
  AOI221_X1 U88814 ( .B1(n120063), .B2(n119232), .C1(n120057), .C2(n118425), 
        .A(n115341), .ZN(n115315) );
  AOI221_X1 U88815 ( .B1(n120087), .B2(n119040), .C1(n120081), .C2(n118604), 
        .A(n115339), .ZN(n115316) );
  NOR4_X1 U88816 ( .A1(n115333), .A2(n115334), .A3(n115335), .A4(n115336), 
        .ZN(n115317) );
  NAND4_X1 U88817 ( .A1(n115287), .A2(n115288), .A3(n115289), .A4(n115290), 
        .ZN(n5457) );
  AOI221_X1 U88818 ( .B1(n120063), .B2(n119233), .C1(n120057), .C2(n118426), 
        .A(n115313), .ZN(n115287) );
  AOI221_X1 U88819 ( .B1(n120087), .B2(n119041), .C1(n120081), .C2(n118605), 
        .A(n115311), .ZN(n115288) );
  NOR4_X1 U88820 ( .A1(n115305), .A2(n115306), .A3(n115307), .A4(n115308), 
        .ZN(n115289) );
  NAND4_X1 U88821 ( .A1(n115259), .A2(n115260), .A3(n115261), .A4(n115262), 
        .ZN(n5459) );
  AOI221_X1 U88822 ( .B1(n120063), .B2(n119234), .C1(n120057), .C2(n118427), 
        .A(n115285), .ZN(n115259) );
  AOI221_X1 U88823 ( .B1(n120087), .B2(n119042), .C1(n120081), .C2(n118606), 
        .A(n115283), .ZN(n115260) );
  NOR4_X1 U88824 ( .A1(n115277), .A2(n115278), .A3(n115279), .A4(n115280), 
        .ZN(n115261) );
  NAND4_X1 U88825 ( .A1(n115231), .A2(n115232), .A3(n115233), .A4(n115234), 
        .ZN(n5461) );
  AOI221_X1 U88826 ( .B1(n120063), .B2(n119235), .C1(n120057), .C2(n118428), 
        .A(n115257), .ZN(n115231) );
  AOI221_X1 U88827 ( .B1(n120087), .B2(n119043), .C1(n120081), .C2(n118607), 
        .A(n115255), .ZN(n115232) );
  NOR4_X1 U88828 ( .A1(n115249), .A2(n115250), .A3(n115251), .A4(n115252), 
        .ZN(n115233) );
  NAND4_X1 U88829 ( .A1(n115203), .A2(n115204), .A3(n115205), .A4(n115206), 
        .ZN(n5463) );
  AOI221_X1 U88830 ( .B1(n120063), .B2(n119236), .C1(n120057), .C2(n118429), 
        .A(n115229), .ZN(n115203) );
  AOI221_X1 U88831 ( .B1(n120087), .B2(n119044), .C1(n120081), .C2(n118608), 
        .A(n115227), .ZN(n115204) );
  NOR4_X1 U88832 ( .A1(n115221), .A2(n115222), .A3(n115223), .A4(n115224), 
        .ZN(n115205) );
  NAND4_X1 U88833 ( .A1(n115175), .A2(n115176), .A3(n115177), .A4(n115178), 
        .ZN(n5465) );
  AOI221_X1 U88834 ( .B1(n120063), .B2(n119237), .C1(n120057), .C2(n118430), 
        .A(n115201), .ZN(n115175) );
  AOI221_X1 U88835 ( .B1(n120087), .B2(n119045), .C1(n120081), .C2(n118609), 
        .A(n115199), .ZN(n115176) );
  NOR4_X1 U88836 ( .A1(n115193), .A2(n115194), .A3(n115195), .A4(n115196), 
        .ZN(n115177) );
  AND3_X1 U88837 ( .A1(WR), .A2(ENABLE), .A3(ADD_WR[4]), .ZN(n114302) );
  INV_X1 U88838 ( .A(RESET), .ZN(n113892) );
  INV_X1 U88839 ( .A(DATAIN[60]), .ZN(n113771) );
  INV_X1 U88840 ( .A(DATAIN[61]), .ZN(n113770) );
  INV_X1 U88841 ( .A(DATAIN[62]), .ZN(n113769) );
  INV_X1 U88842 ( .A(DATAIN[63]), .ZN(n113768) );
  INV_X1 U88843 ( .A(DATAIN[0]), .ZN(n113891) );
  INV_X1 U88844 ( .A(DATAIN[1]), .ZN(n113889) );
  INV_X1 U88845 ( .A(DATAIN[2]), .ZN(n113887) );
  INV_X1 U88846 ( .A(DATAIN[3]), .ZN(n113885) );
  INV_X1 U88847 ( .A(DATAIN[4]), .ZN(n113883) );
  INV_X1 U88848 ( .A(DATAIN[5]), .ZN(n113881) );
  INV_X1 U88849 ( .A(DATAIN[6]), .ZN(n113879) );
  INV_X1 U88850 ( .A(DATAIN[7]), .ZN(n113877) );
  INV_X1 U88851 ( .A(DATAIN[8]), .ZN(n113875) );
  INV_X1 U88852 ( .A(DATAIN[9]), .ZN(n113873) );
  INV_X1 U88853 ( .A(DATAIN[10]), .ZN(n113871) );
  INV_X1 U88854 ( .A(DATAIN[11]), .ZN(n113869) );
  INV_X1 U88855 ( .A(DATAIN[12]), .ZN(n113867) );
  INV_X1 U88856 ( .A(DATAIN[13]), .ZN(n113865) );
  INV_X1 U88857 ( .A(DATAIN[14]), .ZN(n113863) );
  INV_X1 U88858 ( .A(DATAIN[15]), .ZN(n113861) );
  INV_X1 U88859 ( .A(DATAIN[16]), .ZN(n113859) );
  INV_X1 U88860 ( .A(DATAIN[17]), .ZN(n113857) );
  INV_X1 U88861 ( .A(DATAIN[18]), .ZN(n113855) );
  INV_X1 U88862 ( .A(DATAIN[19]), .ZN(n113853) );
  INV_X1 U88863 ( .A(DATAIN[20]), .ZN(n113851) );
  INV_X1 U88864 ( .A(DATAIN[21]), .ZN(n113849) );
  INV_X1 U88865 ( .A(DATAIN[22]), .ZN(n113847) );
  INV_X1 U88866 ( .A(DATAIN[23]), .ZN(n113845) );
  INV_X1 U88867 ( .A(DATAIN[24]), .ZN(n113843) );
  INV_X1 U88868 ( .A(DATAIN[25]), .ZN(n113841) );
  INV_X1 U88869 ( .A(DATAIN[26]), .ZN(n113839) );
  INV_X1 U88870 ( .A(DATAIN[27]), .ZN(n113837) );
  INV_X1 U88871 ( .A(DATAIN[28]), .ZN(n113835) );
  INV_X1 U88872 ( .A(DATAIN[29]), .ZN(n113833) );
  INV_X1 U88873 ( .A(DATAIN[30]), .ZN(n113831) );
  INV_X1 U88874 ( .A(DATAIN[31]), .ZN(n113829) );
  INV_X1 U88875 ( .A(DATAIN[32]), .ZN(n113827) );
  INV_X1 U88876 ( .A(DATAIN[33]), .ZN(n113825) );
  INV_X1 U88877 ( .A(DATAIN[34]), .ZN(n113823) );
  INV_X1 U88878 ( .A(DATAIN[35]), .ZN(n113821) );
  INV_X1 U88879 ( .A(DATAIN[36]), .ZN(n113819) );
  INV_X1 U88880 ( .A(DATAIN[37]), .ZN(n113817) );
  INV_X1 U88881 ( .A(DATAIN[38]), .ZN(n113815) );
  INV_X1 U88882 ( .A(DATAIN[39]), .ZN(n113813) );
  INV_X1 U88883 ( .A(DATAIN[40]), .ZN(n113811) );
  INV_X1 U88884 ( .A(DATAIN[41]), .ZN(n113809) );
  INV_X1 U88885 ( .A(DATAIN[42]), .ZN(n113807) );
  INV_X1 U88886 ( .A(DATAIN[43]), .ZN(n113805) );
  INV_X1 U88887 ( .A(DATAIN[44]), .ZN(n113803) );
  INV_X1 U88888 ( .A(DATAIN[45]), .ZN(n113801) );
  INV_X1 U88889 ( .A(DATAIN[46]), .ZN(n113799) );
  INV_X1 U88890 ( .A(DATAIN[47]), .ZN(n113797) );
  INV_X1 U88891 ( .A(DATAIN[48]), .ZN(n113795) );
  INV_X1 U88892 ( .A(DATAIN[49]), .ZN(n113793) );
  INV_X1 U88893 ( .A(DATAIN[50]), .ZN(n113791) );
  INV_X1 U88894 ( .A(DATAIN[51]), .ZN(n113789) );
  INV_X1 U88895 ( .A(DATAIN[52]), .ZN(n113787) );
  INV_X1 U88896 ( .A(DATAIN[53]), .ZN(n113785) );
  INV_X1 U88897 ( .A(DATAIN[54]), .ZN(n113783) );
  INV_X1 U88898 ( .A(DATAIN[55]), .ZN(n113781) );
  INV_X1 U88899 ( .A(DATAIN[56]), .ZN(n113779) );
  INV_X1 U88900 ( .A(DATAIN[57]), .ZN(n113777) );
  INV_X1 U88901 ( .A(DATAIN[58]), .ZN(n113775) );
  INV_X1 U88902 ( .A(DATAIN[59]), .ZN(n113773) );
  INV_X1 U88903 ( .A(ADD_WR[3]), .ZN(n113988) );
  INV_X1 U88904 ( .A(ADD_WR[0]), .ZN(n113987) );
  INV_X1 U88905 ( .A(ADD_WR[1]), .ZN(n114376) );
  INV_X1 U88906 ( .A(ADD_RD2[1]), .ZN(n117973) );
  INV_X1 U88907 ( .A(ADD_RD1[2]), .ZN(n116475) );
  INV_X1 U88908 ( .A(ADD_RD2[2]), .ZN(n117971) );
  INV_X1 U88909 ( .A(ADD_RD1[1]), .ZN(n116478) );
  INV_X1 U88910 ( .A(ADD_WR[2]), .ZN(n114375) );
  AND3_X1 U88911 ( .A1(ENABLE), .A2(n114138), .A3(WR), .ZN(n113989) );
  INV_X1 U88912 ( .A(ADD_WR[4]), .ZN(n114138) );
  CLKBUF_X1 U88913 ( .A(n116532), .Z(n119849) );
  CLKBUF_X1 U88914 ( .A(n116531), .Z(n119855) );
  CLKBUF_X1 U88915 ( .A(n116529), .Z(n119861) );
  CLKBUF_X1 U88916 ( .A(n116528), .Z(n119867) );
  CLKBUF_X1 U88917 ( .A(n116527), .Z(n119873) );
  CLKBUF_X1 U88918 ( .A(n116526), .Z(n119879) );
  CLKBUF_X1 U88919 ( .A(n116523), .Z(n119885) );
  CLKBUF_X1 U88920 ( .A(n116522), .Z(n119891) );
  CLKBUF_X1 U88921 ( .A(n116521), .Z(n119897) );
  CLKBUF_X1 U88922 ( .A(n116520), .Z(n119903) );
  CLKBUF_X1 U88923 ( .A(n116519), .Z(n119909) );
  CLKBUF_X1 U88924 ( .A(n116518), .Z(n119915) );
  CLKBUF_X1 U88925 ( .A(n116517), .Z(n119921) );
  CLKBUF_X1 U88926 ( .A(n116516), .Z(n119927) );
  CLKBUF_X1 U88927 ( .A(n116515), .Z(n119933) );
  CLKBUF_X1 U88928 ( .A(n116514), .Z(n119939) );
  CLKBUF_X1 U88929 ( .A(n116513), .Z(n119945) );
  CLKBUF_X1 U88930 ( .A(n116508), .Z(n119951) );
  CLKBUF_X1 U88931 ( .A(n116507), .Z(n119957) );
  CLKBUF_X1 U88932 ( .A(n116505), .Z(n119963) );
  CLKBUF_X1 U88933 ( .A(n116504), .Z(n119969) );
  CLKBUF_X1 U88934 ( .A(n116503), .Z(n119975) );
  CLKBUF_X1 U88935 ( .A(n116502), .Z(n119981) );
  CLKBUF_X1 U88936 ( .A(n116500), .Z(n119987) );
  CLKBUF_X1 U88937 ( .A(n116499), .Z(n119993) );
  CLKBUF_X1 U88938 ( .A(n116497), .Z(n119999) );
  CLKBUF_X1 U88939 ( .A(n116495), .Z(n120005) );
  CLKBUF_X1 U88940 ( .A(n116493), .Z(n120011) );
  CLKBUF_X1 U88941 ( .A(n116492), .Z(n120017) );
  CLKBUF_X1 U88942 ( .A(n116491), .Z(n120023) );
  CLKBUF_X1 U88943 ( .A(n116490), .Z(n120029) );
  CLKBUF_X1 U88944 ( .A(n116488), .Z(n120035) );
  CLKBUF_X1 U88945 ( .A(n116487), .Z(n120041) );
  CLKBUF_X1 U88946 ( .A(n114703), .Z(n120047) );
  CLKBUF_X1 U88947 ( .A(n114702), .Z(n120053) );
  CLKBUF_X1 U88948 ( .A(n114700), .Z(n120059) );
  CLKBUF_X1 U88949 ( .A(n114698), .Z(n120065) );
  CLKBUF_X1 U88950 ( .A(n114697), .Z(n120071) );
  CLKBUF_X1 U88951 ( .A(n114696), .Z(n120077) );
  CLKBUF_X1 U88952 ( .A(n114693), .Z(n120083) );
  CLKBUF_X1 U88953 ( .A(n114691), .Z(n120089) );
  CLKBUF_X1 U88954 ( .A(n114690), .Z(n120095) );
  CLKBUF_X1 U88955 ( .A(n114689), .Z(n120101) );
  CLKBUF_X1 U88956 ( .A(n114688), .Z(n120107) );
  CLKBUF_X1 U88957 ( .A(n114687), .Z(n120113) );
  CLKBUF_X1 U88958 ( .A(n114686), .Z(n120119) );
  CLKBUF_X1 U88959 ( .A(n114685), .Z(n120125) );
  CLKBUF_X1 U88960 ( .A(n114684), .Z(n120131) );
  CLKBUF_X1 U88961 ( .A(n114683), .Z(n120137) );
  CLKBUF_X1 U88962 ( .A(n114682), .Z(n120143) );
  CLKBUF_X1 U88963 ( .A(n114676), .Z(n120149) );
  CLKBUF_X1 U88964 ( .A(n114675), .Z(n120155) );
  CLKBUF_X1 U88965 ( .A(n114673), .Z(n120161) );
  CLKBUF_X1 U88966 ( .A(n114672), .Z(n120167) );
  CLKBUF_X1 U88967 ( .A(n114670), .Z(n120173) );
  CLKBUF_X1 U88968 ( .A(n114669), .Z(n120179) );
  CLKBUF_X1 U88969 ( .A(n114667), .Z(n120185) );
  CLKBUF_X1 U88970 ( .A(n114666), .Z(n120191) );
  CLKBUF_X1 U88971 ( .A(n114664), .Z(n120197) );
  CLKBUF_X1 U88972 ( .A(n114662), .Z(n120203) );
  CLKBUF_X1 U88973 ( .A(n114660), .Z(n120209) );
  CLKBUF_X1 U88974 ( .A(n114659), .Z(n120215) );
  CLKBUF_X1 U88975 ( .A(n114658), .Z(n120221) );
  CLKBUF_X1 U88976 ( .A(n114657), .Z(n120227) );
  CLKBUF_X1 U88977 ( .A(n114655), .Z(n120233) );
  CLKBUF_X1 U88978 ( .A(n114654), .Z(n120239) );
  CLKBUF_X1 U88979 ( .A(n114645), .Z(n120245) );
  CLKBUF_X1 U88980 ( .A(n114579), .Z(n120258) );
  CLKBUF_X1 U88981 ( .A(n114576), .Z(n120271) );
  CLKBUF_X1 U88982 ( .A(n114575), .Z(n120277) );
  CLKBUF_X1 U88983 ( .A(n114511), .Z(n120283) );
  CLKBUF_X1 U88984 ( .A(n114445), .Z(n120296) );
  CLKBUF_X1 U88985 ( .A(n114379), .Z(n120309) );
  CLKBUF_X1 U88986 ( .A(n114373), .Z(n120322) );
  CLKBUF_X1 U88987 ( .A(n114372), .Z(n120328) );
  CLKBUF_X1 U88988 ( .A(n114307), .Z(n120334) );
  CLKBUF_X1 U88989 ( .A(n114304), .Z(n120347) );
  CLKBUF_X1 U88990 ( .A(n114303), .Z(n120353) );
  CLKBUF_X1 U88991 ( .A(n114301), .Z(n120359) );
  CLKBUF_X1 U88992 ( .A(n114300), .Z(n120365) );
  CLKBUF_X1 U88993 ( .A(n114236), .Z(n120371) );
  CLKBUF_X1 U88994 ( .A(n114214), .Z(n120384) );
  CLKBUF_X1 U88995 ( .A(n114213), .Z(n120390) );
  CLKBUF_X1 U88996 ( .A(n114212), .Z(n120396) );
  CLKBUF_X1 U88997 ( .A(n114211), .Z(n120402) );
  CLKBUF_X1 U88998 ( .A(n114147), .Z(n120408) );
  CLKBUF_X1 U88999 ( .A(n114143), .Z(n120421) );
  CLKBUF_X1 U89000 ( .A(n114142), .Z(n120427) );
  CLKBUF_X1 U89001 ( .A(n114140), .Z(n120433) );
  CLKBUF_X1 U89002 ( .A(n114139), .Z(n120439) );
  CLKBUF_X1 U89003 ( .A(n114137), .Z(n120445) );
  CLKBUF_X1 U89004 ( .A(n114136), .Z(n120451) );
  CLKBUF_X1 U89005 ( .A(n114135), .Z(n120457) );
  CLKBUF_X1 U89006 ( .A(n114134), .Z(n120463) );
  CLKBUF_X1 U89007 ( .A(n114133), .Z(n120469) );
  CLKBUF_X1 U89008 ( .A(n114132), .Z(n120475) );
  CLKBUF_X1 U89009 ( .A(n114131), .Z(n120481) );
  CLKBUF_X1 U89010 ( .A(n114130), .Z(n120487) );
  CLKBUF_X1 U89011 ( .A(n114129), .Z(n120493) );
  CLKBUF_X1 U89012 ( .A(n114128), .Z(n120499) );
  CLKBUF_X1 U89013 ( .A(n114124), .Z(n120505) );
  CLKBUF_X1 U89014 ( .A(n114122), .Z(n120511) );
  CLKBUF_X1 U89015 ( .A(n114057), .Z(n120517) );
  CLKBUF_X1 U89016 ( .A(n114053), .Z(n120530) );
  CLKBUF_X1 U89017 ( .A(n114052), .Z(n120536) );
  CLKBUF_X1 U89018 ( .A(n113991), .Z(n120542) );
  CLKBUF_X1 U89019 ( .A(n113982), .Z(n120555) );
  CLKBUF_X1 U89020 ( .A(n113980), .Z(n120561) );
  CLKBUF_X1 U89021 ( .A(n113916), .Z(n120567) );
  CLKBUF_X1 U89022 ( .A(n113912), .Z(n120580) );
  CLKBUF_X1 U89023 ( .A(n113911), .Z(n120586) );
  CLKBUF_X1 U89024 ( .A(n113910), .Z(n120592) );
  CLKBUF_X1 U89025 ( .A(n113909), .Z(n120598) );
  CLKBUF_X1 U89026 ( .A(n113904), .Z(n120604) );
  CLKBUF_X1 U89027 ( .A(n113902), .Z(n120610) );
  CLKBUF_X1 U89028 ( .A(n113897), .Z(n120616) );
  CLKBUF_X1 U89029 ( .A(n113895), .Z(n120622) );
  CLKBUF_X1 U89030 ( .A(n113892), .Z(n120628) );
  CLKBUF_X1 U89031 ( .A(n113767), .Z(n120826) );
endmodule

