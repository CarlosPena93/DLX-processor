
module registerfile_generic_n_bit32_data_bit64 ( CLK, RESET, ENABLE, RD1, RD2, 
        WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [5:0] ADD_WR;
  input [5:0] ADD_RD1;
  input [5:0] ADD_RD2;
  input [63:0] DATAIN;
  output [63:0] OUT1;
  output [63:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7489, n7505, n7521, n7537,
         n7553, n7569, n7585, n7601, n7617, n7633, n7649, n7665, n7681, n7697,
         n7713, n7729, n7745, n7761, n7777, n7793, n7809, n7825, n7841, n7857,
         n7873, n7889, n7905, n7921, n7937, n7953, n7969, n7985, n8001, n8017,
         n8033, n8049, n8065, n8081, n8097, n8113, n8129, n8145, n8161, n8177,
         n8193, n8209, n8225, n8241, n8257, n8273, n8289, n8305, n8321, n8337,
         n8353, n8369, n8385, n8401, n8417, n8433, n8449, n8461, n8465, n8477,
         n8481, n8493, n8497, n8509, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8961,
         n8963, n8965, n8967, n8969, n8971, n8973, n8975, n8977, n8979, n8981,
         n8983, n8985, n8987, n8989, n8991, n8993, n8995, n8997, n8999, n9001,
         n9003, n9005, n9007, n9009, n9011, n9013, n9015, n9017, n9019, n9021,
         n9023, n9025, n9027, n9029, n9031, n9033, n9035, n9037, n9039, n9041,
         n9043, n9045, n9047, n9049, n9051, n9053, n9055, n9057, n9059, n9061,
         n9063, n9065, n9067, n9069, n9071, n9073, n9075, n9077, n9079, n9081,
         n9083, n9085, n49228, n49229, n49230, n49231, n49232, n49233, n49234,
         n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
         n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250,
         n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
         n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266,
         n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
         n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282,
         n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290,
         n49291, n49420, n49421, n49422, n49423, n49424, n49425, n49426,
         n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434,
         n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
         n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450,
         n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458,
         n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466,
         n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
         n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482,
         n49483, n50517, n50518, n50519, n50520, n50521, n50522, n50523,
         n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531,
         n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539,
         n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547,
         n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555,
         n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563,
         n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571,
         n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579,
         n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651,
         n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659,
         n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667,
         n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675,
         n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683,
         n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691,
         n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699,
         n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707,
         n54184, n54185, n54186, n54187, n54188, n54189, n54190, n54191,
         n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199,
         n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207,
         n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215,
         n54216, n54217, n54218, n54219, n54220, n54221, n54222, n54223,
         n54224, n54225, n54226, n54227, n54228, n54229, n54230, n54231,
         n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239,
         n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54606,
         n54608, n54609, n54610, n54611, n54612, n54613, n54614, n54615,
         n54616, n54617, n54618, n54619, n54620, n54621, n54622, n54623,
         n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631,
         n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639,
         n54640, n54641, n54642, n54643, n54644, n54645, n54646, n54647,
         n54648, n54649, n54650, n54651, n54652, n54653, n54654, n54655,
         n54656, n54657, n54658, n54659, n54660, n54661, n54662, n54663,
         n54664, n54665, n54666, n54667, n54668, n54669, n54670, n56020,
         n56047, n56074, n56101, n56490, n56531, n56555, n56579, n56597,
         n56603, n56609, n56611, n56621, n56627, n56633, n56635, n56645,
         n56651, n56657, n56659, n56669, n56675, n56681, n56683, n56693,
         n56699, n56705, n56707, n56717, n56723, n56729, n56731, n56741,
         n56747, n56753, n56755, n56765, n56771, n56777, n56779, n56789,
         n56791, n56795, n56801, n56803, n56813, n56815, n56819, n56825,
         n56827, n56837, n56839, n56843, n56849, n56851, n56861, n56863,
         n56867, n56873, n56875, n56885, n56887, n56891, n56897, n56899,
         n56909, n56911, n56915, n56921, n56923, n56933, n56935, n56939,
         n56945, n56947, n56957, n56959, n56963, n56969, n56971, n56981,
         n56983, n56987, n56993, n56995, n57005, n57007, n57011, n57017,
         n57019, n57029, n57031, n57035, n57041, n57043, n57053, n57055,
         n57059, n57065, n57067, n57077, n57079, n57083, n57089, n57091,
         n57101, n57103, n57107, n57113, n57115, n57125, n57127, n57131,
         n57137, n57139, n57149, n57151, n57155, n57161, n57163, n57173,
         n57175, n57179, n57185, n57187, n57197, n57199, n57203, n57209,
         n57211, n57221, n57223, n57227, n57233, n57235, n57245, n57247,
         n57251, n57257, n57259, n57269, n57271, n57275, n57281, n57283,
         n57293, n57295, n57299, n57305, n57307, n57317, n57319, n57323,
         n57329, n57331, n57341, n57343, n57347, n57353, n57355, n57365,
         n57367, n57371, n57377, n57379, n57389, n57391, n57395, n57401,
         n57403, n57413, n57415, n57419, n57425, n57427, n57437, n57439,
         n57443, n57449, n57451, n57461, n57463, n57467, n57473, n57475,
         n57485, n57487, n57491, n57497, n57499, n57509, n57511, n57515,
         n57521, n57523, n57533, n57535, n57539, n57545, n57547, n57557,
         n57559, n57563, n57569, n57571, n57581, n57583, n57587, n57593,
         n57595, n57605, n57607, n57611, n57617, n57619, n57629, n57631,
         n57635, n57641, n57643, n57653, n57659, n57665, n57667, n57677,
         n57683, n57689, n57691, n57701, n57707, n57713, n57715, n57725,
         n57731, n57737, n57739, n57749, n57755, n57761, n57763, n57773,
         n57779, n57785, n57787, n57797, n57803, n57809, n57811, n57821,
         n57827, n57833, n57835, n57845, n57851, n57857, n57859, n57869,
         n57875, n57881, n57883, n57893, n57899, n57905, n57907, n57917,
         n57923, n57929, n57931, n57941, n57947, n57953, n57955, n57965,
         n57971, n57977, n57979, n57989, n57995, n58001, n58003, n58013,
         n58028, n58036, n58041, n58047, n58048, n58049, n58050, n58051,
         n58052, n58053, n58054, n58055, n58056, n58057, n58058, n58059,
         n58060, n58061, n58062, n58063, n58064, n58065, n58066, n58067,
         n58068, n58069, n58070, n58071, n58072, n58073, n58074, n58075,
         n58076, n58077, n58078, n58079, n58080, n58081, n58082, n58083,
         n58084, n58085, n58086, n58087, n58088, n58089, n58090, n58091,
         n58092, n58093, n58094, n58095, n58096, n58097, n58098, n58099,
         n58100, n58101, n58102, n58103, n58104, n58105, n58106, n58107,
         n58108, n58109, n58110, n58112, n58114, n58116, n58118, n58120,
         n58122, n58124, n58126, n58128, n58130, n58132, n58134, n58135,
         n58137, n58139, n58141, n58143, n58145, n58147, n58149, n58151,
         n58153, n58155, n58157, n58159, n58161, n58163, n58165, n58167,
         n58169, n58171, n58173, n58175, n58177, n58179, n58181, n58183,
         n58185, n58187, n58189, n58191, n58193, n58195, n58197, n58199,
         n58201, n58203, n58205, n58207, n58209, n58211, n58213, n58215,
         n58217, n58219, n58221, n58223, n58225, n58227, n58229, n58231,
         n58232, n58233, n58234, n58235, n58236, n58237, n58238, n58239,
         n58240, n58241, n58242, n58243, n58244, n58245, n58246, n58247,
         n58248, n58249, n58250, n58251, n58252, n58253, n58254, n58255,
         n58256, n58257, n58258, n58259, n58260, n58261, n58262, n58263,
         n58264, n58265, n58266, n58267, n58268, n58269, n58270, n58271,
         n58272, n58273, n58274, n58275, n58276, n58277, n58278, n58279,
         n58280, n58281, n58282, n58283, n58284, n58285, n58286, n58287,
         n58288, n58289, n58290, n58291, n58292, n58293, n58294, n58295,
         n58297, n58299, n58301, n58303, n58304, n58305, n58306, n58307,
         n58308, n58309, n58310, n58311, n58312, n58313, n58314, n58315,
         n58316, n58317, n58318, n58319, n58320, n58321, n58322, n58323,
         n58324, n58325, n58326, n58327, n58328, n58329, n58330, n58331,
         n58332, n58333, n58334, n58335, n58336, n58337, n58338, n58339,
         n58340, n58341, n58342, n58343, n58344, n58345, n58346, n58347,
         n58348, n58349, n58350, n58351, n58352, n58353, n58354, n58355,
         n58356, n58357, n58358, n58359, n58360, n58361, n58362, n58363,
         n58364, n58365, n58366, n58367, n58368, n58369, n58370, n58375,
         n58376, n58377, n58378, n58379, n58380, n58381, n58382, n58383,
         n58384, n58385, n58386, n58387, n58388, n58389, n58390, n58391,
         n58392, n58393, n58394, n58395, n58396, n58397, n58398, n58399,
         n58400, n58401, n58402, n58403, n58404, n58405, n58406, n58407,
         n58408, n58409, n58410, n58411, n58412, n58413, n58414, n58415,
         n58416, n58417, n58418, n58419, n58420, n58421, n58422, n58423,
         n58424, n58425, n58426, n58427, n58428, n58429, n58430, n58431,
         n58432, n58433, n58434, n58435, n58436, n58437, n58438, n58439,
         n58440, n58441, n58442, n58443, n58444, n58445, n58446, n58447,
         n58448, n58449, n58450, n58451, n58452, n58453, n58454, n58455,
         n58456, n58457, n58458, n58459, n58460, n58461, n58462, n58463,
         n58464, n58465, n58466, n58467, n58468, n58469, n58470, n58471,
         n58472, n58473, n58474, n58475, n58476, n58477, n58478, n58479,
         n58480, n58481, n58482, n58483, n58484, n58485, n58486, n58487,
         n58488, n58489, n58490, n58491, n58492, n58493, n58494, n58495,
         n58496, n58497, n58498, n58627, n58628, n58629, n58630, n58631,
         n58632, n58633, n58634, n58635, n58636, n58637, n58638, n58639,
         n58640, n58641, n58642, n58643, n58644, n58645, n58646, n58647,
         n58648, n58649, n58650, n58651, n58652, n58653, n58654, n58667,
         n58668, n58669, n58670, n58671, n58672, n58673, n58674, n58675,
         n58676, n58677, n58678, n58679, n58680, n58681, n58682, n58683,
         n58684, n58685, n58686, n58687, n58688, n58689, n58690, n58691,
         n58692, n58693, n58694, n58695, n58696, n58697, n58698, n58699,
         n58700, n58701, n58702, n58703, n58704, n58705, n58706, n58707,
         n58708, n58709, n58710, n58711, n58712, n58713, n58714, n58715,
         n58716, n58717, n58718, n58731, n58732, n58733, n58734, n58735,
         n58736, n58737, n58738, n58739, n58740, n58741, n58742, n58779,
         n58780, n58781, n58782, n58783, n58784, n58785, n58786, n58787,
         n58788, n58789, n58790, n58791, n58792, n58793, n58794, n58795,
         n58796, n58797, n58798, n58799, n58800, n58801, n58802, n58803,
         n58804, n58805, n58806, n58807, n58808, n58809, n58810, n58811,
         n58812, n58813, n58814, n58815, n58816, n58817, n58818, n58819,
         n58820, n58821, n58822, n58823, n58824, n58825, n58826, n58827,
         n58828, n58829, n58830, n58831, n58832, n58833, n58834, n58835,
         n58836, n58837, n58838, n58839, n58840, n58841, n58842, n58960,
         n59022, n59024, n59026, n59029, n59030, n59031, n59032, n59033,
         n59034, n59035, n59036, n59037, n59038, n59039, n59040, n59041,
         n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049,
         n59050, n59051, n59052, n59053, n59054, n59055, n59056, n59057,
         n59058, n59059, n59060, n59061, n59062, n59063, n59064, n59065,
         n59066, n59067, n59068, n59069, n59070, n59071, n59072, n59073,
         n59074, n59075, n59076, n59077, n59078, n59079, n59080, n59081,
         n59082, n59083, n59084, n59085, n59086, n59087, n59088, n59089,
         n59090, n59091, n59092, n61957, n61958, n61959, n61960, n61961,
         n61962, n61963, n61964, n61965, n61966, n61967, n61968, n61969,
         n61970, n61971, n61972, n61973, n61974, n61975, n61976, n61977,
         n61978, n61979, n61980, n61981, n61982, n61983, n61984, n61985,
         n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993,
         n61994, n61995, n61996, n61997, n61998, n61999, n62000, n62001,
         n62002, n62003, n62004, n62005, n62006, n62007, n62008, n62009,
         n62010, n62011, n62012, n62013, n62014, n62015, n62016, n62017,
         n62018, n62019, n62020, n62021, n62022, n62023, n62024, n62025,
         n62026, n62027, n62028, n62029, n62030, n62031, n62032, n62033,
         n62034, n62035, n62036, n62037, n62038, n62039, n62040, n62041,
         n62042, n62043, n62044, n62045, n62046, n62047, n62048, n62049,
         n62050, n62051, n62052, n62053, n62054, n62055, n62056, n62057,
         n62058, n62059, n62060, n62061, n62062, n62063, n62064, n62065,
         n62066, n62067, n62068, n62069, n62070, n62071, n62072, n62073,
         n62074, n62075, n62076, n62077, n62078, n62079, n62080, n62081,
         n62082, n62083, n62084, n62085, n62086, n62087, n62088, n62089,
         n62090, n62091, n62092, n62093, n62094, n62095, n62096, n62097,
         n62098, n62099, n62100, n62101, n62102, n62103, n62104, n62105,
         n62106, n62107, n62108, n62109, n62110, n62111, n62112, n62113,
         n62114, n62115, n62116, n62117, n62118, n62119, n62120, n62121,
         n62122, n62123, n62124, n62125, n62126, n62127, n62128, n62129,
         n62130, n62131, n62132, n62133, n62134, n62135, n62136, n62137,
         n62138, n62139, n62140, n62141, n62142, n62143, n62144, n62145,
         n62146, n62147, n62148, n62149, n62150, n62151, n62152, n62153,
         n62154, n62155, n62156, n62157, n62158, n62159, n62160, n62161,
         n62162, n62163, n62164, n62165, n62166, n62167, n62168, n62169,
         n62170, n62171, n62172, n62173, n62174, n62175, n62176, n62177,
         n62178, n62179, n62180, n62181, n62182, n62183, n62184, n62185,
         n62186, n62187, n62188, n62189, n62190, n62191, n62192, n62193,
         n62194, n62195, n62196, n62197, n62198, n62199, n62200, n62201,
         n62202, n62203, n62204, n62205, n62206, n62207, n62208, n62209,
         n62210, n62211, n62212, n62213, n62214, n62215, n62216, n62217,
         n62218, n62219, n62220, n62221, n62222, n62223, n62224, n62225,
         n62226, n62227, n62228, n62229, n62230, n62231, n62232, n62233,
         n62234, n62235, n62236, n62237, n62238, n62239, n62240, n62241,
         n62242, n62243, n62244, n62245, n62246, n62247, n62248, n62249,
         n62250, n62251, n62252, n62253, n62254, n62255, n62256, n62257,
         n62258, n62259, n62260, n62261, n62262, n62263, n62264, n62265,
         n62266, n62267, n62268, n62269, n62270, n62271, n62272, n62273,
         n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281,
         n62282, n62283, n62284, n62285, n62286, n62287, n62288, n62289,
         n62290, n62291, n62292, n62293, n62294, n62295, n62296, n62297,
         n62298, n62299, n62300, n62301, n62302, n62303, n62304, n62305,
         n62306, n62307, n62308, n62309, n62310, n62311, n62312, n62313,
         n62314, n62315, n62316, n62317, n62318, n62319, n62320, n62321,
         n62322, n62323, n62324, n62325, n62326, n62327, n62328, n62329,
         n62330, n62331, n62332, n62333, n62334, n62335, n62336, n62337,
         n62338, n62339, n62340, n62341, n62342, n62343, n62344, n62345,
         n62346, n62347, n62348, n62349, n62350, n62351, n62352, n62353,
         n62354, n62355, n62356, n62357, n62358, n62359, n62360, n62361,
         n62362, n62363, n62364, n62365, n62366, n62367, n62368, n62369,
         n62370, n62371, n62372, n62373, n62374, n62375, n62376, n62377,
         n62378, n62379, n62380, n62381, n62382, n62383, n62384, n62385,
         n62386, n62387, n62388, n62389, n62390, n62391, n62392, n62393,
         n62394, n62395, n62396, n62397, n62398, n62399, n62400, n62401,
         n62402, n62403, n62404, n62405, n62406, n62407, n62408, n62409,
         n62410, n62411, n62412, n62413, n62414, n62415, n62416, n62417,
         n62418, n62419, n62420, n62421, n62422, n62423, n62424, n62425,
         n62426, n62427, n62428, n62429, n62430, n62431, n62432, n62433,
         n62434, n62435, n62436, n62437, n62438, n62439, n62440, n62441,
         n62442, n62443, n62444, n62445, n62446, n62447, n62448, n62449,
         n62450, n62451, n62452, n62453, n62454, n62455, n62456, n62457,
         n62458, n62459, n62460, n62461, n62462, n62463, n62464, n62465,
         n62466, n62467, n62468, n62469, n62470, n62471, n62472, n62473,
         n62474, n62475, n62476, n62477, n62478, n62479, n62480, n62481,
         n62482, n62483, n62484, n62485, n62486, n62487, n62488, n62489,
         n62490, n62491, n62492, n62493, n62494, n62495, n62496, n62497,
         n62498, n62499, n62500, n62501, n62502, n62503, n62504, n62505,
         n62506, n62507, n62508, n62509, n62510, n62511, n62512, n62513,
         n62514, n62515, n62516, n62517, n62518, n62519, n62520, n62521,
         n62522, n62523, n62524, n62525, n62526, n62527, n62528, n62529,
         n62530, n62531, n62532, n62533, n62534, n62535, n62536, n62537,
         n62538, n62539, n62540, n62541, n62542, n62543, n62544, n62545,
         n62546, n62547, n62548, n62549, n62550, n62551, n62552, n62553,
         n62554, n62555, n62556, n62557, n62558, n62559, n62560, n62561,
         n62562, n62563, n62564, n62565, n62566, n62567, n62568, n62569,
         n62570, n62571, n62572, n62573, n62574, n62575, n62576, n62577,
         n62578, n62579, n62580, n62581, n62582, n62583, n62584, n62585,
         n62586, n62587, n62588, n62589, n62590, n62591, n62592, n62593,
         n62594, n62595, n62596, n62597, n62598, n62599, n62600, n62601,
         n62602, n62603, n62604, n62605, n62606, n62607, n62608, n62609,
         n62610, n62611, n62612, n62613, n62614, n62615, n62616, n62617,
         n62618, n62619, n62620, n62621, n62622, n62623, n62624, n62625,
         n62626, n62627, n62628, n62629, n62630, n62631, n62632, n62633,
         n62634, n62635, n62636, n62637, n62638, n62639, n62640, n62641,
         n62642, n62643, n62644, n62645, n62646, n62647, n62648, n62649,
         n62650, n62651, n62652, n62653, n62654, n62655, n62656, n62657,
         n62658, n62659, n62660, n62661, n62662, n62663, n62664, n62665,
         n62666, n62667, n62668, n62669, n62670, n62671, n62672, n62673,
         n62674, n62675, n62676, n62677, n62678, n62679, n62680, n62681,
         n62682, n62683, n62684, n62685, n62686, n62687, n62688, n62689,
         n62690, n62691, n62692, n62693, n62694, n62695, n62696, n62697,
         n62698, n62699, n62700, n62701, n62702, n62703, n62704, n62705,
         n62706, n62707, n62708, n62709, n62710, n62711, n62712, n62713,
         n62714, n62715, n62716, n62717, n62718, n62719, n62720, n62721,
         n62722, n62723, n62724, n62725, n62726, n62727, n62728, n62729,
         n62730, n62731, n62732, n62733, n62734, n62735, n62736, n62737,
         n62738, n62739, n62740, n62741, n62742, n62743, n62744, n62745,
         n62746, n62747, n62748, n62749, n62750, n62751, n62752, n62753,
         n62754, n62755, n62756, n62757, n62758, n62759, n62760, n62761,
         n62762, n62763, n62764, n62765, n62766, n62767, n62768, n62769,
         n62770, n62771, n62772, n62773, n62774, n62775, n62776, n62777,
         n62778, n62779, n62780, n62781, n62782, n62783, n62784, n62785,
         n62786, n62787, n62788, n62789, n62790, n62791, n62792, n62793,
         n62794, n62795, n62796, n62797, n62798, n62799, n62800, n62801,
         n62802, n62803, n62804, n62805, n62806, n62807, n62808, n62809,
         n62810, n62811, n62812, n62813, n62814, n62815, n62816, n62817,
         n62818, n62819, n62820, n62821, n62822, n62823, n62824, n62825,
         n62826, n62827, n62828, n62829, n62830, n62831, n62832, n62833,
         n62834, n62835, n62836, n62837, n62838, n62839, n62840, n62841,
         n62842, n62843, n62844, n62845, n62846, n62847, n62848, n62849,
         n62850, n62851, n62852, n62853, n62854, n62855, n62856, n62857,
         n62858, n62859, n62860, n62861, n62862, n62863, n62864, n62865,
         n62866, n62867, n62868, n62869, n62870, n62871, n62872, n62873,
         n62874, n62875, n62876, n62877, n62878, n62879, n62880, n62881,
         n62882, n62883, n62884, n62885, n62886, n62887, n62888, n62889,
         n62890, n62891, n62892, n62893, n62894, n62895, n62896, n62897,
         n62898, n62899, n62900, n62901, n62902, n62903, n62904, n62905,
         n62906, n62907, n62908, n62909, n62910, n62911, n62912, n62913,
         n62914, n62915, n62916, n62917, n62918, n62919, n62920, n62921,
         n62922, n62923, n62924, n62925, n62926, n62927, n62928, n62929,
         n62930, n62931, n62932, n62933, n62934, n62935, n62936, n62937,
         n62938, n62939, n62940, n62941, n62942, n62943, n62944, n62945,
         n62946, n62947, n62948, n62949, n62950, n62951, n62952, n62953,
         n62954, n62955, n62956, n62957, n62958, n62959, n62960, n62961,
         n62962, n62963, n62964, n62965, n62966, n62967, n62968, n62969,
         n62970, n62971, n62972, n62973, n62974, n62975, n62976, n62977,
         n62978, n62979, n62980, n62981, n62982, n62983, n62984, n62985,
         n62986, n62987, n62988, n62989, n62990, n62991, n62992, n62993,
         n62994, n62995, n62996, n62997, n62998, n62999, n63000, n63001,
         n63002, n63003, n63004, n63005, n63006, n63007, n63008, n63009,
         n63010, n63011, n63012, n63013, n63014, n63015, n63016, n63017,
         n63018, n63019, n63020, n63021, n63022, n63023, n63024, n63025,
         n63026, n63027, n63028, n63029, n63030, n63031, n63032, n63033,
         n63034, n63035, n63036, n63037, n63038, n63039, n63040, n63041,
         n63042, n63043, n63044, n63045, n63046, n63047, n63048, n63049,
         n63050, n63051, n63052, n63053, n63054, n63055, n63056, n63057,
         n63058, n63059, n63060, n63061, n63062, n63063, n63064, n63065,
         n63066, n63067, n63068, n63069, n63070, n63071, n63072, n63073,
         n63074, n63075, n63076, n63077, n63078, n63079, n63080, n63081,
         n63082, n63083, n63084, n63085, n63086, n63087, n63088, n63089,
         n63090, n63091, n63092, n63093, n63094, n63095, n63096, n63097,
         n63098, n63099, n63100, n63101, n63102, n63103, n63104, n63105,
         n63106, n63107, n63108, n63109, n63110, n63111, n63112, n63113,
         n63114, n63115, n63116, n63117, n63118, n63119, n63120, n63121,
         n63122, n63123, n63124, n63125, n63126, n63127, n63128, n63129,
         n63130, n63131, n63132, n63133, n63134, n63135, n63136, n63137,
         n63138, n63139, n63140, n63141, n63142, n63143, n63144, n63145,
         n63146, n63147, n63148, n63149, n63150, n63151, n63152, n63153,
         n63154, n63155, n63156, n63157, n63158, n63159, n63160, n63161,
         n63162, n63163, n63164, n63165, n63166, n63167, n63168, n63169,
         n63170, n63171, n63172, n63173, n63174, n63175, n63176, n63177,
         n63178, n63179, n63180, n63181, n63182, n63183, n63184, n63185,
         n63186, n63187, n63188, n63189, n63190, n63191, n63192, n63193,
         n63194, n63195, n63196, n63197, n63198, n63199, n63200, n63201,
         n63202, n63203, n63204, n63205, n63206, n63207, n63208, n63209,
         n63210, n63211, n63212, n63213, n63214, n63215, n63216, n63217,
         n63218, n63219, n63220, n63221, n63222, n63223, n63224, n63225,
         n63226, n63227, n63228, n63229, n63230, n63231, n63232, n63233,
         n63234, n63235, n63236, n63237, n63238, n63239, n63240, n63241,
         n63242, n63243, n63244, n63245, n63246, n63247, n63248, n63249,
         n63250, n63251, n63252, n63253, n63254, n63255, n63256, n63257,
         n63258, n63259, n63260, n63261, n63262, n63263, n63264, n63265,
         n63266, n63267, n63268, n63269, n63270, n63271, n63272, n63273,
         n63274, n63275, n63276, n63277, n63278, n63279, n63280, n63281,
         n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289,
         n63290, n63291, n63292, n63293, n63294, n63295, n63296, n63297,
         n63298, n63299, n63300, n63301, n63302, n63303, n63304, n63305,
         n63306, n63307, n63308, n63309, n63310, n63311, n63312, n63313,
         n63314, n63315, n63316, n63317, n63318, n63319, n63320, n63321,
         n63322, n63323, n63324, n63325, n63326, n63327, n63328, n63329,
         n63330, n63331, n63332, n63333, n63334, n63335, n63336, n63337,
         n63338, n63339, n63340, n63341, n63342, n63343, n63344, n63345,
         n63346, n63347, n63348, n63349, n63350, n63351, n63352, n63353,
         n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361,
         n63362, n63363, n63364, n63365, n63366, n63367, n63368, n63369,
         n63370, n63371, n63372, n63373, n63374, n63375, n63376, n63377,
         n63378, n63379, n63380, n63381, n63382, n63383, n63384, n63385,
         n63386, n63387, n63388, n63389, n63390, n63391, n63392, n63393,
         n63394, n63395, n63396, n63397, n63398, n63399, n63400, n63401,
         n63402, n63403, n63404, n63405, n63406, n63407, n63408, n63409,
         n63410, n63411, n63412, n63413, n63414, n63415, n63416, n63417,
         n63418, n63419, n63420, n63421, n63422, n63423, n63424, n63425,
         n63426, n63427, n63428, n63429, n63430, n63431, n63432, n63433,
         n63434, n63435, n63436, n63437, n63438, n63439, n63440, n63441,
         n63442, n63443, n63444, n63445, n63446, n63447, n63448, n63449,
         n63450, n63451, n63452, n63453, n63454, n63455, n63456, n63457,
         n63458, n63459, n63460, n63461, n63462, n63463, n63464, n63465,
         n63466, n63467, n63468, n63469, n63470, n63471, n63472, n63473,
         n63474, n63475, n63476, n63477, n63478, n63479, n63480, n63481,
         n63482, n63483, n63484, n63485, n63486, n63487, n63488, n63489,
         n63490, n63491, n63492, n63493, n63494, n63495, n63496, n63497,
         n63498, n63499, n63500, n63501, n63502, n63503, n63504, n63505,
         n63506, n63507, n63508, n63509, n63510, n63511, n63512, n63513,
         n63514, n63515, n63516, n63517, n63518, n63519, n63520, n63521,
         n63522, n63523, n63524, n63525, n63526, n63527, n63528, n63529,
         n63530, n63531, n63532, n63533, n63534, n63535, n63536, n63537,
         n63538, n63539, n63540, n63541, n63542, n63543, n63544, n63545,
         n63546, n63547, n63548, n63549, n63550, n63551, n63552, n63553,
         n63554, n63555, n63556, n63557, n63558, n63559, n63560, n63561,
         n63562, n63563, n63564, n63565, n63566, n63567, n63568, n63569,
         n63570, n63571, n63572, n63573, n63574, n63575, n63576, n63577,
         n63578, n63579, n63580, n63581, n63582, n63583, n63584, n63585,
         n63586, n63587, n63588, n63589, n63590, n63591, n63592, n63593,
         n63594, n63595, n63596, n63597, n63598, n63599, n63600, n63601,
         n63602, n63603, n63604, n63605, n63606, n63607, n63608, n63609,
         n63610, n63611, n63612, n63613, n63614, n63615, n63616, n63617,
         n63618, n63619, n63620, n63621, n63622, n63623, n63624, n63625,
         n63626, n63627, n63628, n63629, n63630, n63631, n63632, n63633,
         n63634, n63635, n63636, n63637, n63638, n63639, n63640, n63641,
         n63642, n63643, n63644, n63645, n63646, n63647, n63648, n63649,
         n63650, n63651, n63652, n63653, n63654, n63655, n63656, n63657,
         n63658, n63659, n63660, n63661, n63662, n63663, n63664, n63665,
         n63666, n63667, n63668, n63669, n63670, n63671, n63672, n63673,
         n63674, n63675, n63676, n63677, n63678, n63679, n63680, n63681,
         n63682, n63683, n63684, n63685, n63686, n63687, n63688, n63689,
         n63690, n63691, n63692, n63693, n63694, n63695, n63696, n63697,
         n63698, n63699, n63700, n63701, n63702, n63703, n63704, n63705,
         n63706, n63707, n63708, n63709, n63710, n63711, n63712, n63713,
         n63714, n63715, n63716, n63717, n63718, n63719, n63720, n63721,
         n63722, n63723, n63724, n63725, n63726, n63727, n63728, n63729,
         n63730, n63731, n63732, n63733, n63734, n63735, n63736, n63737,
         n63738, n63739, n63740, n63741, n63742, n63743, n63744, n63745,
         n63746, n63747, n63748, n63749, n63750, n63751, n63752, n63753,
         n63754, n63755, n63756, n63757, n63758, n63759, n63760, n63761,
         n63762, n63763, n63764, n63765, n63766, n63767, n63768, n63769,
         n63770, n63771, n63772, n63773, n63774, n63775, n63776, n63777,
         n63778, n63780, n63781, n63782, n63783, n63784, n63785, n63786,
         n63787, n63788, n63790, n63791, n63792, n63793, n63794, n63795,
         n63797, n63798, n63799, n63800, n63801, n63802, n63803, n63804,
         n63805, n63806, n63807, n63808, n63809, n63810, n63811, n63812,
         n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820,
         n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828,
         n63829, n63830, n63831, n63833, n63835, n63836, n63837, n63838,
         n63839, n63840, n63841, n63842, n63843, n63844, n63845, n63846,
         n63847, n63848, n63849, n63850, n63851, n63852, n63854, n63856,
         n63857, n63858, n63859, n63860, n63861, n63862, n63863, n63864,
         n63865, n63866, n63867, n63868, n63869, n63870, n63871, n63872,
         n63873, n63875, n63877, n63878, n63879, n63880, n63881, n63882,
         n63883, n63884, n63885, n63886, n63887, n63888, n63889, n63890,
         n63891, n63892, n63893, n63894, n63896, n63897, n63898, n63899,
         n63900, n63901, n63902, n63903, n63904, n63905, n63906, n63907,
         n63908, n63909, n63910, n63911, n63912, n63913, n63914, n63916,
         n63917, n63918, n63919, n63920, n63921, n63922, n63923, n63924,
         n63925, n63926, n63927, n63928, n63929, n63930, n63931, n63932,
         n63933, n63934, n63936, n63937, n63938, n63939, n63940, n63941,
         n63942, n63943, n63944, n63945, n63946, n63947, n63948, n63949,
         n63950, n63951, n63952, n63953, n63954, n63956, n63957, n63958,
         n63959, n63960, n63961, n63962, n63963, n63964, n63965, n63966,
         n63967, n63968, n63969, n63970, n63971, n63972, n63973, n63974,
         n63976, n63977, n63978, n63979, n63980, n63981, n63982, n63983,
         n63984, n63985, n63986, n63987, n63988, n63989, n63990, n63991,
         n63992, n63993, n63994, n63996, n63997, n63998, n63999, n64000,
         n64001, n64002, n64003, n64004, n64005, n64006, n64007, n64008,
         n64009, n64010, n64011, n64012, n64013, n64014, n64016, n64017,
         n64018, n64019, n64020, n64021, n64022, n64023, n64024, n64025,
         n64026, n64027, n64028, n64029, n64030, n64031, n64032, n64033,
         n64034, n64036, n64037, n64038, n64039, n64040, n64041, n64042,
         n64043, n64044, n64045, n64046, n64047, n64048, n64049, n64050,
         n64051, n64052, n64053, n64054, n64056, n64057, n64058, n64059,
         n64060, n64061, n64062, n64063, n64064, n64065, n64066, n64067,
         n64068, n64069, n64070, n64071, n64072, n64073, n64074, n64076,
         n64077, n64078, n64079, n64080, n64081, n64082, n64083, n64084,
         n64085, n64086, n64087, n64088, n64089, n64090, n64091, n64092,
         n64093, n64094, n64096, n64097, n64098, n64099, n64100, n64101,
         n64102, n64103, n64104, n64105, n64106, n64107, n64108, n64109,
         n64110, n64111, n64112, n64113, n64114, n64116, n64117, n64118,
         n64119, n64120, n64121, n64122, n64123, n64124, n64125, n64126,
         n64127, n64128, n64129, n64130, n64131, n64132, n64133, n64134,
         n64136, n64137, n64138, n64139, n64140, n64141, n64142, n64143,
         n64144, n64145, n64146, n64147, n64148, n64149, n64150, n64151,
         n64152, n64153, n64154, n64156, n64157, n64158, n64159, n64160,
         n64161, n64162, n64163, n64164, n64165, n64166, n64167, n64168,
         n64169, n64170, n64171, n64172, n64173, n64174, n64176, n64177,
         n64178, n64179, n64180, n64181, n64182, n64183, n64184, n64185,
         n64186, n64187, n64188, n64189, n64190, n64191, n64192, n64193,
         n64194, n64196, n64197, n64198, n64199, n64200, n64201, n64202,
         n64203, n64204, n64205, n64206, n64207, n64208, n64209, n64210,
         n64211, n64212, n64213, n64214, n64216, n64217, n64218, n64219,
         n64220, n64221, n64222, n64223, n64224, n64225, n64226, n64227,
         n64228, n64229, n64230, n64231, n64232, n64233, n64234, n64236,
         n64237, n64238, n64239, n64240, n64241, n64242, n64243, n64244,
         n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64252,
         n64253, n64254, n64256, n64257, n64258, n64259, n64260, n64261,
         n64262, n64263, n64264, n64265, n64266, n64267, n64268, n64269,
         n64270, n64271, n64272, n64273, n64274, n64276, n64277, n64278,
         n64279, n64280, n64281, n64282, n64283, n64284, n64285, n64286,
         n64287, n64288, n64289, n64290, n64291, n64292, n64293, n64294,
         n64296, n64297, n64298, n64299, n64300, n64301, n64302, n64303,
         n64304, n64305, n64306, n64307, n64308, n64309, n64310, n64311,
         n64312, n64313, n64314, n64316, n64317, n64318, n64319, n64320,
         n64321, n64322, n64323, n64324, n64325, n64326, n64327, n64328,
         n64329, n64330, n64331, n64332, n64333, n64334, n64336, n64337,
         n64338, n64339, n64340, n64341, n64342, n64343, n64344, n64345,
         n64346, n64347, n64348, n64349, n64350, n64351, n64352, n64353,
         n64354, n64356, n64357, n64358, n64359, n64360, n64361, n64362,
         n64363, n64364, n64365, n64366, n64367, n64368, n64369, n64370,
         n64371, n64372, n64373, n64374, n64376, n64377, n64378, n64379,
         n64380, n64381, n64382, n64383, n64384, n64385, n64386, n64387,
         n64388, n64389, n64390, n64391, n64392, n64393, n64394, n64396,
         n64397, n64398, n64399, n64400, n64401, n64402, n64403, n64404,
         n64405, n64406, n64407, n64408, n64409, n64410, n64411, n64412,
         n64413, n64414, n64416, n64417, n64418, n64419, n64420, n64421,
         n64422, n64423, n64424, n64425, n64426, n64427, n64428, n64429,
         n64430, n64431, n64432, n64433, n64434, n64436, n64437, n64438,
         n64439, n64440, n64441, n64442, n64443, n64444, n64445, n64446,
         n64447, n64448, n64449, n64450, n64451, n64452, n64453, n64454,
         n64456, n64457, n64458, n64459, n64460, n64461, n64462, n64463,
         n64464, n64465, n64466, n64467, n64468, n64469, n64470, n64471,
         n64472, n64473, n64474, n64476, n64477, n64478, n64479, n64480,
         n64481, n64482, n64483, n64484, n64485, n64486, n64487, n64488,
         n64489, n64490, n64491, n64492, n64493, n64494, n64496, n64497,
         n64498, n64499, n64500, n64501, n64502, n64503, n64504, n64505,
         n64506, n64507, n64508, n64509, n64510, n64511, n64512, n64513,
         n64514, n64516, n64517, n64518, n64519, n64520, n64521, n64522,
         n64523, n64524, n64525, n64526, n64527, n64528, n64529, n64530,
         n64531, n64532, n64533, n64534, n64536, n64537, n64538, n64539,
         n64540, n64541, n64542, n64543, n64544, n64545, n64546, n64547,
         n64548, n64549, n64550, n64551, n64552, n64553, n64554, n64556,
         n64557, n64558, n64559, n64560, n64561, n64562, n64563, n64564,
         n64565, n64566, n64567, n64568, n64569, n64570, n64571, n64572,
         n64573, n64574, n64576, n64577, n64578, n64579, n64580, n64581,
         n64582, n64583, n64584, n64585, n64586, n64587, n64588, n64589,
         n64590, n64591, n64592, n64593, n64594, n64596, n64597, n64598,
         n64599, n64600, n64601, n64602, n64603, n64604, n64605, n64606,
         n64607, n64608, n64609, n64610, n64611, n64612, n64613, n64614,
         n64616, n64617, n64618, n64619, n64620, n64621, n64622, n64623,
         n64624, n64625, n64626, n64627, n64628, n64629, n64630, n64631,
         n64632, n64633, n64634, n64636, n64637, n64638, n64639, n64640,
         n64641, n64642, n64643, n64644, n64645, n64646, n64647, n64648,
         n64649, n64650, n64651, n64652, n64653, n64654, n64656, n64657,
         n64658, n64659, n64660, n64661, n64662, n64663, n64664, n64665,
         n64666, n64667, n64668, n64669, n64670, n64671, n64672, n64673,
         n64674, n64676, n64677, n64678, n64679, n64680, n64681, n64682,
         n64683, n64684, n64685, n64686, n64687, n64688, n64689, n64690,
         n64691, n64692, n64693, n64694, n64696, n64697, n64698, n64699,
         n64700, n64701, n64702, n64703, n64704, n64705, n64706, n64707,
         n64708, n64709, n64710, n64711, n64712, n64713, n64714, n64716,
         n64717, n64718, n64719, n64720, n64721, n64722, n64723, n64724,
         n64725, n64726, n64727, n64728, n64729, n64730, n64731, n64732,
         n64733, n64734, n64736, n64737, n64738, n64739, n64740, n64741,
         n64742, n64743, n64744, n64745, n64746, n64747, n64748, n64749,
         n64750, n64751, n64752, n64753, n64754, n64756, n64757, n64758,
         n64759, n64760, n64761, n64762, n64763, n64764, n64765, n64766,
         n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774,
         n64776, n64777, n64778, n64779, n64780, n64781, n64782, n64783,
         n64784, n64785, n64786, n64787, n64788, n64789, n64790, n64791,
         n64792, n64793, n64794, n64796, n64797, n64798, n64799, n64800,
         n64801, n64802, n64803, n64804, n64805, n64806, n64807, n64808,
         n64809, n64810, n64811, n64812, n64813, n64814, n64816, n64817,
         n64818, n64819, n64820, n64821, n64822, n64823, n64824, n64825,
         n64826, n64827, n64828, n64829, n64830, n64831, n64832, n64833,
         n64834, n64836, n64837, n64838, n64839, n64840, n64841, n64842,
         n64843, n64844, n64845, n64846, n64847, n64848, n64849, n64850,
         n64851, n64852, n64853, n64854, n64855, n64856, n64857, n64858,
         n64859, n64860, n64861, n64862, n64863, n64864, n64865, n64866,
         n64867, n64868, n64869, n64870, n64871, n64872, n64873, n64874,
         n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882,
         n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890,
         n64891, n64892, n64893, n64894, n64895, n64896, n64897, n64898,
         n64899, n64900, n64901, n64902, n64903, n64904, n64905, n64906,
         n64907, n64908, n64909, n64910, n64911, n64912, n64913, n64914,
         n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922,
         n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930,
         n64931, n64932, n64933, n64934, n64935, n64936, n64937, n64938,
         n64939, n64940, n64941, n64942, n64943, n64944, n64945, n64946,
         n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954,
         n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962,
         n64963, n64964, n64965, n64966, n64967, n64968, n64969, n64970,
         n64971, n64972, n64973, n64974, n64975, n64976, n64977, n64978,
         n64979, n64980, n64981, n64982, n64983, n64984, n64985, n64986,
         n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994,
         n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002,
         n65003, n65004, n65005, n65006, n65007, n65008, n65009, n65010,
         n65011, n65012, n65013, n65014, n65015, n65016, n65017, n65018,
         n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026,
         n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034,
         n65035, n65036, n65037, n65038, n65039, n65040, n65041, n65042,
         n65043, n65044, n65045, n65046, n65047, n65048, n65049, n65050,
         n65051, n65052, n65053, n65054, n65055, n65056, n65057, n65058,
         n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066,
         n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074,
         n65075, n65076, n65077, n65078, n65079, n65080, n65081, n65082,
         n65083, n65084, n65085, n65086, n65087, n65088, n65089, n65090,
         n65091, n65092, n65093, n65094, n65095, n65096, n65098, n65099,
         n65100, n65101, n65102, n65103, n65104, n65105, n65106, n65107,
         n65108, n65109, n65110, n65111, n65112, n65113, n65114, n65115,
         n65116, n65117, n65118, n65119, n65120, n65121, n65122, n65123,
         n65124, n65125, n65126, n65127, n65128, n65129, n65130, n65131,
         n65132, n65133, n65134, n65135, n65136, n65137, n65138, n65139,
         n65140, n65141, n65142, n65143, n65144, n65145, n65146, n65147,
         n65148, n65149, n65150, n65151, n65152, n65153, n65154, n65155,
         n65156, n65157, n65158, n65159, n65160, n65161, n65162, n65163,
         n65164, n65165, n65166, n65167, n65168, n65169, n65170, n65171,
         n65172, n65173, n65174, n65175, n65176, n65177, n65178, n65179,
         n65180, n65181, n65182, n65183, n65184, n65185, n65186, n65187,
         n65188, n65189, n65190, n65191, n65192, n65193, n65194, n65195,
         n65196, n65197, n65198, n65199, n65200, n65201, n65202, n65203,
         n65204, n65205, n65206, n65207, n65208, n65209, n65210, n65211,
         n65212, n65213, n65214, n65215, n65216, n65217, n65218, n65219,
         n65220, n65221, n65222, n65223, n65224, n65225, n65226, n65227,
         n65228, n65229, n65230, n65231, n65232, n65233, n65234, n65235,
         n65236, n65237, n65238, n65239, n65240, n65241, n65242, n65243,
         n65244, n65245, n65246, n65247, n65248, n65249, n65250, n65251,
         n65252, n65253, n65254, n65255, n65256, n65257, n65258, n65259,
         n65260, n65261, n65262, n65263, n65264, n65265, n65266, n65267,
         n65268, n65269, n65270, n65271, n65272, n65273, n65274, n65275,
         n65276, n65277, n65278, n65279, n65280, n65281, n65282, n65283,
         n65284, n65285, n65286, n65287, n65288, n65289, n65290, n65291,
         n65292, n65293, n65294, n65295, n65296, n65297, n65298, n65299,
         n65300, n65301, n65302, n65303, n65304, n65305, n65306, n65307,
         n65308, n65309, n65310, n65311, n65312, n65313, n65314, n65315,
         n65316, n65317, n65318, n65319, n65320, n65321, n65322, n65323,
         n65324, n65325, n65326, n65327, n65328, n65329, n65330, n65331,
         n65332, n65333, n65334, n65335, n65336, n65337, n65338, n65339,
         n65340, n65341, n65342, n65343, n65344, n65345, n65346, n65347,
         n65348, n65349, n65350, n65351, n65352, n65353, n65354, n65355,
         n65356, n65357, n65358, n65359, n65360, n65361, n65362, n65363,
         n65364, n65365, n65366, n65367, n65368, n65369, n65370, n65371,
         n65372, n65373, n65374, n65375, n65376, n65377, n65378, n65379,
         n65380, n65381, n65382, n65383, n65384, n65385, n65386, n65387,
         n65388, n65389, n65390, n65391, n65392, n65393, n65394, n65395,
         n65396, n65397, n65398, n65399, n65400, n65401, n65402, n65403,
         n65404, n65405, n65406, n65407, n65408, n65409, n65410, n65411,
         n65412, n65413, n65414, n65415, n65416, n65417, n65418, n65419,
         n65420, n65421, n65422, n65423, n65424, n65425, n65426, n65427,
         n65428, n65429, n65430, n65431, n65432, n65433, n65434, n65435,
         n65436, n65437, n65438, n65439, n65440, n65441, n65442, n65443,
         n65444, n65445, n65446, n65447, n65448, n65449, n65450, n65451,
         n65452, n65453, n65454, n65455, n65456, n65457, n65458, n65459,
         n65460, n65461, n65462, n65463, n65464, n65465, n65466, n65467,
         n65468, n65469, n65470, n65471, n65472, n65473, n65474, n65475,
         n65476, n65477, n65478, n65479, n65480, n65481, n65482, n65483,
         n65484, n65485, n65486, n65487, n65488, n65489, n65490, n65491,
         n65492, n65493, n65494, n65495, n65496, n65497, n65498, n65499,
         n65500, n65501, n65502, n65503, n65504, n65505, n65506, n65507,
         n65508, n65509, n65510, n65511, n65512, n65513, n65514, n65515,
         n65516, n65517, n65518, n65519, n65520, n65521, n65522, n65523,
         n65524, n65525, n65526, n65527, n65528, n65529, n65530, n65531,
         n65532, n65533, n65534, n65535, n65536, n65537, n65538, n65539,
         n65540, n65541, n65542, n65543, n65544, n65545, n65546, n65547,
         n65548, n65549, n65550, n65551, n65552, n65553, n65554, n65555,
         n65556, n65557, n65558, n65559, n65560, n65561, n65562, n65563,
         n65564, n65565, n65566, n65567, n65568, n65569, n65570, n65571,
         n65572, n65573, n65574, n65575, n65576, n65577, n65578, n65579,
         n65580, n65581, n65582, n65583, n65584, n65585, n65586, n65587,
         n65588, n65589, n65590, n65591, n65592, n65593, n65594, n65595,
         n65596, n65597, n65598, n65599, n65600, n65601, n65602, n65603,
         n65604, n65605, n65606, n65607, n65608, n65609, n65610, n65611,
         n65612, n65613, n65614, n65615, n65616, n65617, n65618, n65619,
         n65620, n65621, n65622, n65623, n65624, n65625, n65626, n65627,
         n65628, n65629, n65630, n65631, n65632, n65633, n65634, n65635,
         n65636, n65637, n65638, n65639, n65640, n65641, n65642, n65643,
         n65644, n65645, n65646, n65647, n65648, n65649, n65650, n65651,
         n65652, n65653, n65654, n65655, n65656, n65657, n65658, n65659,
         n65660, n65661, n65662, n65663, n65664, n65665, n65666, n65667,
         n65668, n65669, n65670, n65671, n65672, n65673, n65674, n65675,
         n65676, n65677, n65678, n65679, n65680, n65681, n65682, n65683,
         n65684, n65685, n65686, n65687, n65688, n65689, n65690, n65691,
         n65692, n65693, n65694, n65695, n65696, n65697, n65698, n65699,
         n65700, n65701, n65702, n65703, n65704, n65705, n65706, n65707,
         n65708, n65709, n65710, n65711, n65712, n65713, n65714, n65715,
         n65716, n65717, n65718, n65719, n65720, n65721, n65722, n65723,
         n65724, n65725, n65726, n65727, n65728, n65729, n65730, n65731,
         n65732, n65733, n65734, n65735, n65736, n65737, n65738, n65739,
         n65740, n65741, n65742, n65743, n65744, n65745, n65746, n65747,
         n65748, n65749, n65750, n65751, n65752, n65753, n65754, n65755,
         n65756, n65757, n65758, n65759, n65760, n65761, n65762, n65763,
         n65764, n65765, n65766, n65767, n65768, n65769, n65770, n65771,
         n65772, n65773, n65774, n65775, n65776, n65777, n65778, n65779,
         n65780, n65781, n65782, n65783, n65784, n65785, n65786, n65787,
         n65788, n65789, n65790, n65791, n65792, n65793, n65794, n65795,
         n65796, n65797, n65798, n65799, n65800, n65801, n65802, n65803,
         n65804, n65805, n65806, n65807, n65808, n65809, n65810, n65811,
         n65812, n65813, n65814, n65815, n65816, n65817, n65818, n65819,
         n65820, n65821, n65822, n65823, n65824, n65825, n65826, n65827,
         n65828, n65829, n65830, n65831, n65832, n65833, n65834, n65835,
         n65836, n65837, n65838, n65839, n65840, n65841, n65842, n65843,
         n65844, n65845, n65846, n65847, n65848, n65849, n65850, n65851,
         n65852, n65853, n65854, n65855, n65856, n65857, n65858, n65859,
         n65860, n65861, n65862, n65863, n65864, n65865, n65866, n65867,
         n65868, n65869, n65870, n65871, n65872, n65873, n65874, n65875,
         n65876, n65877, n65878, n65879, n65880, n65881, n65882, n65883,
         n65884, n65885, n65886, n65887, n65888, n65889, n65890, n65891,
         n65892, n65893, n65894, n65895, n65896, n65897, n65898, n65899,
         n65900, n65901, n65902, n65903, n65904, n65905, n65906, n65907,
         n65908, n65909, n65910, n65911, n65912, n65913, n65914, n65915,
         n65916, n65917, n65918, n65919, n65920, n65921, n65922, n65923,
         n65924, n65925, n65926, n65927, n65928, n65929, n65930, n65931,
         n65932, n65933, n65934, n65935, n65936, n65937, n65938, n65939,
         n65940, n65941, n65942, n65943, n65944, n65945, n65946, n65947,
         n65948, n65949, n65950, n65951, n65952, n65953, n65954, n65955,
         n65956, n65957, n65958, n65959, n65960, n65961, n65962, n65963,
         n65964, n65965, n65966, n65967, n65968, n65969, n65970, n65971,
         n65972, n65973, n65974, n65975, n65976, n65977, n65978, n65979,
         n65980, n65981, n65982, n65983, n65984, n65985, n65986, n65987,
         n65988, n65989, n65990, n65991, n65992, n65993, n65994, n65995,
         n65996, n65997, n65998, n65999, n66000, n66001, n66002, n66003,
         n66004, n66005, n66006, n66007, n66008, n66009, n66010, n66011,
         n66012, n66013, n66014, n66015, n66016, n66017, n66018, n66019,
         n66020, n66021, n66022, n66023, n66024, n66025, n66026, n66027,
         n66028, n66029, n66030, n66031, n66032, n66033, n66034, n66035,
         n66036, n66037, n66038, n66039, n66040, n66041, n66042, n66043,
         n66044, n66045, n66046, n66047, n66048, n66049, n66050, n66051,
         n66052, n66053, n66054, n66055, n66056, n66057, n66058, n66059,
         n66060, n66061, n66062, n66063, n66064, n66065, n66066, n66067,
         n66068, n66069, n66070, n66071, n66072, n66073, n66074, n66075,
         n66076, n66077, n66078, n66079, n66080, n66081, n66082, n66083,
         n66084, n66085, n66086, n66087, n66088, n66089, n66090, n66091,
         n66092, n66093, n66094, n66095, n66096, n66097, n66098, n66099,
         n66100, n66101, n66102, n66103, n66104, n66105, n66106, n66107,
         n66108, n66109, n66110, n66111, n66112, n66113, n66114, n66115,
         n66116, n66117, n66118, n66119, n66120, n66121, n66122, n66123,
         n66124, n66125, n66126, n66127, n66128, n66129, n66130, n66131,
         n66132, n66133, n66134, n66135, n66136, n66137, n66138, n66139,
         n66140, n66141, n66142, n66143, n66144, n66145, n66146, n66147,
         n66148, n66149, n66150, n66151, n66152, n66153, n66154, n66155,
         n66156, n66157, n66158, n66159, n66160, n66161, n66162, n66163,
         n66164, n66165, n66166, n66167, n66168, n66169, n66170, n66171,
         n66172, n66173, n66174, n66175, n66176, n66177, n66178, n66179,
         n66180, n66181, n66182, n66183, n66184, n66185, n66186, n66187,
         n66188, n66189, n66190, n66191, n66192, n66193, n66194, n66195,
         n66196, n66197, n66198, n66199, n66200, n66201, n66202, n66203,
         n66204, n66205, n66206, n66207, n66208, n66209, n66210, n66211,
         n66212, n66213, n66214, n66215, n66216, n66217, n66218, n66219,
         n66220, n66221, n66222, n66223, n66224, n66225, n66226, n66227,
         n66228, n66229, n66230, n66231, n66232, n66233, n66234, n66235,
         n66236, n66237, n66238, n66239, n66240, n66241, n66242, n66243,
         n66244, n66245, n66246, n66247, n66248, n66249, n66250, n66251,
         n66252, n66253, n66254, n66255, n66256, n66257, n66258, n66259,
         n66260, n66261, n66262, n66263, n66264, n66265, n66266, n66267,
         n66268, n66269, n66270, n66271, n66272, n66273, n66274, n66275,
         n66276, n66277, n66278, n66279, n66280, n66281, n66282, n66283,
         n66284, n66285, n66286, n66287, n66288, n66289, n66290, n66291,
         n66292, n66293, n66294, n66295, n66296, n66297, n66298, n66299,
         n66300, n66301, n66305, n66306, n66307, n66308, n66313, n66314,
         n66315, n66316, n66317, n66318, n66319, n66320, n66321, n66322,
         n66323, n66324, n66325, n66326, n66327, n66328, n66329, n66330,
         n66331, n66332, n66333, n66334, n66335, n66336, n66337, n66338,
         n66339, n66340, n66341, n66342, n66343, n66344, n66345, n66346,
         n66347, n66348, n66349, n66350, n66351, n66352, n66353, n66354,
         n66355, n66356, n66357, n66358, n66359, n66360, n66361, n66362,
         n66363, n66364, n66365, n66366, n66367, n66368, n66369, n66370,
         n66371, n66372, n66494, n66495, n66496, n66497, n66498, n66499,
         n66500, n66501, n66502, n66503, n66504, n66505, n66506, n66507,
         n66508, n66509, n66510, n66511, n66512, n66513, n66514, n66515,
         n66516, n66517, n66518, n66519, n66520, n66521, n66522, n66523,
         n66524, n66525, n66526, n66527, n66528, n66529, n66530, n66531,
         n66532, n66533, n66534, n66535, n66536, n66537, n66538, n66539,
         n66540, n66541, n66542, n66543, n66544, n66545, n66546, n66547,
         n66548, n66549, n66550, n67260, n67261, n67262, n67263, n67264,
         n67265, n67266, n67267, n67268, n67269, n67270, n67271, n67272,
         n67273, n67274, n67275, n67276, n67277, n67278, n67279, n67280,
         n67281, n67282, n67283, n67284, n67285, n67286, n67287, n67288,
         n67289, n67290, n67291, n67292, n67293, n67294, n67295, n67296,
         n67297, n67298, n67299, n67300, n67301, n67302, n67303, n67304,
         n67305, n67306, n67307, n67308, n67309, n67310, n67311, n67312,
         n67313, n67314, n67315, n67316, n67317, n67318, n67319, n67320,
         n67321, n67322, n67323, n67324, n67325, n67326, n67327, n67328,
         n67329, n67330, n67331, n67332, n67333, n67334, n67335, n67336,
         n67337, n67338, n67339, n67340, n67341, n67342, n67343, n67344,
         n67345, n67346, n67347, n67348, n67349, n67350, n67351, n67352,
         n67353, n67354, n67355, n67356, n67357, n67358, n67359, n67360,
         n67361, n67362, n67363, n67364, n67365, n67366, n67367, n67368,
         n67369, n67370, n67371, n67372, n67373, n67374, n67375, n67376,
         n67377, n67378, n67379, n67380, n67381, n67382, n67383, n67384,
         n67385, n67386, n67387, n67388, n67389, n67390, n67391, n67392,
         n67393, n67394, n67395, n67396, n67397, n67398, n67399, n67400,
         n67401, n67402, n67403, n67404, n67405, n67406, n67407, n67408,
         n67409, n67410, n67411, n67412, n67413, n67414, n67415, n67416,
         n67417, n67418, n67419, n67420, n67421, n67422, n67423, n67424,
         n67425, n67426, n67427, n67428, n67429, n67430, n67431, n67432,
         n67433, n67434, n67435, n67436, n67437, n67438, n67439, n67440,
         n67441, n67442, n67443, n67444, n67445, n67446, n67447, n67448,
         n67449, n67450, n67451, n67452, n67453, n67454, n67455, n67456,
         n67457, n67458, n67459, n67460, n67461, n67462, n67463, n67464,
         n67465, n67466, n67467, n67468, n67469, n67470, n67471, n67472,
         n67473, n67474, n67475, n67476, n67477, n67478, n67479, n67480,
         n67481, n67482, n67483, n67484, n67485, n67486, n67487, n67488,
         n67489, n67490, n67491, n67492, n67493, n67494, n67495, n67496,
         n67497, n67498, n67499, n67500, n67501, n67502, n67503, n67504,
         n67505, n67506, n67507, n67508, n67509, n67510, n67511, n67512,
         n67513, n67514, n67515, n67516, n67517, n67518, n67519, n67520,
         n67521, n67522, n67523, n67524, n67525, n67526, n67527, n67528,
         n67529, n67530, n67531, n67532, n67533, n67534, n67535, n67536,
         n67537, n67538, n67539, n67540, n67541, n67542, n67543, n67544,
         n67545, n67546, n67547, n67548, n67549, n67550, n67551, n67552,
         n67553, n67554, n67555, n67556, n67557, n67558, n67559, n67560,
         n67561, n67562, n67563, n67564, n67565, n67566, n67567, n67568,
         n67569, n67570, n67571, n67572, n67573, n67574, n67575, n67576,
         n67577, n67578, n67579, n67580, n67581, n67582, n67583, n67584,
         n67585, n67586, n67587, n67588, n67589, n67590, n67591, n67592,
         n67593, n67594, n67595, n67596, n67597, n67598, n67599, n67600,
         n67601, n67602, n67603, n67604, n67605, n67606, n67607, n67608,
         n67609, n67610, n67611, n67612, n67613, n67614, n67615, n67616,
         n67617, n67618, n67619, n67620, n67621, n67622, n67623, n67624,
         n67625, n67626, n67627, n67628, n67629, n67630, n67631, n67632,
         n67633, n67634, n67635, n67636, n67637, n67638, n67639, n67640,
         n67641, n67642, n67643, n67644, n67645, n67646, n67647, n67648,
         n67649, n67650, n67651, n67652, n67653, n67654, n67655, n67656,
         n67657, n67658, n67659, n67660, n67661, n67662, n67663, n67664,
         n67665, n67666, n67667, n67668, n67669, n67670, n67671, n67672,
         n67673, n67674, n67675, n67676, n67677, n67678, n67679, n67680,
         n67681, n67682, n67683, n67684, n67685, n67686, n67687, n67688,
         n67689, n67690, n67691, n67692, n67693, n67694, n67695, n67696,
         n67697, n67698, n67699, n67700, n67701, n67702, n67703, n67704,
         n67705, n67706, n67707, n67708, n67709, n67710, n67711, n67712,
         n67713, n67714, n67715, n67716, n67717, n67718, n67719, n67720,
         n67721, n67722, n67723, n67724, n67725, n67726, n67727, n67728,
         n67729, n67730, n67731, n67732, n67733, n67734, n67735, n67736,
         n67737, n67738, n67739, n67740, n67741, n67742, n67743, n67744,
         n67745, n67746, n67747, n67748, n67749, n67750, n67751, n67752,
         n67753, n67754, n67755, n67756, n67757, n67758, n67759, n67760,
         n67761, n67762, n67763, n67764, n67765, n67766, n67767, n67768,
         n67769, n67770, n67771, n67772, n67773, n67774, n67775, n67776,
         n67777, n67778, n67779, n67780, n67781, n67782, n67783, n67784,
         n67785, n67786, n67787, n67788, n67789, n67790, n67791, n67792,
         n67793, n67794, n67795, n67796, n67797, n67798, n67799, n67800,
         n67801, n67802, n67803, n67804, n67805, n67806, n67807, n67808,
         n67809, n67810, n67811, n67812, n67813, n67814, n67815, n67816,
         n67817, n67818, n67819, n67820, n67821, n67822, n67823, n67824,
         n67825, n67826, n67827, n67828, n67829, n67830, n67831, n67832,
         n67833, n67834, n67835, n67836, n67837, n67838, n67839, n67840,
         n67841, n67842, n67843, n67844, n67845, n67846, n67847, n67848,
         n67849, n67850, n67851, n67852, n67853, n67854, n67855, n67856,
         n67857, n67858, n67859, n67860, n67861, n67862, n67863, n67864,
         n67865, n67866, n67867, n67868, n67869, n67870, n67871, n67872,
         n67873, n67874, n67875, n67876, n67877, n67878, n67879, n67880,
         n67881, n67882, n67883, n67884, n67885, n67886, n67887, n67888,
         n67889, n67890, n67891, n67892, n67893, n67894, n67895, n67896,
         n67897, n67898, n67899, n67900, n67901, n67902, n67903, n67904,
         n67905, n67906, n67907, n67908, n67909, n67910, n67911, n67912,
         n67913, n67914, n67915, n67916, n67917, n67918, n67919, n67920,
         n67921, n67922, n67923, n67924, n67925, n67926, n67927, n67928,
         n67929, n67930, n67931, n67932, n67933, n67934, n67935, n67936,
         n67937, n67938, n67939, n67940, n67941, n67942, n67943, n67944,
         n67945, n67946, n67947, n67948, n67949, n67950, n67951, n67952,
         n67953, n67954, n67955, n67956, n67957, n67958, n67959, n67960,
         n67961, n67962, n67963, n67964, n67965, n67966, n67967, n67968,
         n67969, n67970, n67971, n67972, n67973, n67974, n67975, n67976,
         n67977, n67978, n67979, n67980, n67981, n67982, n67983, n67984,
         n67985, n67986, n67987, n67988, n67989, n67990, n67991, n67992,
         n67993, n67994, n67995, n67996, n67997, n67998, n67999, n68000,
         n68001, n68002, n68003, n68004, n68005, n68006, n68007, n68008,
         n68009, n68010, n68011, n68012, n68013, n68014, n68015, n68016,
         n68017, n68018, n68019, n68020, n68021, n68022, n68023, n68024,
         n68025, n68026, n68027, n68028, n68029, n68030, n68031, n68032,
         n68033, n68034, n68035, n68036, n68037, n68038, n68039, n68040,
         n68041, n68042, n68043, n68044, n68045, n68046, n68047, n68048,
         n68049, n68050, n68051, n68052, n68053, n68054, n68055, n68056,
         n68057, n68058, n68059, n68060, n68061, n68062, n68063, n68064,
         n68065, n68066, n68067, n68068, n68069, n68070, n68071, n68072,
         n68073, n68074, n68075, n68076, n68077, n68078, n68079, n68080,
         n68081, n68082, n68083, n68084, n68085, n68086, n68087, n68088,
         n68089, n68090, n68091, n68092, n68093, n68094, n68095, n68096,
         n68097, n68098, n68099, n68100, n68101, n68102, n68103, n68104,
         n68105, n68106, n68107, n68108, n68109, n68110, n68111, n68112,
         n68113, n68114, n68115, n68116, n68117, n68118, n68119, n68120,
         n68121, n68122, n68123, n68124, n68125, n68126, n68127, n68128,
         n68129, n68130, n68131, n68132, n68133, n68134, n68135, n68136,
         n68137, n68138, n68139, n68140, n68141, n68142, n68143, n68144,
         n68145, n68146, n68147, n68148, n68149, n68150, n68151, n68152,
         n68153, n68154, n68155, n68156, n68157, n68158, n68159, n68160,
         n68161, n68162, n68163, n68164, n68165, n68166, n68167, n68168,
         n68169, n68170, n68171, n68172, n68173, n68174, n68175, n68176,
         n68177, n68178, n68179, n68180, n68181, n68182, n68183, n68184,
         n68185, n68186, n68187, n68188, n68189, n68190, n68191, n68192,
         n68193, n68194, n68195, n68196, n68197, n68198, n68199, n68200,
         n68201, n68202, n68203, n68204, n68205, n68206, n68207, n68208,
         n68209, n68210, n68211, n68212, n68213, n68214, n68215, n68216,
         n68217, n68218, n68219, n68220, n68221, n68222, n68223, n68224,
         n68225, n68226, n68227, n68228, n68229, n68230, n68231, n68232,
         n68233, n68234, n68235, n68236, n68237, n68238, n68239, n68240,
         n68241, n68242, n68243, n68244, n68245, n68246, n68247, n68248,
         n68249, n68250, n68251, n68252, n68253, n68254, n68255, n68256,
         n68257, n68258, n68259, n68260, n68261, n68262;

  DFF_X1 \OUT1_reg[59]  ( .D(n5493), .CK(CLK), .Q(OUT1[59]) );
  DFF_X1 \OUT1_reg[58]  ( .D(n5491), .CK(CLK), .Q(OUT1[58]) );
  DFF_X1 \OUT1_reg[57]  ( .D(n5489), .CK(CLK), .Q(OUT1[57]) );
  DFF_X1 \OUT1_reg[56]  ( .D(n5487), .CK(CLK), .Q(OUT1[56]) );
  DFF_X1 \OUT1_reg[55]  ( .D(n5485), .CK(CLK), .Q(OUT1[55]) );
  DFF_X1 \OUT1_reg[54]  ( .D(n5483), .CK(CLK), .Q(OUT1[54]) );
  DFF_X1 \OUT1_reg[53]  ( .D(n5481), .CK(CLK), .Q(OUT1[53]) );
  DFF_X1 \OUT1_reg[52]  ( .D(n5479), .CK(CLK), .Q(OUT1[52]) );
  DFF_X1 \OUT1_reg[51]  ( .D(n5477), .CK(CLK), .Q(OUT1[51]) );
  DFF_X1 \OUT1_reg[50]  ( .D(n5475), .CK(CLK), .Q(OUT1[50]) );
  DFF_X1 \OUT1_reg[49]  ( .D(n5473), .CK(CLK), .Q(OUT1[49]) );
  DFF_X1 \OUT1_reg[48]  ( .D(n5471), .CK(CLK), .Q(OUT1[48]) );
  DFF_X1 \OUT1_reg[47]  ( .D(n5469), .CK(CLK), .Q(OUT1[47]) );
  DFF_X1 \OUT1_reg[46]  ( .D(n5467), .CK(CLK), .Q(OUT1[46]) );
  DFF_X1 \OUT1_reg[45]  ( .D(n5465), .CK(CLK), .Q(OUT1[45]) );
  DFF_X1 \OUT1_reg[44]  ( .D(n5463), .CK(CLK), .Q(OUT1[44]) );
  DFF_X1 \OUT1_reg[43]  ( .D(n5461), .CK(CLK), .Q(OUT1[43]) );
  DFF_X1 \OUT1_reg[42]  ( .D(n5459), .CK(CLK), .Q(OUT1[42]) );
  DFF_X1 \OUT1_reg[41]  ( .D(n5457), .CK(CLK), .Q(OUT1[41]) );
  DFF_X1 \OUT1_reg[40]  ( .D(n5455), .CK(CLK), .Q(OUT1[40]) );
  DFF_X1 \OUT1_reg[39]  ( .D(n5453), .CK(CLK), .Q(OUT1[39]) );
  DFF_X1 \OUT1_reg[38]  ( .D(n5451), .CK(CLK), .Q(OUT1[38]) );
  DFF_X1 \OUT1_reg[37]  ( .D(n5449), .CK(CLK), .Q(OUT1[37]) );
  DFF_X1 \OUT1_reg[36]  ( .D(n5447), .CK(CLK), .Q(OUT1[36]) );
  DFF_X1 \OUT1_reg[35]  ( .D(n5445), .CK(CLK), .Q(OUT1[35]) );
  DFF_X1 \OUT1_reg[34]  ( .D(n5443), .CK(CLK), .Q(OUT1[34]) );
  DFF_X1 \OUT1_reg[33]  ( .D(n5441), .CK(CLK), .Q(OUT1[33]) );
  DFF_X1 \OUT1_reg[32]  ( .D(n5439), .CK(CLK), .Q(OUT1[32]) );
  DFF_X1 \OUT1_reg[31]  ( .D(n5437), .CK(CLK), .Q(OUT1[31]) );
  DFF_X1 \OUT1_reg[30]  ( .D(n5435), .CK(CLK), .Q(OUT1[30]) );
  DFF_X1 \OUT1_reg[29]  ( .D(n5433), .CK(CLK), .Q(OUT1[29]) );
  DFF_X1 \OUT1_reg[28]  ( .D(n5431), .CK(CLK), .Q(OUT1[28]) );
  DFF_X1 \OUT1_reg[27]  ( .D(n5429), .CK(CLK), .Q(OUT1[27]) );
  DFF_X1 \OUT1_reg[26]  ( .D(n5427), .CK(CLK), .Q(OUT1[26]) );
  DFF_X1 \OUT1_reg[25]  ( .D(n5425), .CK(CLK), .Q(OUT1[25]) );
  DFF_X1 \OUT1_reg[24]  ( .D(n5423), .CK(CLK), .Q(OUT1[24]) );
  DFF_X1 \OUT1_reg[23]  ( .D(n5421), .CK(CLK), .Q(OUT1[23]) );
  DFF_X1 \OUT1_reg[22]  ( .D(n5419), .CK(CLK), .Q(OUT1[22]) );
  DFF_X1 \OUT1_reg[21]  ( .D(n5417), .CK(CLK), .Q(OUT1[21]) );
  DFF_X1 \OUT1_reg[20]  ( .D(n5415), .CK(CLK), .Q(OUT1[20]) );
  DFF_X1 \OUT1_reg[19]  ( .D(n5413), .CK(CLK), .Q(OUT1[19]) );
  DFF_X1 \OUT1_reg[18]  ( .D(n5411), .CK(CLK), .Q(OUT1[18]) );
  DFF_X1 \OUT1_reg[17]  ( .D(n5409), .CK(CLK), .Q(OUT1[17]) );
  DFF_X1 \OUT1_reg[16]  ( .D(n5407), .CK(CLK), .Q(OUT1[16]) );
  DFF_X1 \OUT1_reg[15]  ( .D(n5405), .CK(CLK), .Q(OUT1[15]) );
  DFF_X1 \OUT1_reg[14]  ( .D(n5403), .CK(CLK), .Q(OUT1[14]) );
  DFF_X1 \OUT1_reg[13]  ( .D(n5401), .CK(CLK), .Q(OUT1[13]) );
  DFF_X1 \OUT1_reg[12]  ( .D(n5399), .CK(CLK), .Q(OUT1[12]) );
  DFF_X1 \OUT1_reg[11]  ( .D(n5397), .CK(CLK), .Q(OUT1[11]) );
  DFF_X1 \OUT1_reg[10]  ( .D(n5395), .CK(CLK), .Q(OUT1[10]) );
  DFF_X1 \OUT1_reg[9]  ( .D(n5393), .CK(CLK), .Q(OUT1[9]) );
  DFF_X1 \OUT1_reg[8]  ( .D(n5391), .CK(CLK), .Q(OUT1[8]) );
  DFF_X1 \OUT1_reg[7]  ( .D(n5389), .CK(CLK), .Q(OUT1[7]) );
  DFF_X1 \OUT1_reg[6]  ( .D(n5387), .CK(CLK), .Q(OUT1[6]) );
  DFF_X1 \OUT1_reg[5]  ( .D(n5385), .CK(CLK), .Q(OUT1[5]) );
  DFF_X1 \OUT1_reg[4]  ( .D(n5383), .CK(CLK), .Q(OUT1[4]) );
  DFF_X1 \OUT1_reg[3]  ( .D(n5381), .CK(CLK), .Q(OUT1[3]) );
  DFF_X1 \OUT1_reg[2]  ( .D(n5379), .CK(CLK), .Q(OUT1[2]) );
  DFF_X1 \OUT1_reg[1]  ( .D(n5377), .CK(CLK), .Q(OUT1[1]) );
  DFF_X1 \OUT1_reg[0]  ( .D(n5375), .CK(CLK), .Q(OUT1[0]) );
  DFF_X1 \OUT2_reg[61]  ( .D(n5372), .CK(CLK), .Q(OUT2[61]) );
  DFF_X1 \OUT2_reg[60]  ( .D(n5371), .CK(CLK), .Q(OUT2[60]) );
  DFF_X1 \OUT2_reg[59]  ( .D(n5370), .CK(CLK), .Q(OUT2[59]) );
  DFF_X1 \OUT2_reg[58]  ( .D(n5369), .CK(CLK), .Q(OUT2[58]) );
  DFF_X1 \OUT2_reg[57]  ( .D(n5368), .CK(CLK), .Q(OUT2[57]) );
  DFF_X1 \OUT2_reg[56]  ( .D(n5367), .CK(CLK), .Q(OUT2[56]) );
  DFF_X1 \OUT2_reg[55]  ( .D(n5366), .CK(CLK), .Q(OUT2[55]) );
  DFF_X1 \OUT2_reg[54]  ( .D(n5365), .CK(CLK), .Q(OUT2[54]) );
  DFF_X1 \OUT2_reg[53]  ( .D(n5364), .CK(CLK), .Q(OUT2[53]) );
  DFF_X1 \OUT2_reg[52]  ( .D(n5363), .CK(CLK), .Q(OUT2[52]) );
  DFF_X1 \OUT2_reg[51]  ( .D(n5362), .CK(CLK), .Q(OUT2[51]) );
  DFF_X1 \OUT2_reg[50]  ( .D(n5361), .CK(CLK), .Q(OUT2[50]) );
  DFF_X1 \OUT2_reg[49]  ( .D(n5360), .CK(CLK), .Q(OUT2[49]) );
  DFF_X1 \OUT2_reg[48]  ( .D(n5359), .CK(CLK), .Q(OUT2[48]) );
  DFF_X1 \OUT2_reg[47]  ( .D(n5358), .CK(CLK), .Q(OUT2[47]) );
  DFF_X1 \OUT2_reg[46]  ( .D(n5357), .CK(CLK), .Q(OUT2[46]) );
  DFF_X1 \OUT2_reg[45]  ( .D(n5356), .CK(CLK), .Q(OUT2[45]) );
  DFF_X1 \OUT2_reg[44]  ( .D(n5355), .CK(CLK), .Q(OUT2[44]) );
  DFF_X1 \OUT2_reg[43]  ( .D(n5354), .CK(CLK), .Q(OUT2[43]) );
  DFF_X1 \OUT2_reg[42]  ( .D(n5353), .CK(CLK), .Q(OUT2[42]) );
  DFF_X1 \OUT2_reg[41]  ( .D(n5352), .CK(CLK), .Q(OUT2[41]) );
  DFF_X1 \OUT2_reg[40]  ( .D(n5351), .CK(CLK), .Q(OUT2[40]) );
  DFF_X1 \OUT2_reg[39]  ( .D(n5350), .CK(CLK), .Q(OUT2[39]) );
  DFF_X1 \OUT2_reg[38]  ( .D(n5349), .CK(CLK), .Q(OUT2[38]) );
  DFF_X1 \OUT2_reg[37]  ( .D(n5348), .CK(CLK), .Q(OUT2[37]) );
  DFF_X1 \OUT2_reg[36]  ( .D(n5347), .CK(CLK), .Q(OUT2[36]) );
  DFF_X1 \OUT2_reg[35]  ( .D(n5346), .CK(CLK), .Q(OUT2[35]) );
  DFF_X1 \OUT2_reg[34]  ( .D(n5345), .CK(CLK), .Q(OUT2[34]) );
  DFF_X1 \OUT2_reg[33]  ( .D(n5344), .CK(CLK), .Q(OUT2[33]) );
  DFF_X1 \OUT2_reg[32]  ( .D(n5343), .CK(CLK), .Q(OUT2[32]) );
  DFF_X1 \OUT2_reg[31]  ( .D(n5342), .CK(CLK), .Q(OUT2[31]) );
  DFF_X1 \OUT2_reg[30]  ( .D(n5341), .CK(CLK), .Q(OUT2[30]) );
  DFF_X1 \OUT2_reg[29]  ( .D(n5340), .CK(CLK), .Q(OUT2[29]) );
  DFF_X1 \OUT2_reg[28]  ( .D(n5339), .CK(CLK), .Q(OUT2[28]) );
  DFF_X1 \OUT2_reg[27]  ( .D(n5338), .CK(CLK), .Q(OUT2[27]) );
  DFF_X1 \OUT2_reg[26]  ( .D(n5337), .CK(CLK), .Q(OUT2[26]) );
  DFF_X1 \OUT2_reg[25]  ( .D(n5336), .CK(CLK), .Q(OUT2[25]) );
  DFF_X1 \OUT2_reg[24]  ( .D(n5335), .CK(CLK), .Q(OUT2[24]) );
  DFF_X1 \OUT2_reg[23]  ( .D(n5334), .CK(CLK), .Q(OUT2[23]) );
  DFF_X1 \OUT2_reg[22]  ( .D(n5333), .CK(CLK), .Q(OUT2[22]) );
  DFF_X1 \OUT2_reg[21]  ( .D(n5332), .CK(CLK), .Q(OUT2[21]) );
  DFF_X1 \OUT2_reg[20]  ( .D(n5331), .CK(CLK), .Q(OUT2[20]) );
  DFF_X1 \OUT2_reg[19]  ( .D(n5330), .CK(CLK), .Q(OUT2[19]) );
  DFF_X1 \OUT2_reg[18]  ( .D(n5329), .CK(CLK), .Q(OUT2[18]) );
  DFF_X1 \OUT2_reg[17]  ( .D(n5328), .CK(CLK), .Q(OUT2[17]) );
  DFF_X1 \OUT2_reg[16]  ( .D(n5327), .CK(CLK), .Q(OUT2[16]) );
  DFF_X1 \OUT2_reg[15]  ( .D(n5326), .CK(CLK), .Q(OUT2[15]) );
  DFF_X1 \OUT2_reg[14]  ( .D(n5325), .CK(CLK), .Q(OUT2[14]) );
  DFF_X1 \OUT2_reg[13]  ( .D(n5324), .CK(CLK), .Q(OUT2[13]) );
  DFF_X1 \OUT2_reg[12]  ( .D(n5323), .CK(CLK), .Q(OUT2[12]) );
  DFF_X1 \OUT2_reg[11]  ( .D(n5322), .CK(CLK), .Q(OUT2[11]) );
  DFF_X1 \OUT2_reg[10]  ( .D(n5321), .CK(CLK), .Q(OUT2[10]) );
  DFF_X1 \OUT2_reg[9]  ( .D(n5320), .CK(CLK), .Q(OUT2[9]) );
  DFF_X1 \OUT2_reg[8]  ( .D(n5319), .CK(CLK), .Q(OUT2[8]) );
  DFF_X1 \OUT2_reg[7]  ( .D(n5318), .CK(CLK), .Q(OUT2[7]) );
  DFF_X1 \OUT2_reg[6]  ( .D(n5317), .CK(CLK), .Q(OUT2[6]) );
  DFF_X1 \OUT2_reg[5]  ( .D(n5316), .CK(CLK), .Q(OUT2[5]) );
  DFF_X1 \OUT2_reg[4]  ( .D(n5315), .CK(CLK), .Q(OUT2[4]) );
  DFF_X1 \OUT2_reg[3]  ( .D(n5314), .CK(CLK), .Q(OUT2[3]) );
  DFF_X1 \OUT2_reg[2]  ( .D(n5313), .CK(CLK), .Q(OUT2[2]) );
  DFF_X1 \OUT2_reg[1]  ( .D(n5312), .CK(CLK), .Q(OUT2[1]) );
  DFF_X1 \OUT2_reg[0]  ( .D(n5311), .CK(CLK), .Q(OUT2[0]) );
  DFF_X1 \REGISTERS_reg[21][63]  ( .D(n6142), .CK(CLK), .Q(n58960), .QN(n8497)
         );
  DFF_X1 \REGISTERS_reg[21][62]  ( .D(n6141), .CK(CLK), .Q(n59026), .QN(n8481)
         );
  DFF_X1 \REGISTERS_reg[21][61]  ( .D(n6140), .CK(CLK), .Q(n59024), .QN(n8465)
         );
  DFF_X1 \REGISTERS_reg[21][60]  ( .D(n6139), .CK(CLK), .Q(n59022), .QN(n8449)
         );
  DFF_X1 \REGISTERS_reg[18][63]  ( .D(n6334), .CK(CLK), .QN(n49483) );
  DFF_X1 \REGISTERS_reg[18][62]  ( .D(n6333), .CK(CLK), .QN(n49482) );
  DFF_X1 \REGISTERS_reg[18][61]  ( .D(n6332), .CK(CLK), .QN(n49481) );
  DFF_X1 \REGISTERS_reg[18][60]  ( .D(n6331), .CK(CLK), .QN(n49480) );
  DFF_X1 \REGISTERS_reg[21][59]  ( .D(n6138), .CK(CLK), .Q(n56611), .QN(n8433)
         );
  DFF_X1 \REGISTERS_reg[21][58]  ( .D(n6137), .CK(CLK), .Q(n56635), .QN(n8417)
         );
  DFF_X1 \REGISTERS_reg[21][57]  ( .D(n6136), .CK(CLK), .Q(n56659), .QN(n8401)
         );
  DFF_X1 \REGISTERS_reg[21][56]  ( .D(n6135), .CK(CLK), .Q(n56683), .QN(n8385)
         );
  DFF_X1 \REGISTERS_reg[21][55]  ( .D(n6134), .CK(CLK), .Q(n56707), .QN(n8369)
         );
  DFF_X1 \REGISTERS_reg[21][54]  ( .D(n6133), .CK(CLK), .Q(n56731), .QN(n8353)
         );
  DFF_X1 \REGISTERS_reg[21][53]  ( .D(n6132), .CK(CLK), .Q(n56755), .QN(n8337)
         );
  DFF_X1 \REGISTERS_reg[21][52]  ( .D(n6131), .CK(CLK), .Q(n56779), .QN(n8321)
         );
  DFF_X1 \REGISTERS_reg[21][51]  ( .D(n6130), .CK(CLK), .Q(n56803), .QN(n8305)
         );
  DFF_X1 \REGISTERS_reg[21][50]  ( .D(n6129), .CK(CLK), .Q(n56827), .QN(n8289)
         );
  DFF_X1 \REGISTERS_reg[21][49]  ( .D(n6128), .CK(CLK), .Q(n56851), .QN(n8273)
         );
  DFF_X1 \REGISTERS_reg[21][48]  ( .D(n6127), .CK(CLK), .Q(n56875), .QN(n8257)
         );
  DFF_X1 \REGISTERS_reg[21][47]  ( .D(n6126), .CK(CLK), .Q(n56899), .QN(n8241)
         );
  DFF_X1 \REGISTERS_reg[21][46]  ( .D(n6125), .CK(CLK), .Q(n56923), .QN(n8225)
         );
  DFF_X1 \REGISTERS_reg[21][45]  ( .D(n6124), .CK(CLK), .Q(n56947), .QN(n8209)
         );
  DFF_X1 \REGISTERS_reg[21][44]  ( .D(n6123), .CK(CLK), .Q(n56971), .QN(n8193)
         );
  DFF_X1 \REGISTERS_reg[21][43]  ( .D(n6122), .CK(CLK), .Q(n56995), .QN(n8177)
         );
  DFF_X1 \REGISTERS_reg[21][42]  ( .D(n6121), .CK(CLK), .Q(n57019), .QN(n8161)
         );
  DFF_X1 \REGISTERS_reg[21][41]  ( .D(n6120), .CK(CLK), .Q(n57043), .QN(n8145)
         );
  DFF_X1 \REGISTERS_reg[21][40]  ( .D(n6119), .CK(CLK), .Q(n57067), .QN(n8129)
         );
  DFF_X1 \REGISTERS_reg[21][39]  ( .D(n6118), .CK(CLK), .Q(n57091), .QN(n8113)
         );
  DFF_X1 \REGISTERS_reg[21][38]  ( .D(n6117), .CK(CLK), .Q(n57115), .QN(n8097)
         );
  DFF_X1 \REGISTERS_reg[21][37]  ( .D(n6116), .CK(CLK), .Q(n57139), .QN(n8081)
         );
  DFF_X1 \REGISTERS_reg[21][36]  ( .D(n6115), .CK(CLK), .Q(n57163), .QN(n8065)
         );
  DFF_X1 \REGISTERS_reg[21][35]  ( .D(n6114), .CK(CLK), .Q(n57187), .QN(n8049)
         );
  DFF_X1 \REGISTERS_reg[21][34]  ( .D(n6113), .CK(CLK), .Q(n57211), .QN(n8033)
         );
  DFF_X1 \REGISTERS_reg[21][33]  ( .D(n6112), .CK(CLK), .Q(n57235), .QN(n8017)
         );
  DFF_X1 \REGISTERS_reg[21][32]  ( .D(n6111), .CK(CLK), .Q(n57259), .QN(n8001)
         );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n6110), .CK(CLK), .Q(n57283), .QN(n7985)
         );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n6109), .CK(CLK), .Q(n57307), .QN(n7969)
         );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n6108), .CK(CLK), .Q(n57331), .QN(n7953)
         );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n6107), .CK(CLK), .Q(n57355), .QN(n7937)
         );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n6106), .CK(CLK), .Q(n57379), .QN(n7921)
         );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n6105), .CK(CLK), .Q(n57403), .QN(n7905)
         );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n6104), .CK(CLK), .Q(n57427), .QN(n7889)
         );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n6103), .CK(CLK), .Q(n57451), .QN(n7873)
         );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n6102), .CK(CLK), .Q(n57475), .QN(n7857)
         );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n6101), .CK(CLK), .Q(n57499), .QN(n7841)
         );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n6100), .CK(CLK), .Q(n57523), .QN(n7825)
         );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n6099), .CK(CLK), .Q(n57547), .QN(n7809)
         );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n6098), .CK(CLK), .Q(n57571), .QN(n7793)
         );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n6097), .CK(CLK), .Q(n57595), .QN(n7777)
         );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n6096), .CK(CLK), .Q(n57619), .QN(n7761)
         );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n6095), .CK(CLK), .Q(n57643), .QN(n7745)
         );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n6094), .CK(CLK), .Q(n57667), .QN(n7729)
         );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n6093), .CK(CLK), .Q(n57691), .QN(n7713)
         );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n6092), .CK(CLK), .Q(n57715), .QN(n7697)
         );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n6091), .CK(CLK), .Q(n57739), .QN(n7681)
         );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n6090), .CK(CLK), .Q(n57763), .QN(n7665)
         );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n6089), .CK(CLK), .Q(n57787), .QN(n7649)
         );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n6088), .CK(CLK), .Q(n57811), .QN(n7633)
         );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n6087), .CK(CLK), .Q(n57835), .QN(n7617)
         );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n6086), .CK(CLK), .Q(n57859), .QN(n7601)
         );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n6085), .CK(CLK), .Q(n57883), .QN(n7585)
         );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n6084), .CK(CLK), .Q(n57907), .QN(n7569)
         );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n6083), .CK(CLK), .Q(n57931), .QN(n7553)
         );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n6082), .CK(CLK), .Q(n57955), .QN(n7537)
         );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n6081), .CK(CLK), .Q(n57979), .QN(n7521)
         );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n6080), .CK(CLK), .Q(n58003), .QN(n7505)
         );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n6079), .CK(CLK), .Q(n58041), .QN(n7489)
         );
  DFF_X1 \REGISTERS_reg[18][59]  ( .D(n6330), .CK(CLK), .QN(n49479) );
  DFF_X1 \REGISTERS_reg[18][58]  ( .D(n6329), .CK(CLK), .QN(n49478) );
  DFF_X1 \REGISTERS_reg[18][57]  ( .D(n6328), .CK(CLK), .QN(n49477) );
  DFF_X1 \REGISTERS_reg[18][56]  ( .D(n6327), .CK(CLK), .QN(n49476) );
  DFF_X1 \REGISTERS_reg[18][55]  ( .D(n6326), .CK(CLK), .QN(n49475) );
  DFF_X1 \REGISTERS_reg[18][54]  ( .D(n6325), .CK(CLK), .QN(n49474) );
  DFF_X1 \REGISTERS_reg[18][53]  ( .D(n6324), .CK(CLK), .QN(n49473) );
  DFF_X1 \REGISTERS_reg[18][52]  ( .D(n6323), .CK(CLK), .QN(n49472) );
  DFF_X1 \REGISTERS_reg[18][51]  ( .D(n6322), .CK(CLK), .QN(n49471) );
  DFF_X1 \REGISTERS_reg[18][50]  ( .D(n6321), .CK(CLK), .QN(n49470) );
  DFF_X1 \REGISTERS_reg[18][49]  ( .D(n6320), .CK(CLK), .QN(n49469) );
  DFF_X1 \REGISTERS_reg[18][48]  ( .D(n6319), .CK(CLK), .QN(n49468) );
  DFF_X1 \REGISTERS_reg[18][47]  ( .D(n6318), .CK(CLK), .QN(n49467) );
  DFF_X1 \REGISTERS_reg[18][46]  ( .D(n6317), .CK(CLK), .QN(n49466) );
  DFF_X1 \REGISTERS_reg[18][45]  ( .D(n6316), .CK(CLK), .QN(n49465) );
  DFF_X1 \REGISTERS_reg[18][44]  ( .D(n6315), .CK(CLK), .QN(n49464) );
  DFF_X1 \REGISTERS_reg[18][43]  ( .D(n6314), .CK(CLK), .QN(n49463) );
  DFF_X1 \REGISTERS_reg[18][42]  ( .D(n6313), .CK(CLK), .QN(n49462) );
  DFF_X1 \REGISTERS_reg[18][41]  ( .D(n6312), .CK(CLK), .QN(n49461) );
  DFF_X1 \REGISTERS_reg[18][40]  ( .D(n6311), .CK(CLK), .QN(n49460) );
  DFF_X1 \REGISTERS_reg[18][39]  ( .D(n6310), .CK(CLK), .QN(n49459) );
  DFF_X1 \REGISTERS_reg[18][38]  ( .D(n6309), .CK(CLK), .QN(n49458) );
  DFF_X1 \REGISTERS_reg[18][37]  ( .D(n6308), .CK(CLK), .QN(n49457) );
  DFF_X1 \REGISTERS_reg[18][36]  ( .D(n6307), .CK(CLK), .QN(n49456) );
  DFF_X1 \REGISTERS_reg[18][35]  ( .D(n6306), .CK(CLK), .QN(n49455) );
  DFF_X1 \REGISTERS_reg[18][34]  ( .D(n6305), .CK(CLK), .QN(n49454) );
  DFF_X1 \REGISTERS_reg[18][33]  ( .D(n6304), .CK(CLK), .QN(n49453) );
  DFF_X1 \REGISTERS_reg[18][32]  ( .D(n6303), .CK(CLK), .QN(n49452) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n6302), .CK(CLK), .QN(n49451) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n6301), .CK(CLK), .QN(n49450) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n6300), .CK(CLK), .QN(n49449) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n6299), .CK(CLK), .QN(n49448) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n6298), .CK(CLK), .QN(n49447) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n6297), .CK(CLK), .QN(n49446) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n6296), .CK(CLK), .QN(n49445) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n6295), .CK(CLK), .QN(n49444) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n6294), .CK(CLK), .QN(n49443) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n6293), .CK(CLK), .QN(n49442) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n6292), .CK(CLK), .QN(n49441) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n6291), .CK(CLK), .QN(n49440) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n6290), .CK(CLK), .QN(n49439) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n6289), .CK(CLK), .QN(n49438) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n6288), .CK(CLK), .QN(n49437) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n6287), .CK(CLK), .QN(n49436) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n6286), .CK(CLK), .QN(n49435) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n6285), .CK(CLK), .QN(n49434) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n6284), .CK(CLK), .QN(n49433) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n6283), .CK(CLK), .QN(n49432) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n6282), .CK(CLK), .QN(n49431) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n6281), .CK(CLK), .QN(n49430) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n6280), .CK(CLK), .QN(n49429) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n6279), .CK(CLK), .QN(n49428) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n6278), .CK(CLK), .QN(n49427) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n6277), .CK(CLK), .QN(n49426) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n6276), .CK(CLK), .QN(n49425) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n6275), .CK(CLK), .QN(n49424) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n6274), .CK(CLK), .QN(n49423) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n6273), .CK(CLK), .QN(n49422) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n6272), .CK(CLK), .QN(n49421) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n6271), .CK(CLK), .QN(n49420) );
  DFF_X1 \REGISTERS_reg[13][63]  ( .D(n6654), .CK(CLK), .Q(n66498), .QN(n8509)
         );
  DFF_X1 \REGISTERS_reg[13][62]  ( .D(n6653), .CK(CLK), .Q(n66497), .QN(n8493)
         );
  DFF_X1 \REGISTERS_reg[13][61]  ( .D(n6652), .CK(CLK), .Q(n66496), .QN(n8477)
         );
  DFF_X1 \REGISTERS_reg[13][60]  ( .D(n6651), .CK(CLK), .Q(n66495), .QN(n8461)
         );
  DFF_X1 \REGISTERS_reg[12][63]  ( .D(n6718), .CK(CLK), .Q(n66550), .QN(n49228) );
  DFF_X1 \REGISTERS_reg[12][62]  ( .D(n6717), .CK(CLK), .Q(n66501), .QN(n49231) );
  DFF_X1 \REGISTERS_reg[12][61]  ( .D(n6716), .CK(CLK), .Q(n66500), .QN(n49230) );
  DFF_X1 \REGISTERS_reg[12][60]  ( .D(n6715), .CK(CLK), .Q(n66499), .QN(n49229) );
  DFF_X1 \REGISTERS_reg[12][59]  ( .D(n6714), .CK(CLK), .Q(n66513), .QN(n49291) );
  DFF_X1 \REGISTERS_reg[12][58]  ( .D(n6713), .CK(CLK), .Q(n66512), .QN(n49290) );
  DFF_X1 \REGISTERS_reg[12][57]  ( .D(n6712), .CK(CLK), .Q(n66511), .QN(n49289) );
  DFF_X1 \REGISTERS_reg[12][56]  ( .D(n6711), .CK(CLK), .Q(n66510), .QN(n49288) );
  DFF_X1 \REGISTERS_reg[12][55]  ( .D(n6710), .CK(CLK), .Q(n66509), .QN(n49287) );
  DFF_X1 \REGISTERS_reg[12][54]  ( .D(n6709), .CK(CLK), .Q(n66508), .QN(n49286) );
  DFF_X1 \REGISTERS_reg[12][53]  ( .D(n6708), .CK(CLK), .Q(n66507), .QN(n49285) );
  DFF_X1 \REGISTERS_reg[12][52]  ( .D(n6707), .CK(CLK), .Q(n66506), .QN(n49284) );
  DFF_X1 \REGISTERS_reg[12][51]  ( .D(n6706), .CK(CLK), .Q(n66505), .QN(n49283) );
  DFF_X1 \REGISTERS_reg[12][50]  ( .D(n6705), .CK(CLK), .Q(n66504), .QN(n49282) );
  DFF_X1 \REGISTERS_reg[12][49]  ( .D(n6704), .CK(CLK), .Q(n66503), .QN(n49281) );
  DFF_X1 \REGISTERS_reg[12][48]  ( .D(n6703), .CK(CLK), .Q(n66502), .QN(n49280) );
  DFF_X1 \REGISTERS_reg[12][47]  ( .D(n6702), .CK(CLK), .Q(n66549), .QN(n49279) );
  DFF_X1 \REGISTERS_reg[12][46]  ( .D(n6701), .CK(CLK), .Q(n66548), .QN(n49278) );
  DFF_X1 \REGISTERS_reg[12][45]  ( .D(n6700), .CK(CLK), .Q(n66547), .QN(n49277) );
  DFF_X1 \REGISTERS_reg[12][44]  ( .D(n6699), .CK(CLK), .Q(n66546), .QN(n49276) );
  DFF_X1 \REGISTERS_reg[12][43]  ( .D(n6698), .CK(CLK), .Q(n66545), .QN(n49275) );
  DFF_X1 \REGISTERS_reg[12][42]  ( .D(n6697), .CK(CLK), .Q(n66544), .QN(n49274) );
  DFF_X1 \REGISTERS_reg[12][41]  ( .D(n6696), .CK(CLK), .Q(n66543), .QN(n49273) );
  DFF_X1 \REGISTERS_reg[12][40]  ( .D(n6695), .CK(CLK), .Q(n66542), .QN(n49272) );
  DFF_X1 \REGISTERS_reg[12][39]  ( .D(n6694), .CK(CLK), .Q(n66541), .QN(n49271) );
  DFF_X1 \REGISTERS_reg[12][38]  ( .D(n6693), .CK(CLK), .Q(n66540), .QN(n49270) );
  DFF_X1 \REGISTERS_reg[12][37]  ( .D(n6692), .CK(CLK), .Q(n66539), .QN(n49269) );
  DFF_X1 \REGISTERS_reg[12][36]  ( .D(n6691), .CK(CLK), .Q(n66538), .QN(n49268) );
  DFF_X1 \REGISTERS_reg[12][35]  ( .D(n6690), .CK(CLK), .Q(n66537), .QN(n49267) );
  DFF_X1 \REGISTERS_reg[12][34]  ( .D(n6689), .CK(CLK), .Q(n66536), .QN(n49266) );
  DFF_X1 \REGISTERS_reg[12][33]  ( .D(n6688), .CK(CLK), .Q(n66535), .QN(n49265) );
  DFF_X1 \REGISTERS_reg[12][32]  ( .D(n6687), .CK(CLK), .Q(n66534), .QN(n49264) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n6686), .CK(CLK), .Q(n66533), .QN(n49263) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n6685), .CK(CLK), .Q(n66532), .QN(n49262) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n6684), .CK(CLK), .Q(n66531), .QN(n49261) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n6683), .CK(CLK), .Q(n66530), .QN(n49260) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n6682), .CK(CLK), .Q(n66529), .QN(n49259) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n6681), .CK(CLK), .Q(n66528), .QN(n49258) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n6680), .CK(CLK), .Q(n66527), .QN(n49257) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n6679), .CK(CLK), .Q(n66526), .QN(n49256) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n6678), .CK(CLK), .Q(n66525), .QN(n49255) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n6677), .CK(CLK), .Q(n66524), .QN(n49254) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n6676), .CK(CLK), .Q(n66523), .QN(n49253) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n6675), .CK(CLK), .Q(n66522), .QN(n49252) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n6674), .CK(CLK), .Q(n66521), .QN(n49251) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n6673), .CK(CLK), .Q(n66520), .QN(n49250) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n6672), .CK(CLK), .Q(n66519), .QN(n49249) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n6671), .CK(CLK), .Q(n66518), .QN(n49248) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n6670), .CK(CLK), .Q(n66517), .QN(n49247) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n6669), .CK(CLK), .Q(n66516), .QN(n49246) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n6668), .CK(CLK), .Q(n66515), .QN(n49245) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n6667), .CK(CLK), .Q(n66514), .QN(n49244) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n6666), .CK(CLK), .Q(n64855), .QN(n49243) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n6665), .CK(CLK), .Q(n64875), .QN(n49242) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n6664), .CK(CLK), .Q(n64895), .QN(n49241)
         );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n6663), .CK(CLK), .Q(n64915), .QN(n49240)
         );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n6662), .CK(CLK), .Q(n64935), .QN(n49239)
         );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n6661), .CK(CLK), .Q(n64955), .QN(n49238)
         );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n6660), .CK(CLK), .Q(n64975), .QN(n49237)
         );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n6659), .CK(CLK), .Q(n64995), .QN(n49236)
         );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n6658), .CK(CLK), .Q(n65015), .QN(n49235)
         );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n6657), .CK(CLK), .Q(n65035), .QN(n49234)
         );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n6656), .CK(CLK), .Q(n65055), .QN(n49233)
         );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n6655), .CK(CLK), .Q(n65084), .QN(n49232)
         );
  DFF_X1 \REGISTERS_reg[26][63]  ( .D(n5822), .CK(CLK), .Q(n50647), .QN(n54606) );
  DFF_X1 \REGISTERS_reg[26][62]  ( .D(n5821), .CK(CLK), .Q(n50646), .QN(n54608) );
  DFF_X1 \REGISTERS_reg[26][61]  ( .D(n5820), .CK(CLK), .Q(n50645), .QN(n54609) );
  DFF_X1 \REGISTERS_reg[26][60]  ( .D(n5819), .CK(CLK), .Q(n50644), .QN(n54610) );
  DFF_X1 \REGISTERS_reg[10][62]  ( .D(n6845), .CK(CLK), .Q(n50579), .QN(n54184) );
  DFF_X1 \REGISTERS_reg[10][61]  ( .D(n6844), .CK(CLK), .Q(n50578), .QN(n54185) );
  DFF_X1 \REGISTERS_reg[10][60]  ( .D(n6843), .CK(CLK), .Q(n50577), .QN(n54186) );
  DFF_X1 \REGISTERS_reg[26][59]  ( .D(n5818), .CK(CLK), .Q(n50707), .QN(n54611) );
  DFF_X1 \REGISTERS_reg[26][58]  ( .D(n5817), .CK(CLK), .Q(n50706), .QN(n54612) );
  DFF_X1 \REGISTERS_reg[26][57]  ( .D(n5816), .CK(CLK), .Q(n50705), .QN(n54613) );
  DFF_X1 \REGISTERS_reg[26][56]  ( .D(n5815), .CK(CLK), .Q(n50704), .QN(n54614) );
  DFF_X1 \REGISTERS_reg[26][55]  ( .D(n5814), .CK(CLK), .Q(n50703), .QN(n54615) );
  DFF_X1 \REGISTERS_reg[26][54]  ( .D(n5813), .CK(CLK), .Q(n50702), .QN(n54616) );
  DFF_X1 \REGISTERS_reg[26][53]  ( .D(n5812), .CK(CLK), .Q(n50701), .QN(n54617) );
  DFF_X1 \REGISTERS_reg[26][52]  ( .D(n5811), .CK(CLK), .Q(n50700), .QN(n54618) );
  DFF_X1 \REGISTERS_reg[26][51]  ( .D(n5810), .CK(CLK), .Q(n50699), .QN(n54619) );
  DFF_X1 \REGISTERS_reg[26][50]  ( .D(n5809), .CK(CLK), .Q(n50698), .QN(n54620) );
  DFF_X1 \REGISTERS_reg[26][49]  ( .D(n5808), .CK(CLK), .Q(n50697), .QN(n54621) );
  DFF_X1 \REGISTERS_reg[26][48]  ( .D(n5807), .CK(CLK), .Q(n50696), .QN(n54622) );
  DFF_X1 \REGISTERS_reg[26][47]  ( .D(n5806), .CK(CLK), .Q(n50695), .QN(n54623) );
  DFF_X1 \REGISTERS_reg[26][46]  ( .D(n5805), .CK(CLK), .Q(n50694), .QN(n54624) );
  DFF_X1 \REGISTERS_reg[26][45]  ( .D(n5804), .CK(CLK), .Q(n50693), .QN(n54625) );
  DFF_X1 \REGISTERS_reg[26][44]  ( .D(n5803), .CK(CLK), .Q(n50692), .QN(n54626) );
  DFF_X1 \REGISTERS_reg[26][43]  ( .D(n5802), .CK(CLK), .Q(n50691), .QN(n54627) );
  DFF_X1 \REGISTERS_reg[26][42]  ( .D(n5801), .CK(CLK), .Q(n50690), .QN(n54628) );
  DFF_X1 \REGISTERS_reg[26][41]  ( .D(n5800), .CK(CLK), .Q(n50689), .QN(n54629) );
  DFF_X1 \REGISTERS_reg[26][40]  ( .D(n5799), .CK(CLK), .Q(n50688), .QN(n54630) );
  DFF_X1 \REGISTERS_reg[26][39]  ( .D(n5798), .CK(CLK), .Q(n50687), .QN(n54631) );
  DFF_X1 \REGISTERS_reg[26][38]  ( .D(n5797), .CK(CLK), .Q(n50686), .QN(n54632) );
  DFF_X1 \REGISTERS_reg[26][37]  ( .D(n5796), .CK(CLK), .Q(n50685), .QN(n54633) );
  DFF_X1 \REGISTERS_reg[26][36]  ( .D(n5795), .CK(CLK), .Q(n50684), .QN(n54634) );
  DFF_X1 \REGISTERS_reg[26][35]  ( .D(n5794), .CK(CLK), .Q(n50683), .QN(n54635) );
  DFF_X1 \REGISTERS_reg[26][34]  ( .D(n5793), .CK(CLK), .Q(n50682), .QN(n54636) );
  DFF_X1 \REGISTERS_reg[26][33]  ( .D(n5792), .CK(CLK), .Q(n50681), .QN(n54637) );
  DFF_X1 \REGISTERS_reg[26][32]  ( .D(n5791), .CK(CLK), .Q(n50680), .QN(n54638) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n5790), .CK(CLK), .Q(n50679), .QN(n54639) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n5789), .CK(CLK), .Q(n50678), .QN(n54640) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n5788), .CK(CLK), .Q(n50677), .QN(n54641) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n5787), .CK(CLK), .Q(n50676), .QN(n54642) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n5786), .CK(CLK), .Q(n50675), .QN(n54643) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n5785), .CK(CLK), .Q(n50674), .QN(n54644) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n5784), .CK(CLK), .Q(n50673), .QN(n54645) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n5783), .CK(CLK), .Q(n50672), .QN(n54646) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n5782), .CK(CLK), .Q(n50671), .QN(n54647) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n5781), .CK(CLK), .Q(n50670), .QN(n54648) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n5780), .CK(CLK), .Q(n50669), .QN(n54649) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n5779), .CK(CLK), .Q(n50668), .QN(n54650) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n5778), .CK(CLK), .Q(n50667), .QN(n54651) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n5777), .CK(CLK), .Q(n50666), .QN(n54652) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n5776), .CK(CLK), .Q(n50665), .QN(n54653) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n5775), .CK(CLK), .Q(n50664), .QN(n54654) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n5774), .CK(CLK), .Q(n50663), .QN(n54655) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n5773), .CK(CLK), .Q(n50662), .QN(n54656) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n5772), .CK(CLK), .Q(n50661), .QN(n54657) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n5771), .CK(CLK), .Q(n50660), .QN(n54658) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n5770), .CK(CLK), .Q(n50659), .QN(n54659) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n5769), .CK(CLK), .Q(n50658), .QN(n54660) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n5768), .CK(CLK), .Q(n50657), .QN(n54661)
         );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n5767), .CK(CLK), .Q(n50656), .QN(n54662)
         );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n5766), .CK(CLK), .Q(n50655), .QN(n54663)
         );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n5765), .CK(CLK), .Q(n50654), .QN(n54664)
         );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n5764), .CK(CLK), .Q(n50653), .QN(n54665)
         );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n5763), .CK(CLK), .Q(n50652), .QN(n54666)
         );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n5762), .CK(CLK), .Q(n50651), .QN(n54667)
         );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n5761), .CK(CLK), .Q(n50650), .QN(n54668)
         );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n5760), .CK(CLK), .Q(n50649), .QN(n54669)
         );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n5759), .CK(CLK), .Q(n50648), .QN(n54670)
         );
  DFF_X1 \REGISTERS_reg[10][59]  ( .D(n6842), .CK(CLK), .Q(n50576), .QN(n54187) );
  DFF_X1 \REGISTERS_reg[10][58]  ( .D(n6841), .CK(CLK), .Q(n50575), .QN(n54188) );
  DFF_X1 \REGISTERS_reg[10][57]  ( .D(n6840), .CK(CLK), .Q(n50574), .QN(n54189) );
  DFF_X1 \REGISTERS_reg[10][56]  ( .D(n6839), .CK(CLK), .Q(n50573), .QN(n54190) );
  DFF_X1 \REGISTERS_reg[10][55]  ( .D(n6838), .CK(CLK), .Q(n50572), .QN(n54191) );
  DFF_X1 \REGISTERS_reg[10][54]  ( .D(n6837), .CK(CLK), .Q(n50571), .QN(n54192) );
  DFF_X1 \REGISTERS_reg[10][53]  ( .D(n6836), .CK(CLK), .Q(n50570), .QN(n54193) );
  DFF_X1 \REGISTERS_reg[10][52]  ( .D(n6835), .CK(CLK), .Q(n50569), .QN(n54194) );
  DFF_X1 \REGISTERS_reg[10][51]  ( .D(n6834), .CK(CLK), .Q(n50568), .QN(n54195) );
  DFF_X1 \REGISTERS_reg[10][50]  ( .D(n6833), .CK(CLK), .Q(n50567), .QN(n54196) );
  DFF_X1 \REGISTERS_reg[10][49]  ( .D(n6832), .CK(CLK), .Q(n50566), .QN(n54197) );
  DFF_X1 \REGISTERS_reg[10][48]  ( .D(n6831), .CK(CLK), .Q(n50565), .QN(n54198) );
  DFF_X1 \REGISTERS_reg[10][47]  ( .D(n6830), .CK(CLK), .Q(n50564), .QN(n54199) );
  DFF_X1 \REGISTERS_reg[10][46]  ( .D(n6829), .CK(CLK), .Q(n50563), .QN(n54200) );
  DFF_X1 \REGISTERS_reg[10][45]  ( .D(n6828), .CK(CLK), .Q(n50562), .QN(n54201) );
  DFF_X1 \REGISTERS_reg[10][44]  ( .D(n6827), .CK(CLK), .Q(n50561), .QN(n54202) );
  DFF_X1 \REGISTERS_reg[10][43]  ( .D(n6826), .CK(CLK), .Q(n50560), .QN(n54203) );
  DFF_X1 \REGISTERS_reg[10][42]  ( .D(n6825), .CK(CLK), .Q(n50559), .QN(n54204) );
  DFF_X1 \REGISTERS_reg[10][41]  ( .D(n6824), .CK(CLK), .Q(n50558), .QN(n54205) );
  DFF_X1 \REGISTERS_reg[10][40]  ( .D(n6823), .CK(CLK), .Q(n50557), .QN(n54206) );
  DFF_X1 \REGISTERS_reg[10][39]  ( .D(n6822), .CK(CLK), .Q(n50556), .QN(n54207) );
  DFF_X1 \REGISTERS_reg[10][38]  ( .D(n6821), .CK(CLK), .Q(n50555), .QN(n54208) );
  DFF_X1 \REGISTERS_reg[10][37]  ( .D(n6820), .CK(CLK), .Q(n50554), .QN(n54209) );
  DFF_X1 \REGISTERS_reg[10][36]  ( .D(n6819), .CK(CLK), .Q(n50553), .QN(n54210) );
  DFF_X1 \REGISTERS_reg[10][35]  ( .D(n6818), .CK(CLK), .Q(n50552), .QN(n54211) );
  DFF_X1 \REGISTERS_reg[10][34]  ( .D(n6817), .CK(CLK), .Q(n50551), .QN(n54212) );
  DFF_X1 \REGISTERS_reg[10][33]  ( .D(n6816), .CK(CLK), .Q(n50550), .QN(n54213) );
  DFF_X1 \REGISTERS_reg[10][32]  ( .D(n6815), .CK(CLK), .Q(n50549), .QN(n54214) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n6814), .CK(CLK), .Q(n50548), .QN(n54215) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n6813), .CK(CLK), .Q(n50547), .QN(n54216) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n6812), .CK(CLK), .Q(n50546), .QN(n54217) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n6811), .CK(CLK), .Q(n50545), .QN(n54218) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n6810), .CK(CLK), .Q(n50544), .QN(n54219) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n6809), .CK(CLK), .Q(n50543), .QN(n54220) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n6808), .CK(CLK), .Q(n50542), .QN(n54221) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n6807), .CK(CLK), .Q(n50541), .QN(n54222) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n6806), .CK(CLK), .Q(n50540), .QN(n54223) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n6805), .CK(CLK), .Q(n50539), .QN(n54224) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n6804), .CK(CLK), .Q(n50538), .QN(n54225) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n6803), .CK(CLK), .Q(n50537), .QN(n54226) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n6802), .CK(CLK), .Q(n50536), .QN(n54227) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n6801), .CK(CLK), .Q(n50535), .QN(n54228) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n6800), .CK(CLK), .Q(n50534), .QN(n54229) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n6799), .CK(CLK), .Q(n50533), .QN(n54230) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n6798), .CK(CLK), .Q(n50532), .QN(n54231) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n6797), .CK(CLK), .Q(n50531), .QN(n54232) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n6796), .CK(CLK), .Q(n50530), .QN(n54233) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n6795), .CK(CLK), .Q(n50529), .QN(n54234) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n6794), .CK(CLK), .Q(n50528), .QN(n54235) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n6793), .CK(CLK), .Q(n50527), .QN(n54236) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n6792), .CK(CLK), .Q(n50526), .QN(n54237)
         );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n6791), .CK(CLK), .Q(n50525), .QN(n54238)
         );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n6790), .CK(CLK), .Q(n50524), .QN(n54239)
         );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n6789), .CK(CLK), .Q(n50523), .QN(n54240)
         );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n6788), .CK(CLK), .Q(n50522), .QN(n54241)
         );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n6787), .CK(CLK), .Q(n50521), .QN(n54242)
         );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n6786), .CK(CLK), .Q(n50520), .QN(n54243)
         );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n6785), .CK(CLK), .Q(n50519), .QN(n54244)
         );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n6784), .CK(CLK), .Q(n50518), .QN(n54245)
         );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n6783), .CK(CLK), .Q(n50517), .QN(n54246)
         );
  DFF_X1 \OUT2_reg[63]  ( .D(n5374), .CK(CLK), .Q(OUT2[63]) );
  DFF_X1 \OUT2_reg[62]  ( .D(n5373), .CK(CLK), .Q(OUT2[62]) );
  NOR3_X2 U45435 ( .A1(n67434), .A2(ADD_RD2[2]), .A3(n66301), .ZN(n66283) );
  NAND3_X1 U45452 ( .A1(n62490), .A2(n62491), .A3(n62492), .ZN(n62088) );
  NAND3_X1 U45453 ( .A1(n62492), .A2(n62491), .A3(ADD_WR[0]), .ZN(n62156) );
  NAND3_X1 U45454 ( .A1(n62492), .A2(n62490), .A3(ADD_WR[3]), .ZN(n62625) );
  NAND3_X1 U45455 ( .A1(ADD_WR[0]), .A2(n62492), .A3(ADD_WR[3]), .ZN(n62692)
         );
  NAND3_X1 U45456 ( .A1(n62490), .A2(n62491), .A3(n63295), .ZN(n63025) );
  NAND3_X1 U45457 ( .A1(ADD_WR[0]), .A2(n62491), .A3(n63295), .ZN(n63092) );
  NAND3_X1 U45458 ( .A1(ADD_WR[3]), .A2(n62490), .A3(n63295), .ZN(n63428) );
  NAND3_X1 U45459 ( .A1(ADD_WR[3]), .A2(ADD_WR[0]), .A3(n63295), .ZN(n63495)
         );
  NAND3_X1 U45461 ( .A1(ENABLE), .A2(n68057), .A3(RD2), .ZN(n65112) );
  DFF_X1 \REGISTERS_reg[31][63]  ( .D(n5502), .CK(CLK), .Q(n58378), .QN(n63765) );
  DFF_X1 \REGISTERS_reg[31][62]  ( .D(n5500), .CK(CLK), .Q(n58377), .QN(n63820) );
  DFF_X1 \REGISTERS_reg[31][61]  ( .D(n5498), .CK(CLK), .Q(n58376), .QN(n63841) );
  DFF_X1 \REGISTERS_reg[31][60]  ( .D(n5496), .CK(CLK), .Q(n58375), .QN(n63862) );
  DFF_X1 \REGISTERS_reg[30][63]  ( .D(n5566), .CK(CLK), .Q(n66308), .QN(n63699) );
  DFF_X1 \REGISTERS_reg[30][62]  ( .D(n5565), .CK(CLK), .Q(n66307), .QN(n63701) );
  DFF_X1 \REGISTERS_reg[30][61]  ( .D(n5564), .CK(CLK), .Q(n66306), .QN(n63702) );
  DFF_X1 \REGISTERS_reg[30][60]  ( .D(n5563), .CK(CLK), .Q(n66305), .QN(n63703) );
  DFF_X1 \REGISTERS_reg[29][63]  ( .D(n5630), .CK(CLK), .QN(n63633) );
  DFF_X1 \REGISTERS_reg[29][62]  ( .D(n5629), .CK(CLK), .QN(n63635) );
  DFF_X1 \REGISTERS_reg[29][61]  ( .D(n5628), .CK(CLK), .QN(n63636) );
  DFF_X1 \REGISTERS_reg[29][60]  ( .D(n5627), .CK(CLK), .QN(n63637) );
  DFF_X1 \REGISTERS_reg[28][63]  ( .D(n5694), .CK(CLK), .QN(n63567) );
  DFF_X1 \REGISTERS_reg[28][62]  ( .D(n5693), .CK(CLK), .QN(n63569) );
  DFF_X1 \REGISTERS_reg[28][61]  ( .D(n5692), .CK(CLK), .QN(n63570) );
  DFF_X1 \REGISTERS_reg[28][60]  ( .D(n5691), .CK(CLK), .QN(n63571) );
  DFF_X1 \REGISTERS_reg[27][63]  ( .D(n5758), .CK(CLK), .QN(n63501) );
  DFF_X1 \REGISTERS_reg[27][62]  ( .D(n5757), .CK(CLK), .QN(n63503) );
  DFF_X1 \REGISTERS_reg[27][61]  ( .D(n5756), .CK(CLK), .QN(n63504) );
  DFF_X1 \REGISTERS_reg[27][60]  ( .D(n5755), .CK(CLK), .QN(n63505) );
  DFF_X1 \REGISTERS_reg[25][63]  ( .D(n5886), .CK(CLK), .Q(n8959), .QN(n63430)
         );
  DFF_X1 \REGISTERS_reg[25][62]  ( .D(n5885), .CK(CLK), .Q(n8961), .QN(n63432)
         );
  DFF_X1 \REGISTERS_reg[25][61]  ( .D(n5884), .CK(CLK), .Q(n8963), .QN(n63433)
         );
  DFF_X1 \REGISTERS_reg[25][60]  ( .D(n5883), .CK(CLK), .Q(n8965), .QN(n63434)
         );
  DFF_X1 \REGISTERS_reg[23][63]  ( .D(n6014), .CK(CLK), .QN(n63297) );
  DFF_X1 \REGISTERS_reg[23][62]  ( .D(n6013), .CK(CLK), .QN(n63299) );
  DFF_X1 \REGISTERS_reg[23][61]  ( .D(n6012), .CK(CLK), .QN(n63300) );
  DFF_X1 \REGISTERS_reg[23][60]  ( .D(n6011), .CK(CLK), .QN(n63301) );
  DFF_X1 \REGISTERS_reg[19][63]  ( .D(n6270), .CK(CLK), .QN(n63096) );
  DFF_X1 \REGISTERS_reg[19][62]  ( .D(n6269), .CK(CLK), .QN(n63098) );
  DFF_X1 \REGISTERS_reg[19][61]  ( .D(n6268), .CK(CLK), .QN(n63099) );
  DFF_X1 \REGISTERS_reg[19][60]  ( .D(n6267), .CK(CLK), .QN(n63100) );
  DFF_X1 \REGISTERS_reg[24][63]  ( .D(n5950), .CK(CLK), .QN(n63363) );
  DFF_X1 \REGISTERS_reg[24][62]  ( .D(n5949), .CK(CLK), .QN(n63365) );
  DFF_X1 \REGISTERS_reg[24][61]  ( .D(n5948), .CK(CLK), .QN(n63366) );
  DFF_X1 \REGISTERS_reg[24][60]  ( .D(n5947), .CK(CLK), .QN(n63367) );
  DFF_X1 \REGISTERS_reg[17][63]  ( .D(n6398), .CK(CLK), .Q(n58234), .QN(n63027) );
  DFF_X1 \REGISTERS_reg[17][62]  ( .D(n6397), .CK(CLK), .Q(n58233), .QN(n63029) );
  DFF_X1 \REGISTERS_reg[17][61]  ( .D(n6396), .CK(CLK), .Q(n58232), .QN(n63030) );
  DFF_X1 \REGISTERS_reg[17][60]  ( .D(n6395), .CK(CLK), .Q(n58231), .QN(n63031) );
  DFF_X1 \REGISTERS_reg[16][63]  ( .D(n6462), .CK(CLK), .Q(n58370), .QN(n62960) );
  DFF_X1 \REGISTERS_reg[16][62]  ( .D(n6461), .CK(CLK), .Q(n58369), .QN(n62962) );
  DFF_X1 \REGISTERS_reg[16][61]  ( .D(n6460), .CK(CLK), .Q(n58368), .QN(n62963) );
  DFF_X1 \REGISTERS_reg[16][60]  ( .D(n6459), .CK(CLK), .Q(n58367), .QN(n62964) );
  DFF_X1 \REGISTERS_reg[22][63]  ( .D(n6078), .CK(CLK), .Q(n58718), .QN(n63230) );
  DFF_X1 \REGISTERS_reg[22][62]  ( .D(n6077), .CK(CLK), .Q(n58717), .QN(n63232) );
  DFF_X1 \REGISTERS_reg[22][61]  ( .D(n6076), .CK(CLK), .Q(n58716), .QN(n63233) );
  DFF_X1 \REGISTERS_reg[22][60]  ( .D(n6075), .CK(CLK), .Q(n58715), .QN(n63234) );
  DFF_X1 \REGISTERS_reg[20][63]  ( .D(n6206), .CK(CLK), .Q(n58301), .QN(n63162) );
  DFF_X1 \REGISTERS_reg[20][62]  ( .D(n6205), .CK(CLK), .Q(n58299), .QN(n63164) );
  DFF_X1 \REGISTERS_reg[20][61]  ( .D(n6204), .CK(CLK), .Q(n58297), .QN(n63165) );
  DFF_X1 \REGISTERS_reg[20][60]  ( .D(n6203), .CK(CLK), .Q(n58295), .QN(n63166) );
  DFF_X1 \REGISTERS_reg[10][63]  ( .D(n6846), .CK(CLK), .QN(n62694) );
  DFF_X1 \REGISTERS_reg[0][63]  ( .D(n7486), .CK(CLK), .Q(n56490), .QN(n61958)
         );
  DFF_X1 \REGISTERS_reg[0][62]  ( .D(n7485), .CK(CLK), .Q(n56531), .QN(n61961)
         );
  DFF_X1 \REGISTERS_reg[0][61]  ( .D(n7484), .CK(CLK), .Q(n56555), .QN(n61963)
         );
  DFF_X1 \REGISTERS_reg[0][60]  ( .D(n7483), .CK(CLK), .Q(n56579), .QN(n61965)
         );
  DFF_X1 \REGISTERS_reg[7][63]  ( .D(n7038), .CK(CLK), .Q(n58050), .QN(n62494)
         );
  DFF_X1 \REGISTERS_reg[7][62]  ( .D(n7037), .CK(CLK), .Q(n58049), .QN(n62496)
         );
  DFF_X1 \REGISTERS_reg[7][61]  ( .D(n7036), .CK(CLK), .Q(n58048), .QN(n62497)
         );
  DFF_X1 \REGISTERS_reg[7][60]  ( .D(n7035), .CK(CLK), .Q(n58047), .QN(n62498)
         );
  DFF_X1 \REGISTERS_reg[5][63]  ( .D(n7166), .CK(CLK), .Q(n58782), .QN(n62358)
         );
  DFF_X1 \REGISTERS_reg[5][62]  ( .D(n7165), .CK(CLK), .Q(n58781), .QN(n62360)
         );
  DFF_X1 \REGISTERS_reg[5][61]  ( .D(n7164), .CK(CLK), .Q(n58780), .QN(n62361)
         );
  DFF_X1 \REGISTERS_reg[5][60]  ( .D(n7163), .CK(CLK), .Q(n58779), .QN(n62362)
         );
  DFF_X1 \REGISTERS_reg[3][63]  ( .D(n7294), .CK(CLK), .QN(n62225) );
  DFF_X1 \REGISTERS_reg[3][62]  ( .D(n7293), .CK(CLK), .QN(n62227) );
  DFF_X1 \REGISTERS_reg[3][61]  ( .D(n7292), .CK(CLK), .QN(n62228) );
  DFF_X1 \REGISTERS_reg[3][60]  ( .D(n7291), .CK(CLK), .QN(n62229) );
  DFF_X1 \REGISTERS_reg[2][63]  ( .D(n7358), .CK(CLK), .QN(n62158) );
  DFF_X1 \REGISTERS_reg[2][62]  ( .D(n7357), .CK(CLK), .QN(n62160) );
  DFF_X1 \REGISTERS_reg[2][61]  ( .D(n7356), .CK(CLK), .QN(n62161) );
  DFF_X1 \REGISTERS_reg[2][60]  ( .D(n7355), .CK(CLK), .QN(n62162) );
  DFF_X1 \REGISTERS_reg[31][59]  ( .D(n5494), .CK(CLK), .Q(n58438), .QN(n63883) );
  DFF_X1 \REGISTERS_reg[31][58]  ( .D(n5492), .CK(CLK), .Q(n58437), .QN(n63903) );
  DFF_X1 \REGISTERS_reg[31][57]  ( .D(n5490), .CK(CLK), .Q(n58436), .QN(n63923) );
  DFF_X1 \REGISTERS_reg[31][56]  ( .D(n5488), .CK(CLK), .Q(n58435), .QN(n63943) );
  DFF_X1 \REGISTERS_reg[31][55]  ( .D(n5486), .CK(CLK), .Q(n58434), .QN(n63963) );
  DFF_X1 \REGISTERS_reg[31][54]  ( .D(n5484), .CK(CLK), .Q(n58433), .QN(n63983) );
  DFF_X1 \REGISTERS_reg[31][53]  ( .D(n5482), .CK(CLK), .Q(n58432), .QN(n64003) );
  DFF_X1 \REGISTERS_reg[31][52]  ( .D(n5480), .CK(CLK), .Q(n58431), .QN(n64023) );
  DFF_X1 \REGISTERS_reg[31][51]  ( .D(n5478), .CK(CLK), .Q(n58430), .QN(n64043) );
  DFF_X1 \REGISTERS_reg[31][50]  ( .D(n5476), .CK(CLK), .Q(n58429), .QN(n64063) );
  DFF_X1 \REGISTERS_reg[31][49]  ( .D(n5474), .CK(CLK), .Q(n58428), .QN(n64083) );
  DFF_X1 \REGISTERS_reg[31][48]  ( .D(n5472), .CK(CLK), .Q(n58427), .QN(n64103) );
  DFF_X1 \REGISTERS_reg[31][47]  ( .D(n5470), .CK(CLK), .Q(n58426), .QN(n64123) );
  DFF_X1 \REGISTERS_reg[31][46]  ( .D(n5468), .CK(CLK), .Q(n58425), .QN(n64143) );
  DFF_X1 \REGISTERS_reg[31][45]  ( .D(n5466), .CK(CLK), .Q(n58424), .QN(n64163) );
  DFF_X1 \REGISTERS_reg[31][44]  ( .D(n5464), .CK(CLK), .Q(n58423), .QN(n64183) );
  DFF_X1 \REGISTERS_reg[31][43]  ( .D(n5462), .CK(CLK), .Q(n58422), .QN(n64203) );
  DFF_X1 \REGISTERS_reg[31][42]  ( .D(n5460), .CK(CLK), .Q(n58421), .QN(n64223) );
  DFF_X1 \REGISTERS_reg[31][41]  ( .D(n5458), .CK(CLK), .Q(n58420), .QN(n64243) );
  DFF_X1 \REGISTERS_reg[31][40]  ( .D(n5456), .CK(CLK), .Q(n58419), .QN(n64263) );
  DFF_X1 \REGISTERS_reg[31][39]  ( .D(n5454), .CK(CLK), .Q(n58418), .QN(n64283) );
  DFF_X1 \REGISTERS_reg[31][38]  ( .D(n5452), .CK(CLK), .Q(n58417), .QN(n64303) );
  DFF_X1 \REGISTERS_reg[31][37]  ( .D(n5450), .CK(CLK), .Q(n58416), .QN(n64323) );
  DFF_X1 \REGISTERS_reg[31][36]  ( .D(n5448), .CK(CLK), .Q(n58415), .QN(n64343) );
  DFF_X1 \REGISTERS_reg[31][35]  ( .D(n5446), .CK(CLK), .Q(n58414), .QN(n64363) );
  DFF_X1 \REGISTERS_reg[31][34]  ( .D(n5444), .CK(CLK), .Q(n58413), .QN(n64383) );
  DFF_X1 \REGISTERS_reg[31][33]  ( .D(n5442), .CK(CLK), .Q(n58412), .QN(n64403) );
  DFF_X1 \REGISTERS_reg[31][32]  ( .D(n5440), .CK(CLK), .Q(n58411), .QN(n64423) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n5438), .CK(CLK), .Q(n58410), .QN(n64443) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n5436), .CK(CLK), .Q(n58409), .QN(n64463) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n5434), .CK(CLK), .Q(n58408), .QN(n64483) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n5432), .CK(CLK), .Q(n58407), .QN(n64503) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n5430), .CK(CLK), .Q(n58406), .QN(n64523) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n5428), .CK(CLK), .Q(n58405), .QN(n64543) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n5426), .CK(CLK), .Q(n58404), .QN(n64563) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n5424), .CK(CLK), .Q(n58403), .QN(n64583) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n5422), .CK(CLK), .Q(n58402), .QN(n64603) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n5420), .CK(CLK), .Q(n58401), .QN(n64623) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n5418), .CK(CLK), .Q(n58400), .QN(n64643) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n5416), .CK(CLK), .Q(n58399), .QN(n64663) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n5414), .CK(CLK), .Q(n58398), .QN(n64683) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n5412), .CK(CLK), .Q(n58397), .QN(n64703) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n5410), .CK(CLK), .Q(n58396), .QN(n64723) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n5408), .CK(CLK), .Q(n58395), .QN(n64743) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n5406), .CK(CLK), .Q(n58394), .QN(n64763) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n5404), .CK(CLK), .Q(n58393), .QN(n64783) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n5402), .CK(CLK), .Q(n58392), .QN(n64803) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n5400), .CK(CLK), .Q(n58391), .QN(n64823) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n5398), .CK(CLK), .Q(n58390), .QN(n64843) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n5396), .CK(CLK), .Q(n58389), .QN(n64863) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n5394), .CK(CLK), .Q(n58388), .QN(n64883)
         );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n5392), .CK(CLK), .Q(n58387), .QN(n64903)
         );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n5390), .CK(CLK), .Q(n58386), .QN(n64923)
         );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n5388), .CK(CLK), .Q(n58385), .QN(n64943)
         );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n5386), .CK(CLK), .Q(n58384), .QN(n64963)
         );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n5384), .CK(CLK), .Q(n58383), .QN(n64983)
         );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n5382), .CK(CLK), .Q(n58382), .QN(n65003)
         );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n5380), .CK(CLK), .Q(n58381), .QN(n65023)
         );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n5378), .CK(CLK), .Q(n58380), .QN(n65043)
         );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n5376), .CK(CLK), .Q(n58379), .QN(n65063)
         );
  DFF_X1 \REGISTERS_reg[6][63]  ( .D(n7102), .CK(CLK), .QN(n62424) );
  DFF_X1 \REGISTERS_reg[6][62]  ( .D(n7101), .CK(CLK), .QN(n62426) );
  DFF_X1 \REGISTERS_reg[6][61]  ( .D(n7100), .CK(CLK), .QN(n62427) );
  DFF_X1 \REGISTERS_reg[6][60]  ( .D(n7099), .CK(CLK), .QN(n62428) );
  DFF_X1 \REGISTERS_reg[4][63]  ( .D(n7230), .CK(CLK), .Q(n59092), .QN(n62291)
         );
  DFF_X1 \REGISTERS_reg[4][62]  ( .D(n7229), .CK(CLK), .Q(n59091), .QN(n62293)
         );
  DFF_X1 \REGISTERS_reg[4][61]  ( .D(n7228), .CK(CLK), .Q(n59090), .QN(n62294)
         );
  DFF_X1 \REGISTERS_reg[4][60]  ( .D(n7227), .CK(CLK), .Q(n59089), .QN(n62295)
         );
  DFF_X1 \REGISTERS_reg[1][63]  ( .D(n7422), .CK(CLK), .QN(n62091) );
  DFF_X1 \REGISTERS_reg[1][62]  ( .D(n7421), .CK(CLK), .QN(n62093) );
  DFF_X1 \REGISTERS_reg[1][61]  ( .D(n7420), .CK(CLK), .QN(n62094) );
  DFF_X1 \REGISTERS_reg[1][60]  ( .D(n7419), .CK(CLK), .QN(n62095) );
  DFF_X1 \REGISTERS_reg[8][63]  ( .D(n6974), .CK(CLK), .Q(n58303), .QN(n62560)
         );
  DFF_X1 \REGISTERS_reg[8][62]  ( .D(n6973), .CK(CLK), .Q(n58306), .QN(n62562)
         );
  DFF_X1 \REGISTERS_reg[8][61]  ( .D(n6972), .CK(CLK), .Q(n58305), .QN(n62563)
         );
  DFF_X1 \REGISTERS_reg[8][60]  ( .D(n6971), .CK(CLK), .Q(n58304), .QN(n62564)
         );
  DFF_X1 \REGISTERS_reg[14][63]  ( .D(n6590), .CK(CLK), .Q(n58783), .QN(n62827) );
  DFF_X1 \REGISTERS_reg[14][62]  ( .D(n6589), .CK(CLK), .Q(n58786), .QN(n62829) );
  DFF_X1 \REGISTERS_reg[14][61]  ( .D(n6588), .CK(CLK), .Q(n58785), .QN(n62830) );
  DFF_X1 \REGISTERS_reg[14][60]  ( .D(n6587), .CK(CLK), .Q(n58784), .QN(n62831) );
  DFF_X1 \REGISTERS_reg[30][59]  ( .D(n5562), .CK(CLK), .Q(n66372), .QN(n63704) );
  DFF_X1 \REGISTERS_reg[30][58]  ( .D(n5561), .CK(CLK), .Q(n66371), .QN(n63705) );
  DFF_X1 \REGISTERS_reg[30][57]  ( .D(n5560), .CK(CLK), .Q(n66370), .QN(n63706) );
  DFF_X1 \REGISTERS_reg[30][56]  ( .D(n5559), .CK(CLK), .Q(n66369), .QN(n63707) );
  DFF_X1 \REGISTERS_reg[30][55]  ( .D(n5558), .CK(CLK), .Q(n66368), .QN(n63708) );
  DFF_X1 \REGISTERS_reg[30][54]  ( .D(n5557), .CK(CLK), .Q(n66367), .QN(n63709) );
  DFF_X1 \REGISTERS_reg[30][53]  ( .D(n5556), .CK(CLK), .Q(n66366), .QN(n63710) );
  DFF_X1 \REGISTERS_reg[30][52]  ( .D(n5555), .CK(CLK), .Q(n66365), .QN(n63711) );
  DFF_X1 \REGISTERS_reg[30][51]  ( .D(n5554), .CK(CLK), .Q(n66364), .QN(n63712) );
  DFF_X1 \REGISTERS_reg[30][50]  ( .D(n5553), .CK(CLK), .Q(n66363), .QN(n63713) );
  DFF_X1 \REGISTERS_reg[30][49]  ( .D(n5552), .CK(CLK), .Q(n66362), .QN(n63714) );
  DFF_X1 \REGISTERS_reg[30][48]  ( .D(n5551), .CK(CLK), .Q(n66361), .QN(n63715) );
  DFF_X1 \REGISTERS_reg[30][47]  ( .D(n5550), .CK(CLK), .Q(n66360), .QN(n63716) );
  DFF_X1 \REGISTERS_reg[30][46]  ( .D(n5549), .CK(CLK), .Q(n66359), .QN(n63717) );
  DFF_X1 \REGISTERS_reg[30][45]  ( .D(n5548), .CK(CLK), .Q(n66358), .QN(n63718) );
  DFF_X1 \REGISTERS_reg[30][44]  ( .D(n5547), .CK(CLK), .Q(n66357), .QN(n63719) );
  DFF_X1 \REGISTERS_reg[30][43]  ( .D(n5546), .CK(CLK), .Q(n66356), .QN(n63720) );
  DFF_X1 \REGISTERS_reg[30][42]  ( .D(n5545), .CK(CLK), .Q(n66355), .QN(n63721) );
  DFF_X1 \REGISTERS_reg[30][41]  ( .D(n5544), .CK(CLK), .Q(n66354), .QN(n63722) );
  DFF_X1 \REGISTERS_reg[30][40]  ( .D(n5543), .CK(CLK), .Q(n66353), .QN(n63723) );
  DFF_X1 \REGISTERS_reg[30][39]  ( .D(n5542), .CK(CLK), .Q(n66352), .QN(n63724) );
  DFF_X1 \REGISTERS_reg[30][38]  ( .D(n5541), .CK(CLK), .Q(n66351), .QN(n63725) );
  DFF_X1 \REGISTERS_reg[30][37]  ( .D(n5540), .CK(CLK), .Q(n66350), .QN(n63726) );
  DFF_X1 \REGISTERS_reg[30][36]  ( .D(n5539), .CK(CLK), .Q(n66349), .QN(n63727) );
  DFF_X1 \REGISTERS_reg[30][35]  ( .D(n5538), .CK(CLK), .Q(n66348), .QN(n63728) );
  DFF_X1 \REGISTERS_reg[30][34]  ( .D(n5537), .CK(CLK), .Q(n66347), .QN(n63729) );
  DFF_X1 \REGISTERS_reg[30][33]  ( .D(n5536), .CK(CLK), .Q(n66346), .QN(n63730) );
  DFF_X1 \REGISTERS_reg[30][32]  ( .D(n5535), .CK(CLK), .Q(n66345), .QN(n63731) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n5534), .CK(CLK), .Q(n66344), .QN(n63732) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n5533), .CK(CLK), .Q(n66343), .QN(n63733) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n5532), .CK(CLK), .Q(n66342), .QN(n63734) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n5531), .CK(CLK), .Q(n66341), .QN(n63735) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n5530), .CK(CLK), .Q(n66340), .QN(n63736) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n5529), .CK(CLK), .Q(n66339), .QN(n63737) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n5528), .CK(CLK), .Q(n66338), .QN(n63738) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n5527), .CK(CLK), .Q(n66337), .QN(n63739) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n5526), .CK(CLK), .Q(n66336), .QN(n63740) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n5525), .CK(CLK), .Q(n66335), .QN(n63741) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n5524), .CK(CLK), .Q(n66334), .QN(n63742) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n5523), .CK(CLK), .Q(n66333), .QN(n63743) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n5522), .CK(CLK), .Q(n66332), .QN(n63744) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n5521), .CK(CLK), .Q(n66331), .QN(n63745) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n5520), .CK(CLK), .Q(n66330), .QN(n63746) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n5519), .CK(CLK), .Q(n66329), .QN(n63747) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n5518), .CK(CLK), .Q(n66328), .QN(n63748) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n5517), .CK(CLK), .Q(n66327), .QN(n63749) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n5516), .CK(CLK), .Q(n66326), .QN(n63750) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n5515), .CK(CLK), .Q(n66325), .QN(n63751) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n5514), .CK(CLK), .Q(n66324), .QN(n63752) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n5513), .CK(CLK), .Q(n66323), .QN(n63753) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n5512), .CK(CLK), .Q(n66322), .QN(n63754)
         );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n5511), .CK(CLK), .Q(n66321), .QN(n63755)
         );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n5510), .CK(CLK), .Q(n66320), .QN(n63756)
         );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n5509), .CK(CLK), .Q(n66319), .QN(n63757)
         );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n5508), .CK(CLK), .Q(n66318), .QN(n63758)
         );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n5507), .CK(CLK), .Q(n66317), .QN(n63759)
         );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n5506), .CK(CLK), .Q(n66316), .QN(n63760)
         );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n5505), .CK(CLK), .Q(n66315), .QN(n63761)
         );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n5504), .CK(CLK), .Q(n66314), .QN(n63762)
         );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n5503), .CK(CLK), .Q(n66313), .QN(n63763)
         );
  DFF_X1 \REGISTERS_reg[29][59]  ( .D(n5626), .CK(CLK), .QN(n63638) );
  DFF_X1 \REGISTERS_reg[29][58]  ( .D(n5625), .CK(CLK), .QN(n63639) );
  DFF_X1 \REGISTERS_reg[29][57]  ( .D(n5624), .CK(CLK), .QN(n63640) );
  DFF_X1 \REGISTERS_reg[29][56]  ( .D(n5623), .CK(CLK), .QN(n63641) );
  DFF_X1 \REGISTERS_reg[29][55]  ( .D(n5622), .CK(CLK), .QN(n63642) );
  DFF_X1 \REGISTERS_reg[29][54]  ( .D(n5621), .CK(CLK), .QN(n63643) );
  DFF_X1 \REGISTERS_reg[29][53]  ( .D(n5620), .CK(CLK), .QN(n63644) );
  DFF_X1 \REGISTERS_reg[29][52]  ( .D(n5619), .CK(CLK), .QN(n63645) );
  DFF_X1 \REGISTERS_reg[29][51]  ( .D(n5618), .CK(CLK), .QN(n63646) );
  DFF_X1 \REGISTERS_reg[29][50]  ( .D(n5617), .CK(CLK), .QN(n63647) );
  DFF_X1 \REGISTERS_reg[29][49]  ( .D(n5616), .CK(CLK), .QN(n63648) );
  DFF_X1 \REGISTERS_reg[29][48]  ( .D(n5615), .CK(CLK), .QN(n63649) );
  DFF_X1 \REGISTERS_reg[29][47]  ( .D(n5614), .CK(CLK), .QN(n63650) );
  DFF_X1 \REGISTERS_reg[29][46]  ( .D(n5613), .CK(CLK), .QN(n63651) );
  DFF_X1 \REGISTERS_reg[29][45]  ( .D(n5612), .CK(CLK), .QN(n63652) );
  DFF_X1 \REGISTERS_reg[29][44]  ( .D(n5611), .CK(CLK), .QN(n63653) );
  DFF_X1 \REGISTERS_reg[29][43]  ( .D(n5610), .CK(CLK), .QN(n63654) );
  DFF_X1 \REGISTERS_reg[29][42]  ( .D(n5609), .CK(CLK), .QN(n63655) );
  DFF_X1 \REGISTERS_reg[29][41]  ( .D(n5608), .CK(CLK), .QN(n63656) );
  DFF_X1 \REGISTERS_reg[29][40]  ( .D(n5607), .CK(CLK), .QN(n63657) );
  DFF_X1 \REGISTERS_reg[29][39]  ( .D(n5606), .CK(CLK), .QN(n63658) );
  DFF_X1 \REGISTERS_reg[29][38]  ( .D(n5605), .CK(CLK), .QN(n63659) );
  DFF_X1 \REGISTERS_reg[29][37]  ( .D(n5604), .CK(CLK), .QN(n63660) );
  DFF_X1 \REGISTERS_reg[29][36]  ( .D(n5603), .CK(CLK), .QN(n63661) );
  DFF_X1 \REGISTERS_reg[29][35]  ( .D(n5602), .CK(CLK), .QN(n63662) );
  DFF_X1 \REGISTERS_reg[29][34]  ( .D(n5601), .CK(CLK), .QN(n63663) );
  DFF_X1 \REGISTERS_reg[29][33]  ( .D(n5600), .CK(CLK), .QN(n63664) );
  DFF_X1 \REGISTERS_reg[29][32]  ( .D(n5599), .CK(CLK), .QN(n63665) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n5598), .CK(CLK), .QN(n63666) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n5597), .CK(CLK), .QN(n63667) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n5596), .CK(CLK), .QN(n63668) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n5595), .CK(CLK), .QN(n63669) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n5594), .CK(CLK), .QN(n63670) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n5593), .CK(CLK), .QN(n63671) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n5592), .CK(CLK), .QN(n63672) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n5591), .CK(CLK), .QN(n63673) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n5590), .CK(CLK), .QN(n63674) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n5589), .CK(CLK), .QN(n63675) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n5588), .CK(CLK), .QN(n63676) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n5587), .CK(CLK), .QN(n63677) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n5586), .CK(CLK), .QN(n63678) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n5585), .CK(CLK), .QN(n63679) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n5584), .CK(CLK), .QN(n63680) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n5583), .CK(CLK), .QN(n63681) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n5582), .CK(CLK), .QN(n63682) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n5581), .CK(CLK), .QN(n63683) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n5580), .CK(CLK), .QN(n63684) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n5579), .CK(CLK), .QN(n63685) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n5578), .CK(CLK), .QN(n63686) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n5577), .CK(CLK), .QN(n63687) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n5576), .CK(CLK), .QN(n63688) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n5575), .CK(CLK), .QN(n63689) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n5574), .CK(CLK), .QN(n63690) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n5573), .CK(CLK), .QN(n63691) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n5572), .CK(CLK), .QN(n63692) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n5571), .CK(CLK), .QN(n63693) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n5570), .CK(CLK), .QN(n63694) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n5569), .CK(CLK), .QN(n63695) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n5568), .CK(CLK), .QN(n63696) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n5567), .CK(CLK), .QN(n63697) );
  DFF_X1 \REGISTERS_reg[28][59]  ( .D(n5690), .CK(CLK), .QN(n63572) );
  DFF_X1 \REGISTERS_reg[28][58]  ( .D(n5689), .CK(CLK), .QN(n63573) );
  DFF_X1 \REGISTERS_reg[28][57]  ( .D(n5688), .CK(CLK), .QN(n63574) );
  DFF_X1 \REGISTERS_reg[28][56]  ( .D(n5687), .CK(CLK), .QN(n63575) );
  DFF_X1 \REGISTERS_reg[28][55]  ( .D(n5686), .CK(CLK), .QN(n63576) );
  DFF_X1 \REGISTERS_reg[28][54]  ( .D(n5685), .CK(CLK), .QN(n63577) );
  DFF_X1 \REGISTERS_reg[28][53]  ( .D(n5684), .CK(CLK), .QN(n63578) );
  DFF_X1 \REGISTERS_reg[28][52]  ( .D(n5683), .CK(CLK), .QN(n63579) );
  DFF_X1 \REGISTERS_reg[28][51]  ( .D(n5682), .CK(CLK), .QN(n63580) );
  DFF_X1 \REGISTERS_reg[28][50]  ( .D(n5681), .CK(CLK), .QN(n63581) );
  DFF_X1 \REGISTERS_reg[28][49]  ( .D(n5680), .CK(CLK), .QN(n63582) );
  DFF_X1 \REGISTERS_reg[28][48]  ( .D(n5679), .CK(CLK), .QN(n63583) );
  DFF_X1 \REGISTERS_reg[28][47]  ( .D(n5678), .CK(CLK), .QN(n63584) );
  DFF_X1 \REGISTERS_reg[28][46]  ( .D(n5677), .CK(CLK), .QN(n63585) );
  DFF_X1 \REGISTERS_reg[28][45]  ( .D(n5676), .CK(CLK), .QN(n63586) );
  DFF_X1 \REGISTERS_reg[28][44]  ( .D(n5675), .CK(CLK), .QN(n63587) );
  DFF_X1 \REGISTERS_reg[28][43]  ( .D(n5674), .CK(CLK), .QN(n63588) );
  DFF_X1 \REGISTERS_reg[28][42]  ( .D(n5673), .CK(CLK), .QN(n63589) );
  DFF_X1 \REGISTERS_reg[28][41]  ( .D(n5672), .CK(CLK), .QN(n63590) );
  DFF_X1 \REGISTERS_reg[28][40]  ( .D(n5671), .CK(CLK), .QN(n63591) );
  DFF_X1 \REGISTERS_reg[28][39]  ( .D(n5670), .CK(CLK), .QN(n63592) );
  DFF_X1 \REGISTERS_reg[28][38]  ( .D(n5669), .CK(CLK), .QN(n63593) );
  DFF_X1 \REGISTERS_reg[28][37]  ( .D(n5668), .CK(CLK), .QN(n63594) );
  DFF_X1 \REGISTERS_reg[28][36]  ( .D(n5667), .CK(CLK), .QN(n63595) );
  DFF_X1 \REGISTERS_reg[28][35]  ( .D(n5666), .CK(CLK), .QN(n63596) );
  DFF_X1 \REGISTERS_reg[28][34]  ( .D(n5665), .CK(CLK), .QN(n63597) );
  DFF_X1 \REGISTERS_reg[28][33]  ( .D(n5664), .CK(CLK), .QN(n63598) );
  DFF_X1 \REGISTERS_reg[28][32]  ( .D(n5663), .CK(CLK), .QN(n63599) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n5662), .CK(CLK), .QN(n63600) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n5661), .CK(CLK), .QN(n63601) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n5660), .CK(CLK), .QN(n63602) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n5659), .CK(CLK), .QN(n63603) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n5658), .CK(CLK), .QN(n63604) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n5657), .CK(CLK), .QN(n63605) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n5656), .CK(CLK), .QN(n63606) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n5655), .CK(CLK), .QN(n63607) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n5654), .CK(CLK), .QN(n63608) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n5653), .CK(CLK), .QN(n63609) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n5652), .CK(CLK), .QN(n63610) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n5651), .CK(CLK), .QN(n63611) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n5650), .CK(CLK), .QN(n63612) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n5649), .CK(CLK), .QN(n63613) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n5648), .CK(CLK), .QN(n63614) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n5647), .CK(CLK), .QN(n63615) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n5646), .CK(CLK), .QN(n63616) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n5645), .CK(CLK), .QN(n63617) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n5644), .CK(CLK), .QN(n63618) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n5643), .CK(CLK), .QN(n63619) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n5642), .CK(CLK), .QN(n63620) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n5641), .CK(CLK), .QN(n63621) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n5640), .CK(CLK), .QN(n63622) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n5639), .CK(CLK), .QN(n63623) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n5638), .CK(CLK), .QN(n63624) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n5637), .CK(CLK), .QN(n63625) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n5636), .CK(CLK), .QN(n63626) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n5635), .CK(CLK), .QN(n63627) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n5634), .CK(CLK), .QN(n63628) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n5633), .CK(CLK), .QN(n63629) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n5632), .CK(CLK), .QN(n63630) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n5631), .CK(CLK), .QN(n63631) );
  DFF_X1 \REGISTERS_reg[27][59]  ( .D(n5754), .CK(CLK), .QN(n63506) );
  DFF_X1 \REGISTERS_reg[27][58]  ( .D(n5753), .CK(CLK), .QN(n63507) );
  DFF_X1 \REGISTERS_reg[27][57]  ( .D(n5752), .CK(CLK), .QN(n63508) );
  DFF_X1 \REGISTERS_reg[27][56]  ( .D(n5751), .CK(CLK), .QN(n63509) );
  DFF_X1 \REGISTERS_reg[27][55]  ( .D(n5750), .CK(CLK), .QN(n63510) );
  DFF_X1 \REGISTERS_reg[27][54]  ( .D(n5749), .CK(CLK), .QN(n63511) );
  DFF_X1 \REGISTERS_reg[27][53]  ( .D(n5748), .CK(CLK), .QN(n63512) );
  DFF_X1 \REGISTERS_reg[27][52]  ( .D(n5747), .CK(CLK), .QN(n63513) );
  DFF_X1 \REGISTERS_reg[27][51]  ( .D(n5746), .CK(CLK), .QN(n63514) );
  DFF_X1 \REGISTERS_reg[27][50]  ( .D(n5745), .CK(CLK), .QN(n63515) );
  DFF_X1 \REGISTERS_reg[27][49]  ( .D(n5744), .CK(CLK), .QN(n63516) );
  DFF_X1 \REGISTERS_reg[27][48]  ( .D(n5743), .CK(CLK), .QN(n63517) );
  DFF_X1 \REGISTERS_reg[27][47]  ( .D(n5742), .CK(CLK), .QN(n63518) );
  DFF_X1 \REGISTERS_reg[27][46]  ( .D(n5741), .CK(CLK), .QN(n63519) );
  DFF_X1 \REGISTERS_reg[27][45]  ( .D(n5740), .CK(CLK), .QN(n63520) );
  DFF_X1 \REGISTERS_reg[27][44]  ( .D(n5739), .CK(CLK), .QN(n63521) );
  DFF_X1 \REGISTERS_reg[27][43]  ( .D(n5738), .CK(CLK), .QN(n63522) );
  DFF_X1 \REGISTERS_reg[27][42]  ( .D(n5737), .CK(CLK), .QN(n63523) );
  DFF_X1 \REGISTERS_reg[27][41]  ( .D(n5736), .CK(CLK), .QN(n63524) );
  DFF_X1 \REGISTERS_reg[27][40]  ( .D(n5735), .CK(CLK), .QN(n63525) );
  DFF_X1 \REGISTERS_reg[27][39]  ( .D(n5734), .CK(CLK), .QN(n63526) );
  DFF_X1 \REGISTERS_reg[27][38]  ( .D(n5733), .CK(CLK), .QN(n63527) );
  DFF_X1 \REGISTERS_reg[27][37]  ( .D(n5732), .CK(CLK), .QN(n63528) );
  DFF_X1 \REGISTERS_reg[27][36]  ( .D(n5731), .CK(CLK), .QN(n63529) );
  DFF_X1 \REGISTERS_reg[27][35]  ( .D(n5730), .CK(CLK), .QN(n63530) );
  DFF_X1 \REGISTERS_reg[27][34]  ( .D(n5729), .CK(CLK), .QN(n63531) );
  DFF_X1 \REGISTERS_reg[27][33]  ( .D(n5728), .CK(CLK), .QN(n63532) );
  DFF_X1 \REGISTERS_reg[27][32]  ( .D(n5727), .CK(CLK), .QN(n63533) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n5726), .CK(CLK), .QN(n63534) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n5725), .CK(CLK), .QN(n63535) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n5724), .CK(CLK), .QN(n63536) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n5723), .CK(CLK), .QN(n63537) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n5722), .CK(CLK), .QN(n63538) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n5721), .CK(CLK), .QN(n63539) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n5720), .CK(CLK), .QN(n63540) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n5719), .CK(CLK), .QN(n63541) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n5718), .CK(CLK), .QN(n63542) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n5717), .CK(CLK), .QN(n63543) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n5716), .CK(CLK), .QN(n63544) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n5715), .CK(CLK), .QN(n63545) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n5714), .CK(CLK), .QN(n63546) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n5713), .CK(CLK), .QN(n63547) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n5712), .CK(CLK), .QN(n63548) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n5711), .CK(CLK), .QN(n63549) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n5710), .CK(CLK), .QN(n63550) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n5709), .CK(CLK), .QN(n63551) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n5708), .CK(CLK), .QN(n63552) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n5707), .CK(CLK), .QN(n63553) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n5706), .CK(CLK), .QN(n63554) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n5705), .CK(CLK), .QN(n63555) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n5704), .CK(CLK), .QN(n63556) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n5703), .CK(CLK), .QN(n63557) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n5702), .CK(CLK), .QN(n63558) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n5701), .CK(CLK), .QN(n63559) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n5700), .CK(CLK), .QN(n63560) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n5699), .CK(CLK), .QN(n63561) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n5698), .CK(CLK), .QN(n63562) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n5697), .CK(CLK), .QN(n63563) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n5696), .CK(CLK), .QN(n63564) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n5695), .CK(CLK), .QN(n63565) );
  DFF_X1 \REGISTERS_reg[25][59]  ( .D(n5882), .CK(CLK), .Q(n8967), .QN(n63435)
         );
  DFF_X1 \REGISTERS_reg[25][58]  ( .D(n5881), .CK(CLK), .Q(n8969), .QN(n63436)
         );
  DFF_X1 \REGISTERS_reg[25][57]  ( .D(n5880), .CK(CLK), .Q(n8971), .QN(n63437)
         );
  DFF_X1 \REGISTERS_reg[25][56]  ( .D(n5879), .CK(CLK), .Q(n8973), .QN(n63438)
         );
  DFF_X1 \REGISTERS_reg[25][55]  ( .D(n5878), .CK(CLK), .Q(n8975), .QN(n63439)
         );
  DFF_X1 \REGISTERS_reg[25][54]  ( .D(n5877), .CK(CLK), .Q(n8977), .QN(n63440)
         );
  DFF_X1 \REGISTERS_reg[25][53]  ( .D(n5876), .CK(CLK), .Q(n8979), .QN(n63441)
         );
  DFF_X1 \REGISTERS_reg[25][52]  ( .D(n5875), .CK(CLK), .Q(n8981), .QN(n63442)
         );
  DFF_X1 \REGISTERS_reg[25][51]  ( .D(n5874), .CK(CLK), .Q(n8983), .QN(n63443)
         );
  DFF_X1 \REGISTERS_reg[25][50]  ( .D(n5873), .CK(CLK), .Q(n8985), .QN(n63444)
         );
  DFF_X1 \REGISTERS_reg[25][49]  ( .D(n5872), .CK(CLK), .Q(n8987), .QN(n63445)
         );
  DFF_X1 \REGISTERS_reg[25][48]  ( .D(n5871), .CK(CLK), .Q(n8989), .QN(n63446)
         );
  DFF_X1 \REGISTERS_reg[25][47]  ( .D(n5870), .CK(CLK), .Q(n8991), .QN(n63447)
         );
  DFF_X1 \REGISTERS_reg[25][46]  ( .D(n5869), .CK(CLK), .Q(n8993), .QN(n63448)
         );
  DFF_X1 \REGISTERS_reg[25][45]  ( .D(n5868), .CK(CLK), .Q(n8995), .QN(n63449)
         );
  DFF_X1 \REGISTERS_reg[25][44]  ( .D(n5867), .CK(CLK), .Q(n8997), .QN(n63450)
         );
  DFF_X1 \REGISTERS_reg[25][43]  ( .D(n5866), .CK(CLK), .Q(n8999), .QN(n63451)
         );
  DFF_X1 \REGISTERS_reg[25][42]  ( .D(n5865), .CK(CLK), .Q(n9001), .QN(n63452)
         );
  DFF_X1 \REGISTERS_reg[25][41]  ( .D(n5864), .CK(CLK), .Q(n9003), .QN(n63453)
         );
  DFF_X1 \REGISTERS_reg[25][40]  ( .D(n5863), .CK(CLK), .Q(n9005), .QN(n63454)
         );
  DFF_X1 \REGISTERS_reg[25][39]  ( .D(n5862), .CK(CLK), .Q(n9007), .QN(n63455)
         );
  DFF_X1 \REGISTERS_reg[25][38]  ( .D(n5861), .CK(CLK), .Q(n9009), .QN(n63456)
         );
  DFF_X1 \REGISTERS_reg[25][37]  ( .D(n5860), .CK(CLK), .Q(n9011), .QN(n63457)
         );
  DFF_X1 \REGISTERS_reg[25][36]  ( .D(n5859), .CK(CLK), .Q(n9013), .QN(n63458)
         );
  DFF_X1 \REGISTERS_reg[25][35]  ( .D(n5858), .CK(CLK), .Q(n9015), .QN(n63459)
         );
  DFF_X1 \REGISTERS_reg[25][34]  ( .D(n5857), .CK(CLK), .Q(n9017), .QN(n63460)
         );
  DFF_X1 \REGISTERS_reg[25][33]  ( .D(n5856), .CK(CLK), .Q(n9019), .QN(n63461)
         );
  DFF_X1 \REGISTERS_reg[25][32]  ( .D(n5855), .CK(CLK), .Q(n9021), .QN(n63462)
         );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n5854), .CK(CLK), .Q(n9023), .QN(n63463)
         );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n5853), .CK(CLK), .Q(n9025), .QN(n63464)
         );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n5852), .CK(CLK), .Q(n9027), .QN(n63465)
         );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n5851), .CK(CLK), .Q(n9029), .QN(n63466)
         );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n5850), .CK(CLK), .Q(n9031), .QN(n63467)
         );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n5849), .CK(CLK), .Q(n9033), .QN(n63468)
         );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n5848), .CK(CLK), .Q(n9035), .QN(n63469)
         );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n5847), .CK(CLK), .Q(n9037), .QN(n63470)
         );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n5846), .CK(CLK), .Q(n9039), .QN(n63471)
         );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n5845), .CK(CLK), .Q(n9041), .QN(n63472)
         );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n5844), .CK(CLK), .Q(n9043), .QN(n63473)
         );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n5843), .CK(CLK), .Q(n9045), .QN(n63474)
         );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n5842), .CK(CLK), .Q(n9047), .QN(n63475)
         );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n5841), .CK(CLK), .Q(n9049), .QN(n63476)
         );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n5840), .CK(CLK), .Q(n9051), .QN(n63477)
         );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n5839), .CK(CLK), .Q(n9053), .QN(n63478)
         );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n5838), .CK(CLK), .Q(n9055), .QN(n63479)
         );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n5837), .CK(CLK), .Q(n9057), .QN(n63480)
         );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n5836), .CK(CLK), .Q(n9059), .QN(n63481)
         );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n5835), .CK(CLK), .Q(n9061), .QN(n63482)
         );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n5834), .CK(CLK), .Q(n9063), .QN(n63483)
         );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n5833), .CK(CLK), .Q(n9065), .QN(n63484)
         );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n5832), .CK(CLK), .Q(n9067), .QN(n63485)
         );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n5831), .CK(CLK), .Q(n9069), .QN(n63486)
         );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n5830), .CK(CLK), .Q(n9071), .QN(n63487)
         );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n5829), .CK(CLK), .Q(n9073), .QN(n63488)
         );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n5828), .CK(CLK), .Q(n9075), .QN(n63489)
         );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n5827), .CK(CLK), .Q(n9077), .QN(n63490)
         );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n5826), .CK(CLK), .Q(n9079), .QN(n63491)
         );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n5825), .CK(CLK), .Q(n9081), .QN(n63492)
         );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n5824), .CK(CLK), .Q(n9083), .QN(n63493)
         );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n5823), .CK(CLK), .Q(n9085), .QN(n63494)
         );
  DFF_X1 \REGISTERS_reg[23][59]  ( .D(n6010), .CK(CLK), .QN(n63302) );
  DFF_X1 \REGISTERS_reg[23][58]  ( .D(n6009), .CK(CLK), .QN(n63303) );
  DFF_X1 \REGISTERS_reg[23][57]  ( .D(n6008), .CK(CLK), .QN(n63304) );
  DFF_X1 \REGISTERS_reg[23][56]  ( .D(n6007), .CK(CLK), .QN(n63305) );
  DFF_X1 \REGISTERS_reg[23][55]  ( .D(n6006), .CK(CLK), .QN(n63306) );
  DFF_X1 \REGISTERS_reg[23][54]  ( .D(n6005), .CK(CLK), .QN(n63307) );
  DFF_X1 \REGISTERS_reg[23][53]  ( .D(n6004), .CK(CLK), .QN(n63308) );
  DFF_X1 \REGISTERS_reg[23][52]  ( .D(n6003), .CK(CLK), .QN(n63309) );
  DFF_X1 \REGISTERS_reg[23][51]  ( .D(n6002), .CK(CLK), .QN(n63310) );
  DFF_X1 \REGISTERS_reg[23][50]  ( .D(n6001), .CK(CLK), .QN(n63311) );
  DFF_X1 \REGISTERS_reg[23][49]  ( .D(n6000), .CK(CLK), .QN(n63312) );
  DFF_X1 \REGISTERS_reg[23][48]  ( .D(n5999), .CK(CLK), .QN(n63313) );
  DFF_X1 \REGISTERS_reg[23][47]  ( .D(n5998), .CK(CLK), .QN(n63314) );
  DFF_X1 \REGISTERS_reg[23][46]  ( .D(n5997), .CK(CLK), .QN(n63315) );
  DFF_X1 \REGISTERS_reg[23][45]  ( .D(n5996), .CK(CLK), .QN(n63316) );
  DFF_X1 \REGISTERS_reg[23][44]  ( .D(n5995), .CK(CLK), .QN(n63317) );
  DFF_X1 \REGISTERS_reg[23][43]  ( .D(n5994), .CK(CLK), .QN(n63318) );
  DFF_X1 \REGISTERS_reg[23][42]  ( .D(n5993), .CK(CLK), .QN(n63319) );
  DFF_X1 \REGISTERS_reg[23][41]  ( .D(n5992), .CK(CLK), .QN(n63320) );
  DFF_X1 \REGISTERS_reg[23][40]  ( .D(n5991), .CK(CLK), .QN(n63321) );
  DFF_X1 \REGISTERS_reg[23][39]  ( .D(n5990), .CK(CLK), .QN(n63322) );
  DFF_X1 \REGISTERS_reg[23][38]  ( .D(n5989), .CK(CLK), .QN(n63323) );
  DFF_X1 \REGISTERS_reg[23][37]  ( .D(n5988), .CK(CLK), .QN(n63324) );
  DFF_X1 \REGISTERS_reg[23][36]  ( .D(n5987), .CK(CLK), .QN(n63325) );
  DFF_X1 \REGISTERS_reg[23][35]  ( .D(n5986), .CK(CLK), .QN(n63326) );
  DFF_X1 \REGISTERS_reg[23][34]  ( .D(n5985), .CK(CLK), .QN(n63327) );
  DFF_X1 \REGISTERS_reg[23][33]  ( .D(n5984), .CK(CLK), .QN(n63328) );
  DFF_X1 \REGISTERS_reg[23][32]  ( .D(n5983), .CK(CLK), .QN(n63329) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n5982), .CK(CLK), .QN(n63330) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n5981), .CK(CLK), .QN(n63331) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n5980), .CK(CLK), .QN(n63332) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n5979), .CK(CLK), .QN(n63333) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n5978), .CK(CLK), .QN(n63334) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n5977), .CK(CLK), .QN(n63335) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n5976), .CK(CLK), .QN(n63336) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n5975), .CK(CLK), .QN(n63337) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n5974), .CK(CLK), .QN(n63338) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n5973), .CK(CLK), .QN(n63339) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n5972), .CK(CLK), .QN(n63340) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n5971), .CK(CLK), .QN(n63341) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n5970), .CK(CLK), .QN(n63342) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n5969), .CK(CLK), .QN(n63343) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n5968), .CK(CLK), .QN(n63344) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n5967), .CK(CLK), .QN(n63345) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n5966), .CK(CLK), .QN(n63346) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n5965), .CK(CLK), .QN(n63347) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n5964), .CK(CLK), .QN(n63348) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n5963), .CK(CLK), .QN(n63349) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n5962), .CK(CLK), .QN(n63350) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n5961), .CK(CLK), .QN(n63351) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n5960), .CK(CLK), .QN(n63352) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n5959), .CK(CLK), .QN(n63353) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n5958), .CK(CLK), .QN(n63354) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n5957), .CK(CLK), .QN(n63355) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n5956), .CK(CLK), .QN(n63356) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n5955), .CK(CLK), .QN(n63357) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n5954), .CK(CLK), .QN(n63358) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n5953), .CK(CLK), .QN(n63359) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n5952), .CK(CLK), .QN(n63360) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n5951), .CK(CLK), .QN(n63361) );
  DFF_X1 \REGISTERS_reg[19][59]  ( .D(n6266), .CK(CLK), .QN(n63101) );
  DFF_X1 \REGISTERS_reg[19][58]  ( .D(n6265), .CK(CLK), .QN(n63102) );
  DFF_X1 \REGISTERS_reg[19][57]  ( .D(n6264), .CK(CLK), .QN(n63103) );
  DFF_X1 \REGISTERS_reg[19][56]  ( .D(n6263), .CK(CLK), .QN(n63104) );
  DFF_X1 \REGISTERS_reg[19][55]  ( .D(n6262), .CK(CLK), .QN(n63105) );
  DFF_X1 \REGISTERS_reg[19][54]  ( .D(n6261), .CK(CLK), .QN(n63106) );
  DFF_X1 \REGISTERS_reg[19][53]  ( .D(n6260), .CK(CLK), .QN(n63107) );
  DFF_X1 \REGISTERS_reg[19][52]  ( .D(n6259), .CK(CLK), .QN(n63108) );
  DFF_X1 \REGISTERS_reg[19][51]  ( .D(n6258), .CK(CLK), .QN(n63109) );
  DFF_X1 \REGISTERS_reg[19][50]  ( .D(n6257), .CK(CLK), .QN(n63110) );
  DFF_X1 \REGISTERS_reg[19][49]  ( .D(n6256), .CK(CLK), .QN(n63111) );
  DFF_X1 \REGISTERS_reg[19][48]  ( .D(n6255), .CK(CLK), .QN(n63112) );
  DFF_X1 \REGISTERS_reg[19][47]  ( .D(n6254), .CK(CLK), .QN(n63113) );
  DFF_X1 \REGISTERS_reg[19][46]  ( .D(n6253), .CK(CLK), .QN(n63114) );
  DFF_X1 \REGISTERS_reg[19][45]  ( .D(n6252), .CK(CLK), .QN(n63115) );
  DFF_X1 \REGISTERS_reg[19][44]  ( .D(n6251), .CK(CLK), .QN(n63116) );
  DFF_X1 \REGISTERS_reg[19][43]  ( .D(n6250), .CK(CLK), .QN(n63117) );
  DFF_X1 \REGISTERS_reg[19][42]  ( .D(n6249), .CK(CLK), .QN(n63118) );
  DFF_X1 \REGISTERS_reg[19][41]  ( .D(n6248), .CK(CLK), .QN(n63119) );
  DFF_X1 \REGISTERS_reg[19][40]  ( .D(n6247), .CK(CLK), .QN(n63120) );
  DFF_X1 \REGISTERS_reg[19][39]  ( .D(n6246), .CK(CLK), .QN(n63121) );
  DFF_X1 \REGISTERS_reg[19][38]  ( .D(n6245), .CK(CLK), .QN(n63122) );
  DFF_X1 \REGISTERS_reg[19][37]  ( .D(n6244), .CK(CLK), .QN(n63123) );
  DFF_X1 \REGISTERS_reg[19][36]  ( .D(n6243), .CK(CLK), .QN(n63124) );
  DFF_X1 \REGISTERS_reg[19][35]  ( .D(n6242), .CK(CLK), .QN(n63125) );
  DFF_X1 \REGISTERS_reg[19][34]  ( .D(n6241), .CK(CLK), .QN(n63126) );
  DFF_X1 \REGISTERS_reg[19][33]  ( .D(n6240), .CK(CLK), .QN(n63127) );
  DFF_X1 \REGISTERS_reg[19][32]  ( .D(n6239), .CK(CLK), .QN(n63128) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n6238), .CK(CLK), .QN(n63129) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n6237), .CK(CLK), .QN(n63130) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n6236), .CK(CLK), .QN(n63131) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n6235), .CK(CLK), .QN(n63132) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n6234), .CK(CLK), .QN(n63133) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n6233), .CK(CLK), .QN(n63134) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n6232), .CK(CLK), .QN(n63135) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n6231), .CK(CLK), .QN(n63136) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n6230), .CK(CLK), .QN(n63137) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n6229), .CK(CLK), .QN(n63138) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n6228), .CK(CLK), .QN(n63139) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n6227), .CK(CLK), .QN(n63140) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n6226), .CK(CLK), .QN(n63141) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n6225), .CK(CLK), .QN(n63142) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n6224), .CK(CLK), .QN(n63143) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n6223), .CK(CLK), .QN(n63144) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n6222), .CK(CLK), .QN(n63145) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n6221), .CK(CLK), .QN(n63146) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n6220), .CK(CLK), .QN(n63147) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n6219), .CK(CLK), .QN(n63148) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n6218), .CK(CLK), .QN(n63149) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n6217), .CK(CLK), .QN(n63150) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n6216), .CK(CLK), .QN(n63151) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n6215), .CK(CLK), .QN(n63152) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n6214), .CK(CLK), .QN(n63153) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n6213), .CK(CLK), .QN(n63154) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n6212), .CK(CLK), .QN(n63155) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n6211), .CK(CLK), .QN(n63156) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n6210), .CK(CLK), .QN(n63157) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n6209), .CK(CLK), .QN(n63158) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n6208), .CK(CLK), .QN(n63159) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n6207), .CK(CLK), .QN(n63160) );
  DFF_X1 \REGISTERS_reg[24][59]  ( .D(n5946), .CK(CLK), .QN(n63368) );
  DFF_X1 \REGISTERS_reg[24][58]  ( .D(n5945), .CK(CLK), .QN(n63369) );
  DFF_X1 \REGISTERS_reg[24][57]  ( .D(n5944), .CK(CLK), .QN(n63370) );
  DFF_X1 \REGISTERS_reg[24][56]  ( .D(n5943), .CK(CLK), .QN(n63371) );
  DFF_X1 \REGISTERS_reg[24][55]  ( .D(n5942), .CK(CLK), .QN(n63372) );
  DFF_X1 \REGISTERS_reg[24][54]  ( .D(n5941), .CK(CLK), .QN(n63373) );
  DFF_X1 \REGISTERS_reg[24][53]  ( .D(n5940), .CK(CLK), .QN(n63374) );
  DFF_X1 \REGISTERS_reg[24][52]  ( .D(n5939), .CK(CLK), .QN(n63375) );
  DFF_X1 \REGISTERS_reg[24][51]  ( .D(n5938), .CK(CLK), .QN(n63376) );
  DFF_X1 \REGISTERS_reg[24][50]  ( .D(n5937), .CK(CLK), .QN(n63377) );
  DFF_X1 \REGISTERS_reg[24][49]  ( .D(n5936), .CK(CLK), .QN(n63378) );
  DFF_X1 \REGISTERS_reg[24][48]  ( .D(n5935), .CK(CLK), .QN(n63379) );
  DFF_X1 \REGISTERS_reg[24][47]  ( .D(n5934), .CK(CLK), .QN(n63380) );
  DFF_X1 \REGISTERS_reg[24][46]  ( .D(n5933), .CK(CLK), .QN(n63381) );
  DFF_X1 \REGISTERS_reg[24][45]  ( .D(n5932), .CK(CLK), .QN(n63382) );
  DFF_X1 \REGISTERS_reg[24][44]  ( .D(n5931), .CK(CLK), .QN(n63383) );
  DFF_X1 \REGISTERS_reg[24][43]  ( .D(n5930), .CK(CLK), .QN(n63384) );
  DFF_X1 \REGISTERS_reg[24][42]  ( .D(n5929), .CK(CLK), .QN(n63385) );
  DFF_X1 \REGISTERS_reg[24][41]  ( .D(n5928), .CK(CLK), .QN(n63386) );
  DFF_X1 \REGISTERS_reg[24][40]  ( .D(n5927), .CK(CLK), .QN(n63387) );
  DFF_X1 \REGISTERS_reg[24][39]  ( .D(n5926), .CK(CLK), .QN(n63388) );
  DFF_X1 \REGISTERS_reg[24][38]  ( .D(n5925), .CK(CLK), .QN(n63389) );
  DFF_X1 \REGISTERS_reg[24][37]  ( .D(n5924), .CK(CLK), .QN(n63390) );
  DFF_X1 \REGISTERS_reg[24][36]  ( .D(n5923), .CK(CLK), .QN(n63391) );
  DFF_X1 \REGISTERS_reg[24][35]  ( .D(n5922), .CK(CLK), .QN(n63392) );
  DFF_X1 \REGISTERS_reg[24][34]  ( .D(n5921), .CK(CLK), .QN(n63393) );
  DFF_X1 \REGISTERS_reg[24][33]  ( .D(n5920), .CK(CLK), .QN(n63394) );
  DFF_X1 \REGISTERS_reg[24][32]  ( .D(n5919), .CK(CLK), .QN(n63395) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n5918), .CK(CLK), .QN(n63396) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n5917), .CK(CLK), .QN(n63397) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n5916), .CK(CLK), .QN(n63398) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n5915), .CK(CLK), .QN(n63399) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n5914), .CK(CLK), .QN(n63400) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n5913), .CK(CLK), .QN(n63401) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n5912), .CK(CLK), .QN(n63402) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n5911), .CK(CLK), .QN(n63403) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n5910), .CK(CLK), .QN(n63404) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n5909), .CK(CLK), .QN(n63405) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n5908), .CK(CLK), .QN(n63406) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n5907), .CK(CLK), .QN(n63407) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n5906), .CK(CLK), .QN(n63408) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n5905), .CK(CLK), .QN(n63409) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n5904), .CK(CLK), .QN(n63410) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n5903), .CK(CLK), .QN(n63411) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n5902), .CK(CLK), .QN(n63412) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n5901), .CK(CLK), .QN(n63413) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n5900), .CK(CLK), .QN(n63414) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n5899), .CK(CLK), .QN(n63415) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n5898), .CK(CLK), .QN(n63416) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n5897), .CK(CLK), .QN(n63417) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n5896), .CK(CLK), .QN(n63418) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n5895), .CK(CLK), .QN(n63419) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n5894), .CK(CLK), .QN(n63420) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n5893), .CK(CLK), .QN(n63421) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n5892), .CK(CLK), .QN(n63422) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n5891), .CK(CLK), .QN(n63423) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n5890), .CK(CLK), .QN(n63424) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n5889), .CK(CLK), .QN(n63425) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n5888), .CK(CLK), .QN(n63426) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n5887), .CK(CLK), .QN(n63427) );
  DFF_X1 \REGISTERS_reg[17][59]  ( .D(n6394), .CK(CLK), .Q(n58229), .QN(n63032) );
  DFF_X1 \REGISTERS_reg[17][58]  ( .D(n6393), .CK(CLK), .Q(n58227), .QN(n63033) );
  DFF_X1 \REGISTERS_reg[17][57]  ( .D(n6392), .CK(CLK), .Q(n58225), .QN(n63034) );
  DFF_X1 \REGISTERS_reg[17][56]  ( .D(n6391), .CK(CLK), .Q(n58223), .QN(n63035) );
  DFF_X1 \REGISTERS_reg[17][55]  ( .D(n6390), .CK(CLK), .Q(n58221), .QN(n63036) );
  DFF_X1 \REGISTERS_reg[17][54]  ( .D(n6389), .CK(CLK), .Q(n58219), .QN(n63037) );
  DFF_X1 \REGISTERS_reg[17][53]  ( .D(n6388), .CK(CLK), .Q(n58217), .QN(n63038) );
  DFF_X1 \REGISTERS_reg[17][52]  ( .D(n6387), .CK(CLK), .Q(n58215), .QN(n63039) );
  DFF_X1 \REGISTERS_reg[17][51]  ( .D(n6386), .CK(CLK), .Q(n58213), .QN(n63040) );
  DFF_X1 \REGISTERS_reg[17][50]  ( .D(n6385), .CK(CLK), .Q(n58211), .QN(n63041) );
  DFF_X1 \REGISTERS_reg[17][49]  ( .D(n6384), .CK(CLK), .Q(n58209), .QN(n63042) );
  DFF_X1 \REGISTERS_reg[17][48]  ( .D(n6383), .CK(CLK), .Q(n58207), .QN(n63043) );
  DFF_X1 \REGISTERS_reg[17][47]  ( .D(n6382), .CK(CLK), .Q(n58205), .QN(n63044) );
  DFF_X1 \REGISTERS_reg[17][46]  ( .D(n6381), .CK(CLK), .Q(n58203), .QN(n63045) );
  DFF_X1 \REGISTERS_reg[17][45]  ( .D(n6380), .CK(CLK), .Q(n58201), .QN(n63046) );
  DFF_X1 \REGISTERS_reg[17][44]  ( .D(n6379), .CK(CLK), .Q(n58199), .QN(n63047) );
  DFF_X1 \REGISTERS_reg[17][43]  ( .D(n6378), .CK(CLK), .Q(n58197), .QN(n63048) );
  DFF_X1 \REGISTERS_reg[17][42]  ( .D(n6377), .CK(CLK), .Q(n58195), .QN(n63049) );
  DFF_X1 \REGISTERS_reg[17][41]  ( .D(n6376), .CK(CLK), .Q(n58193), .QN(n63050) );
  DFF_X1 \REGISTERS_reg[17][40]  ( .D(n6375), .CK(CLK), .Q(n58191), .QN(n63051) );
  DFF_X1 \REGISTERS_reg[17][39]  ( .D(n6374), .CK(CLK), .Q(n58189), .QN(n63052) );
  DFF_X1 \REGISTERS_reg[17][38]  ( .D(n6373), .CK(CLK), .Q(n58187), .QN(n63053) );
  DFF_X1 \REGISTERS_reg[17][37]  ( .D(n6372), .CK(CLK), .Q(n58185), .QN(n63054) );
  DFF_X1 \REGISTERS_reg[17][36]  ( .D(n6371), .CK(CLK), .Q(n58183), .QN(n63055) );
  DFF_X1 \REGISTERS_reg[17][35]  ( .D(n6370), .CK(CLK), .Q(n58181), .QN(n63056) );
  DFF_X1 \REGISTERS_reg[17][34]  ( .D(n6369), .CK(CLK), .Q(n58179), .QN(n63057) );
  DFF_X1 \REGISTERS_reg[17][33]  ( .D(n6368), .CK(CLK), .Q(n58177), .QN(n63058) );
  DFF_X1 \REGISTERS_reg[17][32]  ( .D(n6367), .CK(CLK), .Q(n58175), .QN(n63059) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n6366), .CK(CLK), .Q(n58173), .QN(n63060) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n6365), .CK(CLK), .Q(n58171), .QN(n63061) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n6364), .CK(CLK), .Q(n58169), .QN(n63062) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n6363), .CK(CLK), .Q(n58167), .QN(n63063) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n6362), .CK(CLK), .Q(n58165), .QN(n63064) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n6361), .CK(CLK), .Q(n58163), .QN(n63065) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n6360), .CK(CLK), .Q(n58161), .QN(n63066) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n6359), .CK(CLK), .Q(n58159), .QN(n63067) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n6358), .CK(CLK), .Q(n58157), .QN(n63068) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n6357), .CK(CLK), .Q(n58155), .QN(n63069) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n6356), .CK(CLK), .Q(n58153), .QN(n63070) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n6355), .CK(CLK), .Q(n58151), .QN(n63071) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n6354), .CK(CLK), .Q(n58149), .QN(n63072) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n6353), .CK(CLK), .Q(n58147), .QN(n63073) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n6352), .CK(CLK), .Q(n58145), .QN(n63074) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n6351), .CK(CLK), .Q(n58143), .QN(n63075) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n6350), .CK(CLK), .Q(n58141), .QN(n63076) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n6349), .CK(CLK), .Q(n58139), .QN(n63077) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n6348), .CK(CLK), .Q(n58137), .QN(n63078) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n6347), .CK(CLK), .Q(n58135), .QN(n63079) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n6346), .CK(CLK), .Q(n58134), .QN(n63080) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n6345), .CK(CLK), .Q(n58132), .QN(n63081) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n6344), .CK(CLK), .Q(n58130), .QN(n63082)
         );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n6343), .CK(CLK), .Q(n58128), .QN(n63083)
         );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n6342), .CK(CLK), .Q(n58126), .QN(n63084)
         );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n6341), .CK(CLK), .Q(n58124), .QN(n63085)
         );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n6340), .CK(CLK), .Q(n58122), .QN(n63086)
         );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n6339), .CK(CLK), .Q(n58120), .QN(n63087)
         );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n6338), .CK(CLK), .Q(n58118), .QN(n63088)
         );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n6337), .CK(CLK), .Q(n58116), .QN(n63089)
         );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n6336), .CK(CLK), .Q(n58114), .QN(n63090)
         );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n6335), .CK(CLK), .Q(n58112), .QN(n63091)
         );
  DFF_X1 \REGISTERS_reg[16][59]  ( .D(n6458), .CK(CLK), .Q(n58498), .QN(n62965) );
  DFF_X1 \REGISTERS_reg[16][58]  ( .D(n6457), .CK(CLK), .Q(n58497), .QN(n62966) );
  DFF_X1 \REGISTERS_reg[16][57]  ( .D(n6456), .CK(CLK), .Q(n58496), .QN(n62967) );
  DFF_X1 \REGISTERS_reg[16][56]  ( .D(n6455), .CK(CLK), .Q(n58495), .QN(n62968) );
  DFF_X1 \REGISTERS_reg[16][55]  ( .D(n6454), .CK(CLK), .Q(n58494), .QN(n62969) );
  DFF_X1 \REGISTERS_reg[16][54]  ( .D(n6453), .CK(CLK), .Q(n58493), .QN(n62970) );
  DFF_X1 \REGISTERS_reg[16][53]  ( .D(n6452), .CK(CLK), .Q(n58492), .QN(n62971) );
  DFF_X1 \REGISTERS_reg[16][52]  ( .D(n6451), .CK(CLK), .Q(n58491), .QN(n62972) );
  DFF_X1 \REGISTERS_reg[16][51]  ( .D(n6450), .CK(CLK), .Q(n58490), .QN(n62973) );
  DFF_X1 \REGISTERS_reg[16][50]  ( .D(n6449), .CK(CLK), .Q(n58489), .QN(n62974) );
  DFF_X1 \REGISTERS_reg[16][49]  ( .D(n6448), .CK(CLK), .Q(n58488), .QN(n62975) );
  DFF_X1 \REGISTERS_reg[16][48]  ( .D(n6447), .CK(CLK), .Q(n58487), .QN(n62976) );
  DFF_X1 \REGISTERS_reg[16][47]  ( .D(n6446), .CK(CLK), .Q(n58486), .QN(n62977) );
  DFF_X1 \REGISTERS_reg[16][46]  ( .D(n6445), .CK(CLK), .Q(n58485), .QN(n62978) );
  DFF_X1 \REGISTERS_reg[16][45]  ( .D(n6444), .CK(CLK), .Q(n58484), .QN(n62979) );
  DFF_X1 \REGISTERS_reg[16][44]  ( .D(n6443), .CK(CLK), .Q(n58483), .QN(n62980) );
  DFF_X1 \REGISTERS_reg[16][43]  ( .D(n6442), .CK(CLK), .Q(n58482), .QN(n62981) );
  DFF_X1 \REGISTERS_reg[16][42]  ( .D(n6441), .CK(CLK), .Q(n58481), .QN(n62982) );
  DFF_X1 \REGISTERS_reg[16][41]  ( .D(n6440), .CK(CLK), .Q(n58480), .QN(n62983) );
  DFF_X1 \REGISTERS_reg[16][40]  ( .D(n6439), .CK(CLK), .Q(n58479), .QN(n62984) );
  DFF_X1 \REGISTERS_reg[16][39]  ( .D(n6438), .CK(CLK), .Q(n58478), .QN(n62985) );
  DFF_X1 \REGISTERS_reg[16][38]  ( .D(n6437), .CK(CLK), .Q(n58477), .QN(n62986) );
  DFF_X1 \REGISTERS_reg[16][37]  ( .D(n6436), .CK(CLK), .Q(n58476), .QN(n62987) );
  DFF_X1 \REGISTERS_reg[16][36]  ( .D(n6435), .CK(CLK), .Q(n58475), .QN(n62988) );
  DFF_X1 \REGISTERS_reg[16][35]  ( .D(n6434), .CK(CLK), .Q(n58474), .QN(n62989) );
  DFF_X1 \REGISTERS_reg[16][34]  ( .D(n6433), .CK(CLK), .Q(n58473), .QN(n62990) );
  DFF_X1 \REGISTERS_reg[16][33]  ( .D(n6432), .CK(CLK), .Q(n58472), .QN(n62991) );
  DFF_X1 \REGISTERS_reg[16][32]  ( .D(n6431), .CK(CLK), .Q(n58471), .QN(n62992) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n6430), .CK(CLK), .Q(n58470), .QN(n62993) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n6429), .CK(CLK), .Q(n58469), .QN(n62994) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n6428), .CK(CLK), .Q(n58468), .QN(n62995) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n6427), .CK(CLK), .Q(n58467), .QN(n62996) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n6426), .CK(CLK), .Q(n58466), .QN(n62997) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n6425), .CK(CLK), .Q(n58465), .QN(n62998) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n6424), .CK(CLK), .Q(n58464), .QN(n62999) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n6423), .CK(CLK), .Q(n58463), .QN(n63000) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n6422), .CK(CLK), .Q(n58462), .QN(n63001) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n6421), .CK(CLK), .Q(n58461), .QN(n63002) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n6420), .CK(CLK), .Q(n58460), .QN(n63003) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n6419), .CK(CLK), .Q(n58459), .QN(n63004) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n6418), .CK(CLK), .Q(n58458), .QN(n63005) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n6417), .CK(CLK), .Q(n58457), .QN(n63006) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n6416), .CK(CLK), .Q(n58456), .QN(n63007) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n6415), .CK(CLK), .Q(n58455), .QN(n63008) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n6414), .CK(CLK), .Q(n58454), .QN(n63009) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n6413), .CK(CLK), .Q(n58453), .QN(n63010) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n6412), .CK(CLK), .Q(n58452), .QN(n63011) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n6411), .CK(CLK), .Q(n58451), .QN(n63012) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n6410), .CK(CLK), .Q(n58450), .QN(n63013) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n6409), .CK(CLK), .Q(n58449), .QN(n63014) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n6408), .CK(CLK), .Q(n58448), .QN(n63015)
         );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n6407), .CK(CLK), .Q(n58447), .QN(n63016)
         );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n6406), .CK(CLK), .Q(n58446), .QN(n63017)
         );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n6405), .CK(CLK), .Q(n58445), .QN(n63018)
         );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n6404), .CK(CLK), .Q(n58444), .QN(n63019)
         );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n6403), .CK(CLK), .Q(n58443), .QN(n63020)
         );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n6402), .CK(CLK), .Q(n58442), .QN(n63021)
         );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n6401), .CK(CLK), .Q(n58441), .QN(n63022)
         );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n6400), .CK(CLK), .Q(n58440), .QN(n63023)
         );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n6399), .CK(CLK), .Q(n58439), .QN(n63024)
         );
  DFF_X1 \REGISTERS_reg[22][59]  ( .D(n6074), .CK(CLK), .Q(n58714), .QN(n63235) );
  DFF_X1 \REGISTERS_reg[22][58]  ( .D(n6073), .CK(CLK), .Q(n58713), .QN(n63236) );
  DFF_X1 \REGISTERS_reg[22][57]  ( .D(n6072), .CK(CLK), .Q(n58712), .QN(n63237) );
  DFF_X1 \REGISTERS_reg[22][56]  ( .D(n6071), .CK(CLK), .Q(n58711), .QN(n63238) );
  DFF_X1 \REGISTERS_reg[22][55]  ( .D(n6070), .CK(CLK), .Q(n58710), .QN(n63239) );
  DFF_X1 \REGISTERS_reg[22][54]  ( .D(n6069), .CK(CLK), .Q(n58709), .QN(n63240) );
  DFF_X1 \REGISTERS_reg[22][53]  ( .D(n6068), .CK(CLK), .Q(n58708), .QN(n63241) );
  DFF_X1 \REGISTERS_reg[22][52]  ( .D(n6067), .CK(CLK), .Q(n58707), .QN(n63242) );
  DFF_X1 \REGISTERS_reg[22][51]  ( .D(n6066), .CK(CLK), .Q(n58706), .QN(n63243) );
  DFF_X1 \REGISTERS_reg[22][50]  ( .D(n6065), .CK(CLK), .Q(n58705), .QN(n63244) );
  DFF_X1 \REGISTERS_reg[22][49]  ( .D(n6064), .CK(CLK), .Q(n58704), .QN(n63245) );
  DFF_X1 \REGISTERS_reg[22][48]  ( .D(n6063), .CK(CLK), .Q(n58703), .QN(n63246) );
  DFF_X1 \REGISTERS_reg[22][47]  ( .D(n6062), .CK(CLK), .Q(n58702), .QN(n63247) );
  DFF_X1 \REGISTERS_reg[22][46]  ( .D(n6061), .CK(CLK), .Q(n58701), .QN(n63248) );
  DFF_X1 \REGISTERS_reg[22][45]  ( .D(n6060), .CK(CLK), .Q(n58700), .QN(n63249) );
  DFF_X1 \REGISTERS_reg[22][44]  ( .D(n6059), .CK(CLK), .Q(n58699), .QN(n63250) );
  DFF_X1 \REGISTERS_reg[22][43]  ( .D(n6058), .CK(CLK), .Q(n58698), .QN(n63251) );
  DFF_X1 \REGISTERS_reg[22][42]  ( .D(n6057), .CK(CLK), .Q(n58697), .QN(n63252) );
  DFF_X1 \REGISTERS_reg[22][41]  ( .D(n6056), .CK(CLK), .Q(n58696), .QN(n63253) );
  DFF_X1 \REGISTERS_reg[22][40]  ( .D(n6055), .CK(CLK), .Q(n58695), .QN(n63254) );
  DFF_X1 \REGISTERS_reg[22][39]  ( .D(n6054), .CK(CLK), .Q(n58694), .QN(n63255) );
  DFF_X1 \REGISTERS_reg[22][38]  ( .D(n6053), .CK(CLK), .Q(n58693), .QN(n63256) );
  DFF_X1 \REGISTERS_reg[22][37]  ( .D(n6052), .CK(CLK), .Q(n58692), .QN(n63257) );
  DFF_X1 \REGISTERS_reg[22][36]  ( .D(n6051), .CK(CLK), .Q(n58691), .QN(n63258) );
  DFF_X1 \REGISTERS_reg[22][35]  ( .D(n6050), .CK(CLK), .Q(n58690), .QN(n63259) );
  DFF_X1 \REGISTERS_reg[22][34]  ( .D(n6049), .CK(CLK), .Q(n58689), .QN(n63260) );
  DFF_X1 \REGISTERS_reg[22][33]  ( .D(n6048), .CK(CLK), .Q(n58688), .QN(n63261) );
  DFF_X1 \REGISTERS_reg[22][32]  ( .D(n6047), .CK(CLK), .Q(n58687), .QN(n63262) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n6046), .CK(CLK), .Q(n58686), .QN(n63263) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n6045), .CK(CLK), .Q(n58685), .QN(n63264) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n6044), .CK(CLK), .Q(n58684), .QN(n63265) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n6043), .CK(CLK), .Q(n58683), .QN(n63266) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n6042), .CK(CLK), .Q(n58682), .QN(n63267) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n6041), .CK(CLK), .Q(n58681), .QN(n63268) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n6040), .CK(CLK), .Q(n58680), .QN(n63269) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n6039), .CK(CLK), .Q(n58679), .QN(n63270) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n6038), .CK(CLK), .Q(n58678), .QN(n63271) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n6037), .CK(CLK), .Q(n58677), .QN(n63272) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n6036), .CK(CLK), .Q(n58676), .QN(n63273) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n6035), .CK(CLK), .Q(n58675), .QN(n63274) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n6034), .CK(CLK), .Q(n58674), .QN(n63275) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n6033), .CK(CLK), .Q(n58673), .QN(n63276) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n6032), .CK(CLK), .Q(n58672), .QN(n63277) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n6031), .CK(CLK), .Q(n58671), .QN(n63278) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n6030), .CK(CLK), .Q(n58670), .QN(n63279) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n6029), .CK(CLK), .Q(n58669), .QN(n63280) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n6028), .CK(CLK), .Q(n58668), .QN(n63281) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n6027), .CK(CLK), .Q(n58667), .QN(n63282) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n6026), .CK(CLK), .Q(n58742), .QN(n63283) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n6025), .CK(CLK), .Q(n58741), .QN(n63284) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n6024), .CK(CLK), .Q(n58740), .QN(n63285)
         );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n6023), .CK(CLK), .Q(n58739), .QN(n63286)
         );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n6022), .CK(CLK), .Q(n58738), .QN(n63287)
         );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n6021), .CK(CLK), .Q(n58737), .QN(n63288)
         );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n6020), .CK(CLK), .Q(n58736), .QN(n63289)
         );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n6019), .CK(CLK), .Q(n58735), .QN(n63290)
         );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n6018), .CK(CLK), .Q(n58734), .QN(n63291)
         );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n6017), .CK(CLK), .Q(n58733), .QN(n63292)
         );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n6016), .CK(CLK), .Q(n58732), .QN(n63293)
         );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n6015), .CK(CLK), .Q(n58731), .QN(n63294)
         );
  DFF_X1 \REGISTERS_reg[20][59]  ( .D(n6202), .CK(CLK), .Q(n58282), .QN(n63167) );
  DFF_X1 \REGISTERS_reg[20][58]  ( .D(n6201), .CK(CLK), .Q(n58281), .QN(n63168) );
  DFF_X1 \REGISTERS_reg[20][57]  ( .D(n6200), .CK(CLK), .Q(n58280), .QN(n63169) );
  DFF_X1 \REGISTERS_reg[20][56]  ( .D(n6199), .CK(CLK), .Q(n58279), .QN(n63170) );
  DFF_X1 \REGISTERS_reg[20][55]  ( .D(n6198), .CK(CLK), .Q(n58278), .QN(n63171) );
  DFF_X1 \REGISTERS_reg[20][54]  ( .D(n6197), .CK(CLK), .Q(n58277), .QN(n63172) );
  DFF_X1 \REGISTERS_reg[20][53]  ( .D(n6196), .CK(CLK), .Q(n58276), .QN(n63173) );
  DFF_X1 \REGISTERS_reg[20][52]  ( .D(n6195), .CK(CLK), .Q(n58275), .QN(n63174) );
  DFF_X1 \REGISTERS_reg[20][51]  ( .D(n6194), .CK(CLK), .Q(n58274), .QN(n63175) );
  DFF_X1 \REGISTERS_reg[20][50]  ( .D(n6193), .CK(CLK), .Q(n58273), .QN(n63176) );
  DFF_X1 \REGISTERS_reg[20][49]  ( .D(n6192), .CK(CLK), .Q(n58272), .QN(n63177) );
  DFF_X1 \REGISTERS_reg[20][48]  ( .D(n6191), .CK(CLK), .Q(n58271), .QN(n63178) );
  DFF_X1 \REGISTERS_reg[20][47]  ( .D(n6190), .CK(CLK), .Q(n58270), .QN(n63179) );
  DFF_X1 \REGISTERS_reg[20][46]  ( .D(n6189), .CK(CLK), .Q(n58269), .QN(n63180) );
  DFF_X1 \REGISTERS_reg[20][45]  ( .D(n6188), .CK(CLK), .Q(n58268), .QN(n63181) );
  DFF_X1 \REGISTERS_reg[20][44]  ( .D(n6187), .CK(CLK), .Q(n58267), .QN(n63182) );
  DFF_X1 \REGISTERS_reg[20][43]  ( .D(n6186), .CK(CLK), .Q(n58266), .QN(n63183) );
  DFF_X1 \REGISTERS_reg[20][42]  ( .D(n6185), .CK(CLK), .Q(n58265), .QN(n63184) );
  DFF_X1 \REGISTERS_reg[20][41]  ( .D(n6184), .CK(CLK), .Q(n58264), .QN(n63185) );
  DFF_X1 \REGISTERS_reg[20][40]  ( .D(n6183), .CK(CLK), .Q(n58263), .QN(n63186) );
  DFF_X1 \REGISTERS_reg[20][39]  ( .D(n6182), .CK(CLK), .Q(n58262), .QN(n63187) );
  DFF_X1 \REGISTERS_reg[20][38]  ( .D(n6181), .CK(CLK), .Q(n58261), .QN(n63188) );
  DFF_X1 \REGISTERS_reg[20][37]  ( .D(n6180), .CK(CLK), .Q(n58260), .QN(n63189) );
  DFF_X1 \REGISTERS_reg[20][36]  ( .D(n6179), .CK(CLK), .Q(n58259), .QN(n63190) );
  DFF_X1 \REGISTERS_reg[20][35]  ( .D(n6178), .CK(CLK), .Q(n58258), .QN(n63191) );
  DFF_X1 \REGISTERS_reg[20][34]  ( .D(n6177), .CK(CLK), .Q(n58257), .QN(n63192) );
  DFF_X1 \REGISTERS_reg[20][33]  ( .D(n6176), .CK(CLK), .Q(n58256), .QN(n63193) );
  DFF_X1 \REGISTERS_reg[20][32]  ( .D(n6175), .CK(CLK), .Q(n58255), .QN(n63194) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n6174), .CK(CLK), .Q(n58254), .QN(n63195) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n6173), .CK(CLK), .Q(n58253), .QN(n63196) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n6172), .CK(CLK), .Q(n58252), .QN(n63197) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n6171), .CK(CLK), .Q(n58251), .QN(n63198) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n6170), .CK(CLK), .Q(n58250), .QN(n63199) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n6169), .CK(CLK), .Q(n58249), .QN(n63200) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n6168), .CK(CLK), .Q(n58248), .QN(n63201) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n6167), .CK(CLK), .Q(n58247), .QN(n63202) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n6166), .CK(CLK), .Q(n58246), .QN(n63203) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n6165), .CK(CLK), .Q(n58245), .QN(n63204) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n6164), .CK(CLK), .Q(n58244), .QN(n63205) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n6163), .CK(CLK), .Q(n58243), .QN(n63206) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n6162), .CK(CLK), .Q(n58242), .QN(n63207) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n6161), .CK(CLK), .Q(n58241), .QN(n63208) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n6160), .CK(CLK), .Q(n58240), .QN(n63209) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n6159), .CK(CLK), .Q(n58239), .QN(n63210) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n6158), .CK(CLK), .Q(n58238), .QN(n63211) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n6157), .CK(CLK), .Q(n58237), .QN(n63212) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n6156), .CK(CLK), .Q(n58236), .QN(n63213) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n6155), .CK(CLK), .Q(n58235), .QN(n63214) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n6154), .CK(CLK), .Q(n58294), .QN(n63215) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n6153), .CK(CLK), .Q(n58293), .QN(n63216) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n6152), .CK(CLK), .Q(n58292), .QN(n63217)
         );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n6151), .CK(CLK), .Q(n58291), .QN(n63218)
         );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n6150), .CK(CLK), .Q(n58290), .QN(n63219)
         );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n6149), .CK(CLK), .Q(n58289), .QN(n63220)
         );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n6148), .CK(CLK), .Q(n58288), .QN(n63221)
         );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n6147), .CK(CLK), .Q(n58287), .QN(n63222)
         );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n6146), .CK(CLK), .Q(n58286), .QN(n63223)
         );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n6145), .CK(CLK), .Q(n58285), .QN(n63224)
         );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n6144), .CK(CLK), .Q(n58284), .QN(n63225)
         );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n6143), .CK(CLK), .Q(n58283), .QN(n63226)
         );
  DFF_X1 \REGISTERS_reg[11][63]  ( .D(n6782), .CK(CLK), .QN(n62697) );
  DFF_X1 \REGISTERS_reg[11][62]  ( .D(n6781), .CK(CLK), .QN(n62699) );
  DFF_X1 \REGISTERS_reg[11][61]  ( .D(n6780), .CK(CLK), .QN(n62700) );
  DFF_X1 \REGISTERS_reg[11][60]  ( .D(n6779), .CK(CLK), .QN(n62701) );
  DFF_X1 \REGISTERS_reg[9][63]  ( .D(n6910), .CK(CLK), .Q(n8895), .QN(n62627)
         );
  DFF_X1 \REGISTERS_reg[9][62]  ( .D(n6909), .CK(CLK), .Q(n8896), .QN(n62629)
         );
  DFF_X1 \REGISTERS_reg[9][61]  ( .D(n6908), .CK(CLK), .Q(n8897), .QN(n62630)
         );
  DFF_X1 \REGISTERS_reg[9][60]  ( .D(n6907), .CK(CLK), .Q(n8898), .QN(n62631)
         );
  DFF_X1 \REGISTERS_reg[15][63]  ( .D(n6526), .CK(CLK), .Q(n58654), .QN(n62893) );
  DFF_X1 \REGISTERS_reg[15][62]  ( .D(n6525), .CK(CLK), .Q(n58653), .QN(n62895) );
  DFF_X1 \REGISTERS_reg[15][61]  ( .D(n6524), .CK(CLK), .Q(n58652), .QN(n62896) );
  DFF_X1 \REGISTERS_reg[15][60]  ( .D(n6523), .CK(CLK), .Q(n58651), .QN(n62897) );
  DFF_X1 \REGISTERS_reg[0][59]  ( .D(n7482), .CK(CLK), .Q(n56603), .QN(n61967)
         );
  DFF_X1 \REGISTERS_reg[0][58]  ( .D(n7481), .CK(CLK), .Q(n56627), .QN(n61969)
         );
  DFF_X1 \REGISTERS_reg[0][57]  ( .D(n7480), .CK(CLK), .Q(n56651), .QN(n61971)
         );
  DFF_X1 \REGISTERS_reg[0][56]  ( .D(n7479), .CK(CLK), .Q(n56675), .QN(n61973)
         );
  DFF_X1 \REGISTERS_reg[0][55]  ( .D(n7478), .CK(CLK), .Q(n56699), .QN(n61975)
         );
  DFF_X1 \REGISTERS_reg[0][54]  ( .D(n7477), .CK(CLK), .Q(n56723), .QN(n61977)
         );
  DFF_X1 \REGISTERS_reg[0][53]  ( .D(n7476), .CK(CLK), .Q(n56747), .QN(n61979)
         );
  DFF_X1 \REGISTERS_reg[0][52]  ( .D(n7475), .CK(CLK), .Q(n56771), .QN(n61981)
         );
  DFF_X1 \REGISTERS_reg[0][51]  ( .D(n7474), .CK(CLK), .Q(n56795), .QN(n61983)
         );
  DFF_X1 \REGISTERS_reg[0][50]  ( .D(n7473), .CK(CLK), .Q(n56819), .QN(n61985)
         );
  DFF_X1 \REGISTERS_reg[0][49]  ( .D(n7472), .CK(CLK), .Q(n56843), .QN(n61987)
         );
  DFF_X1 \REGISTERS_reg[0][48]  ( .D(n7471), .CK(CLK), .Q(n56867), .QN(n61989)
         );
  DFF_X1 \REGISTERS_reg[0][47]  ( .D(n7470), .CK(CLK), .Q(n56891), .QN(n61991)
         );
  DFF_X1 \REGISTERS_reg[0][46]  ( .D(n7469), .CK(CLK), .Q(n56915), .QN(n61993)
         );
  DFF_X1 \REGISTERS_reg[0][45]  ( .D(n7468), .CK(CLK), .Q(n56939), .QN(n61995)
         );
  DFF_X1 \REGISTERS_reg[0][44]  ( .D(n7467), .CK(CLK), .Q(n56963), .QN(n61997)
         );
  DFF_X1 \REGISTERS_reg[0][43]  ( .D(n7466), .CK(CLK), .Q(n56987), .QN(n61999)
         );
  DFF_X1 \REGISTERS_reg[0][42]  ( .D(n7465), .CK(CLK), .Q(n57011), .QN(n62001)
         );
  DFF_X1 \REGISTERS_reg[0][41]  ( .D(n7464), .CK(CLK), .Q(n57035), .QN(n62003)
         );
  DFF_X1 \REGISTERS_reg[0][40]  ( .D(n7463), .CK(CLK), .Q(n57059), .QN(n62005)
         );
  DFF_X1 \REGISTERS_reg[0][39]  ( .D(n7462), .CK(CLK), .Q(n57083), .QN(n62007)
         );
  DFF_X1 \REGISTERS_reg[0][38]  ( .D(n7461), .CK(CLK), .Q(n57107), .QN(n62009)
         );
  DFF_X1 \REGISTERS_reg[0][37]  ( .D(n7460), .CK(CLK), .Q(n57131), .QN(n62011)
         );
  DFF_X1 \REGISTERS_reg[0][36]  ( .D(n7459), .CK(CLK), .Q(n57155), .QN(n62013)
         );
  DFF_X1 \REGISTERS_reg[0][35]  ( .D(n7458), .CK(CLK), .Q(n57179), .QN(n62015)
         );
  DFF_X1 \REGISTERS_reg[0][34]  ( .D(n7457), .CK(CLK), .Q(n57203), .QN(n62017)
         );
  DFF_X1 \REGISTERS_reg[0][33]  ( .D(n7456), .CK(CLK), .Q(n57227), .QN(n62019)
         );
  DFF_X1 \REGISTERS_reg[0][32]  ( .D(n7455), .CK(CLK), .Q(n57251), .QN(n62021)
         );
  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n7454), .CK(CLK), .Q(n57275), .QN(n62023)
         );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n7453), .CK(CLK), .Q(n57299), .QN(n62025)
         );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n7452), .CK(CLK), .Q(n57323), .QN(n62027)
         );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n7451), .CK(CLK), .Q(n57347), .QN(n62029)
         );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n7450), .CK(CLK), .Q(n57371), .QN(n62031)
         );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n7449), .CK(CLK), .Q(n57395), .QN(n62033)
         );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n7448), .CK(CLK), .Q(n57419), .QN(n62035)
         );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n7447), .CK(CLK), .Q(n57443), .QN(n62037)
         );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n7446), .CK(CLK), .Q(n57467), .QN(n62039)
         );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n7445), .CK(CLK), .Q(n57491), .QN(n62041)
         );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n7444), .CK(CLK), .Q(n57515), .QN(n62043)
         );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n7443), .CK(CLK), .Q(n57539), .QN(n62045)
         );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n7442), .CK(CLK), .Q(n57563), .QN(n62047)
         );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n7441), .CK(CLK), .Q(n57587), .QN(n62049)
         );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n7440), .CK(CLK), .Q(n57611), .QN(n62051)
         );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n7439), .CK(CLK), .Q(n57635), .QN(n62053)
         );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n7438), .CK(CLK), .Q(n57659), .QN(n62055)
         );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n7437), .CK(CLK), .Q(n57683), .QN(n62057)
         );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n7436), .CK(CLK), .Q(n57707), .QN(n62059)
         );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n7435), .CK(CLK), .Q(n57731), .QN(n62061)
         );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n7434), .CK(CLK), .Q(n57755), .QN(n62063)
         );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n7433), .CK(CLK), .Q(n57779), .QN(n62065)
         );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n7432), .CK(CLK), .Q(n57803), .QN(n62067)
         );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n7431), .CK(CLK), .Q(n57827), .QN(n62069)
         );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n7430), .CK(CLK), .Q(n57851), .QN(n62071)
         );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n7429), .CK(CLK), .Q(n57875), .QN(n62073)
         );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n7428), .CK(CLK), .Q(n57899), .QN(n62075)
         );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n7427), .CK(CLK), .Q(n57923), .QN(n62077)
         );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n7426), .CK(CLK), .Q(n57947), .QN(n62079)
         );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n7425), .CK(CLK), .Q(n57971), .QN(n62081)
         );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n7424), .CK(CLK), .Q(n57995), .QN(n62083)
         );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n7423), .CK(CLK), .Q(n58028), .QN(n62085)
         );
  DFF_X1 \REGISTERS_reg[7][59]  ( .D(n7034), .CK(CLK), .Q(n58110), .QN(n62499)
         );
  DFF_X1 \REGISTERS_reg[7][58]  ( .D(n7033), .CK(CLK), .Q(n58109), .QN(n62500)
         );
  DFF_X1 \REGISTERS_reg[7][57]  ( .D(n7032), .CK(CLK), .Q(n58108), .QN(n62501)
         );
  DFF_X1 \REGISTERS_reg[7][56]  ( .D(n7031), .CK(CLK), .Q(n58107), .QN(n62502)
         );
  DFF_X1 \REGISTERS_reg[7][55]  ( .D(n7030), .CK(CLK), .Q(n58106), .QN(n62503)
         );
  DFF_X1 \REGISTERS_reg[7][54]  ( .D(n7029), .CK(CLK), .Q(n58105), .QN(n62504)
         );
  DFF_X1 \REGISTERS_reg[7][53]  ( .D(n7028), .CK(CLK), .Q(n58104), .QN(n62505)
         );
  DFF_X1 \REGISTERS_reg[7][52]  ( .D(n7027), .CK(CLK), .Q(n58103), .QN(n62506)
         );
  DFF_X1 \REGISTERS_reg[7][51]  ( .D(n7026), .CK(CLK), .Q(n58102), .QN(n62507)
         );
  DFF_X1 \REGISTERS_reg[7][50]  ( .D(n7025), .CK(CLK), .Q(n58101), .QN(n62508)
         );
  DFF_X1 \REGISTERS_reg[7][49]  ( .D(n7024), .CK(CLK), .Q(n58100), .QN(n62509)
         );
  DFF_X1 \REGISTERS_reg[7][48]  ( .D(n7023), .CK(CLK), .Q(n58099), .QN(n62510)
         );
  DFF_X1 \REGISTERS_reg[7][47]  ( .D(n7022), .CK(CLK), .Q(n58098), .QN(n62511)
         );
  DFF_X1 \REGISTERS_reg[7][46]  ( .D(n7021), .CK(CLK), .Q(n58097), .QN(n62512)
         );
  DFF_X1 \REGISTERS_reg[7][45]  ( .D(n7020), .CK(CLK), .Q(n58096), .QN(n62513)
         );
  DFF_X1 \REGISTERS_reg[7][44]  ( .D(n7019), .CK(CLK), .Q(n58095), .QN(n62514)
         );
  DFF_X1 \REGISTERS_reg[7][43]  ( .D(n7018), .CK(CLK), .Q(n58094), .QN(n62515)
         );
  DFF_X1 \REGISTERS_reg[7][42]  ( .D(n7017), .CK(CLK), .Q(n58093), .QN(n62516)
         );
  DFF_X1 \REGISTERS_reg[7][41]  ( .D(n7016), .CK(CLK), .Q(n58092), .QN(n62517)
         );
  DFF_X1 \REGISTERS_reg[7][40]  ( .D(n7015), .CK(CLK), .Q(n58091), .QN(n62518)
         );
  DFF_X1 \REGISTERS_reg[7][39]  ( .D(n7014), .CK(CLK), .Q(n58090), .QN(n62519)
         );
  DFF_X1 \REGISTERS_reg[7][38]  ( .D(n7013), .CK(CLK), .Q(n58089), .QN(n62520)
         );
  DFF_X1 \REGISTERS_reg[7][37]  ( .D(n7012), .CK(CLK), .Q(n58088), .QN(n62521)
         );
  DFF_X1 \REGISTERS_reg[7][36]  ( .D(n7011), .CK(CLK), .Q(n58087), .QN(n62522)
         );
  DFF_X1 \REGISTERS_reg[7][35]  ( .D(n7010), .CK(CLK), .Q(n58086), .QN(n62523)
         );
  DFF_X1 \REGISTERS_reg[7][34]  ( .D(n7009), .CK(CLK), .Q(n58085), .QN(n62524)
         );
  DFF_X1 \REGISTERS_reg[7][33]  ( .D(n7008), .CK(CLK), .Q(n58084), .QN(n62525)
         );
  DFF_X1 \REGISTERS_reg[7][32]  ( .D(n7007), .CK(CLK), .Q(n58083), .QN(n62526)
         );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n7006), .CK(CLK), .Q(n58082), .QN(n62527)
         );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n7005), .CK(CLK), .Q(n58081), .QN(n62528)
         );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n7004), .CK(CLK), .Q(n58080), .QN(n62529)
         );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n7003), .CK(CLK), .Q(n58079), .QN(n62530)
         );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n7002), .CK(CLK), .Q(n58078), .QN(n62531)
         );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n7001), .CK(CLK), .Q(n58077), .QN(n62532)
         );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n7000), .CK(CLK), .Q(n58076), .QN(n62533)
         );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n6999), .CK(CLK), .Q(n58075), .QN(n62534)
         );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n6998), .CK(CLK), .Q(n58074), .QN(n62535)
         );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n6997), .CK(CLK), .Q(n58073), .QN(n62536)
         );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n6996), .CK(CLK), .Q(n58072), .QN(n62537)
         );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n6995), .CK(CLK), .Q(n58071), .QN(n62538)
         );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n6994), .CK(CLK), .Q(n58070), .QN(n62539)
         );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n6993), .CK(CLK), .Q(n58069), .QN(n62540)
         );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n6992), .CK(CLK), .Q(n58068), .QN(n62541)
         );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n6991), .CK(CLK), .Q(n58067), .QN(n62542)
         );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n6990), .CK(CLK), .Q(n58066), .QN(n62543)
         );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n6989), .CK(CLK), .Q(n58065), .QN(n62544)
         );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n6988), .CK(CLK), .Q(n58064), .QN(n62545)
         );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n6987), .CK(CLK), .Q(n58063), .QN(n62546)
         );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n6986), .CK(CLK), .Q(n58062), .QN(n62547)
         );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n6985), .CK(CLK), .Q(n58061), .QN(n62548)
         );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n6984), .CK(CLK), .Q(n58060), .QN(n62549)
         );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n6983), .CK(CLK), .Q(n58059), .QN(n62550)
         );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n6982), .CK(CLK), .Q(n58058), .QN(n62551)
         );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n6981), .CK(CLK), .Q(n58057), .QN(n62552)
         );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n6980), .CK(CLK), .Q(n58056), .QN(n62553)
         );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n6979), .CK(CLK), .Q(n58055), .QN(n62554)
         );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n6978), .CK(CLK), .Q(n58054), .QN(n62555)
         );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n6977), .CK(CLK), .Q(n58053), .QN(n62556)
         );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n6976), .CK(CLK), .Q(n58052), .QN(n62557)
         );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n6975), .CK(CLK), .Q(n58051), .QN(n62558)
         );
  DFF_X1 \REGISTERS_reg[5][59]  ( .D(n7162), .CK(CLK), .Q(n58842), .QN(n62363)
         );
  DFF_X1 \REGISTERS_reg[5][58]  ( .D(n7161), .CK(CLK), .Q(n58841), .QN(n62364)
         );
  DFF_X1 \REGISTERS_reg[5][57]  ( .D(n7160), .CK(CLK), .Q(n58840), .QN(n62365)
         );
  DFF_X1 \REGISTERS_reg[5][56]  ( .D(n7159), .CK(CLK), .Q(n58839), .QN(n62366)
         );
  DFF_X1 \REGISTERS_reg[5][55]  ( .D(n7158), .CK(CLK), .Q(n58838), .QN(n62367)
         );
  DFF_X1 \REGISTERS_reg[5][54]  ( .D(n7157), .CK(CLK), .Q(n58837), .QN(n62368)
         );
  DFF_X1 \REGISTERS_reg[5][53]  ( .D(n7156), .CK(CLK), .Q(n58836), .QN(n62369)
         );
  DFF_X1 \REGISTERS_reg[5][52]  ( .D(n7155), .CK(CLK), .Q(n58835), .QN(n62370)
         );
  DFF_X1 \REGISTERS_reg[5][51]  ( .D(n7154), .CK(CLK), .Q(n58834), .QN(n62371)
         );
  DFF_X1 \REGISTERS_reg[5][50]  ( .D(n7153), .CK(CLK), .Q(n58833), .QN(n62372)
         );
  DFF_X1 \REGISTERS_reg[5][49]  ( .D(n7152), .CK(CLK), .Q(n58832), .QN(n62373)
         );
  DFF_X1 \REGISTERS_reg[5][48]  ( .D(n7151), .CK(CLK), .Q(n58831), .QN(n62374)
         );
  DFF_X1 \REGISTERS_reg[5][47]  ( .D(n7150), .CK(CLK), .Q(n58830), .QN(n62375)
         );
  DFF_X1 \REGISTERS_reg[5][46]  ( .D(n7149), .CK(CLK), .Q(n58829), .QN(n62376)
         );
  DFF_X1 \REGISTERS_reg[5][45]  ( .D(n7148), .CK(CLK), .Q(n58828), .QN(n62377)
         );
  DFF_X1 \REGISTERS_reg[5][44]  ( .D(n7147), .CK(CLK), .Q(n58827), .QN(n62378)
         );
  DFF_X1 \REGISTERS_reg[5][43]  ( .D(n7146), .CK(CLK), .Q(n58826), .QN(n62379)
         );
  DFF_X1 \REGISTERS_reg[5][42]  ( .D(n7145), .CK(CLK), .Q(n58825), .QN(n62380)
         );
  DFF_X1 \REGISTERS_reg[5][41]  ( .D(n7144), .CK(CLK), .Q(n58824), .QN(n62381)
         );
  DFF_X1 \REGISTERS_reg[5][40]  ( .D(n7143), .CK(CLK), .Q(n58823), .QN(n62382)
         );
  DFF_X1 \REGISTERS_reg[5][39]  ( .D(n7142), .CK(CLK), .Q(n58822), .QN(n62383)
         );
  DFF_X1 \REGISTERS_reg[5][38]  ( .D(n7141), .CK(CLK), .Q(n58821), .QN(n62384)
         );
  DFF_X1 \REGISTERS_reg[5][37]  ( .D(n7140), .CK(CLK), .Q(n58820), .QN(n62385)
         );
  DFF_X1 \REGISTERS_reg[5][36]  ( .D(n7139), .CK(CLK), .Q(n58819), .QN(n62386)
         );
  DFF_X1 \REGISTERS_reg[5][35]  ( .D(n7138), .CK(CLK), .Q(n58818), .QN(n62387)
         );
  DFF_X1 \REGISTERS_reg[5][34]  ( .D(n7137), .CK(CLK), .Q(n58817), .QN(n62388)
         );
  DFF_X1 \REGISTERS_reg[5][33]  ( .D(n7136), .CK(CLK), .Q(n58816), .QN(n62389)
         );
  DFF_X1 \REGISTERS_reg[5][32]  ( .D(n7135), .CK(CLK), .Q(n58815), .QN(n62390)
         );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n7134), .CK(CLK), .Q(n58814), .QN(n62391)
         );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n7133), .CK(CLK), .Q(n58813), .QN(n62392)
         );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n7132), .CK(CLK), .Q(n58812), .QN(n62393)
         );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n7131), .CK(CLK), .Q(n58811), .QN(n62394)
         );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n7130), .CK(CLK), .Q(n58810), .QN(n62395)
         );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n7129), .CK(CLK), .Q(n58809), .QN(n62396)
         );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n7128), .CK(CLK), .Q(n58808), .QN(n62397)
         );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n7127), .CK(CLK), .Q(n58807), .QN(n62398)
         );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n7126), .CK(CLK), .Q(n58806), .QN(n62399)
         );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n7125), .CK(CLK), .Q(n58805), .QN(n62400)
         );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n7124), .CK(CLK), .Q(n58804), .QN(n62401)
         );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n7123), .CK(CLK), .Q(n58803), .QN(n62402)
         );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n7122), .CK(CLK), .Q(n58802), .QN(n62403)
         );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n7121), .CK(CLK), .Q(n58801), .QN(n62404)
         );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n7120), .CK(CLK), .Q(n58800), .QN(n62405)
         );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n7119), .CK(CLK), .Q(n58799), .QN(n62406)
         );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n7118), .CK(CLK), .Q(n56020), .QN(n62407)
         );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n7117), .CK(CLK), .Q(n56047), .QN(n62408)
         );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n7116), .CK(CLK), .Q(n56074), .QN(n62409)
         );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n7115), .CK(CLK), .Q(n56101), .QN(n62410)
         );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n7114), .CK(CLK), .Q(n58798), .QN(n62411)
         );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n7113), .CK(CLK), .Q(n58797), .QN(n62412)
         );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n7112), .CK(CLK), .Q(n58796), .QN(n62413)
         );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n7111), .CK(CLK), .Q(n58795), .QN(n62414)
         );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n7110), .CK(CLK), .Q(n58794), .QN(n62415)
         );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n7109), .CK(CLK), .Q(n58793), .QN(n62416)
         );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n7108), .CK(CLK), .Q(n58792), .QN(n62417)
         );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n7107), .CK(CLK), .Q(n58791), .QN(n62418)
         );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n7106), .CK(CLK), .Q(n58790), .QN(n62419)
         );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n7105), .CK(CLK), .Q(n58789), .QN(n62420)
         );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n7104), .CK(CLK), .Q(n58788), .QN(n62421)
         );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n7103), .CK(CLK), .Q(n58787), .QN(n62422)
         );
  DFF_X1 \REGISTERS_reg[3][59]  ( .D(n7290), .CK(CLK), .QN(n62230) );
  DFF_X1 \REGISTERS_reg[3][58]  ( .D(n7289), .CK(CLK), .QN(n62231) );
  DFF_X1 \REGISTERS_reg[3][57]  ( .D(n7288), .CK(CLK), .QN(n62232) );
  DFF_X1 \REGISTERS_reg[3][56]  ( .D(n7287), .CK(CLK), .QN(n62233) );
  DFF_X1 \REGISTERS_reg[3][55]  ( .D(n7286), .CK(CLK), .QN(n62234) );
  DFF_X1 \REGISTERS_reg[3][54]  ( .D(n7285), .CK(CLK), .QN(n62235) );
  DFF_X1 \REGISTERS_reg[3][53]  ( .D(n7284), .CK(CLK), .QN(n62236) );
  DFF_X1 \REGISTERS_reg[3][52]  ( .D(n7283), .CK(CLK), .QN(n62237) );
  DFF_X1 \REGISTERS_reg[3][51]  ( .D(n7282), .CK(CLK), .QN(n62238) );
  DFF_X1 \REGISTERS_reg[3][50]  ( .D(n7281), .CK(CLK), .QN(n62239) );
  DFF_X1 \REGISTERS_reg[3][49]  ( .D(n7280), .CK(CLK), .QN(n62240) );
  DFF_X1 \REGISTERS_reg[3][48]  ( .D(n7279), .CK(CLK), .QN(n62241) );
  DFF_X1 \REGISTERS_reg[3][47]  ( .D(n7278), .CK(CLK), .QN(n62242) );
  DFF_X1 \REGISTERS_reg[3][46]  ( .D(n7277), .CK(CLK), .QN(n62243) );
  DFF_X1 \REGISTERS_reg[3][45]  ( .D(n7276), .CK(CLK), .QN(n62244) );
  DFF_X1 \REGISTERS_reg[3][44]  ( .D(n7275), .CK(CLK), .QN(n62245) );
  DFF_X1 \REGISTERS_reg[3][43]  ( .D(n7274), .CK(CLK), .QN(n62246) );
  DFF_X1 \REGISTERS_reg[3][42]  ( .D(n7273), .CK(CLK), .QN(n62247) );
  DFF_X1 \REGISTERS_reg[3][41]  ( .D(n7272), .CK(CLK), .QN(n62248) );
  DFF_X1 \REGISTERS_reg[3][40]  ( .D(n7271), .CK(CLK), .QN(n62249) );
  DFF_X1 \REGISTERS_reg[3][39]  ( .D(n7270), .CK(CLK), .QN(n62250) );
  DFF_X1 \REGISTERS_reg[3][38]  ( .D(n7269), .CK(CLK), .QN(n62251) );
  DFF_X1 \REGISTERS_reg[3][37]  ( .D(n7268), .CK(CLK), .QN(n62252) );
  DFF_X1 \REGISTERS_reg[3][36]  ( .D(n7267), .CK(CLK), .QN(n62253) );
  DFF_X1 \REGISTERS_reg[3][35]  ( .D(n7266), .CK(CLK), .QN(n62254) );
  DFF_X1 \REGISTERS_reg[3][34]  ( .D(n7265), .CK(CLK), .QN(n62255) );
  DFF_X1 \REGISTERS_reg[3][33]  ( .D(n7264), .CK(CLK), .QN(n62256) );
  DFF_X1 \REGISTERS_reg[3][32]  ( .D(n7263), .CK(CLK), .QN(n62257) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n7262), .CK(CLK), .QN(n62258) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n7261), .CK(CLK), .QN(n62259) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n7260), .CK(CLK), .QN(n62260) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n7259), .CK(CLK), .QN(n62261) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n7258), .CK(CLK), .QN(n62262) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n7257), .CK(CLK), .QN(n62263) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n7256), .CK(CLK), .QN(n62264) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n7255), .CK(CLK), .QN(n62265) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n7254), .CK(CLK), .QN(n62266) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n7253), .CK(CLK), .QN(n62267) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n7252), .CK(CLK), .QN(n62268) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n7251), .CK(CLK), .QN(n62269) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n7250), .CK(CLK), .QN(n62270) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n7249), .CK(CLK), .QN(n62271) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n7248), .CK(CLK), .QN(n62272) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n7247), .CK(CLK), .QN(n62273) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n7246), .CK(CLK), .QN(n62274) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n7245), .CK(CLK), .QN(n62275) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n7244), .CK(CLK), .QN(n62276) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n7243), .CK(CLK), .QN(n62277) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n7242), .CK(CLK), .QN(n62278) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n7241), .CK(CLK), .QN(n62279) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n7240), .CK(CLK), .QN(n62280) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n7239), .CK(CLK), .QN(n62281) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n7238), .CK(CLK), .QN(n62282) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n7237), .CK(CLK), .QN(n62283) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n7236), .CK(CLK), .QN(n62284) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n7235), .CK(CLK), .QN(n62285) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n7234), .CK(CLK), .QN(n62286) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n7233), .CK(CLK), .QN(n62287) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n7232), .CK(CLK), .QN(n62288) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n7231), .CK(CLK), .QN(n62289) );
  DFF_X1 \REGISTERS_reg[2][59]  ( .D(n7354), .CK(CLK), .QN(n62163) );
  DFF_X1 \REGISTERS_reg[2][58]  ( .D(n7353), .CK(CLK), .QN(n62164) );
  DFF_X1 \REGISTERS_reg[2][57]  ( .D(n7352), .CK(CLK), .QN(n62165) );
  DFF_X1 \REGISTERS_reg[2][56]  ( .D(n7351), .CK(CLK), .QN(n62166) );
  DFF_X1 \REGISTERS_reg[2][55]  ( .D(n7350), .CK(CLK), .QN(n62167) );
  DFF_X1 \REGISTERS_reg[2][54]  ( .D(n7349), .CK(CLK), .QN(n62168) );
  DFF_X1 \REGISTERS_reg[2][53]  ( .D(n7348), .CK(CLK), .QN(n62169) );
  DFF_X1 \REGISTERS_reg[2][52]  ( .D(n7347), .CK(CLK), .QN(n62170) );
  DFF_X1 \REGISTERS_reg[2][51]  ( .D(n7346), .CK(CLK), .QN(n62171) );
  DFF_X1 \REGISTERS_reg[2][50]  ( .D(n7345), .CK(CLK), .QN(n62172) );
  DFF_X1 \REGISTERS_reg[2][49]  ( .D(n7344), .CK(CLK), .QN(n62173) );
  DFF_X1 \REGISTERS_reg[2][48]  ( .D(n7343), .CK(CLK), .QN(n62174) );
  DFF_X1 \REGISTERS_reg[2][47]  ( .D(n7342), .CK(CLK), .QN(n62175) );
  DFF_X1 \REGISTERS_reg[2][46]  ( .D(n7341), .CK(CLK), .QN(n62176) );
  DFF_X1 \REGISTERS_reg[2][45]  ( .D(n7340), .CK(CLK), .QN(n62177) );
  DFF_X1 \REGISTERS_reg[2][44]  ( .D(n7339), .CK(CLK), .QN(n62178) );
  DFF_X1 \REGISTERS_reg[2][43]  ( .D(n7338), .CK(CLK), .QN(n62179) );
  DFF_X1 \REGISTERS_reg[2][42]  ( .D(n7337), .CK(CLK), .QN(n62180) );
  DFF_X1 \REGISTERS_reg[2][41]  ( .D(n7336), .CK(CLK), .QN(n62181) );
  DFF_X1 \REGISTERS_reg[2][40]  ( .D(n7335), .CK(CLK), .QN(n62182) );
  DFF_X1 \REGISTERS_reg[2][39]  ( .D(n7334), .CK(CLK), .QN(n62183) );
  DFF_X1 \REGISTERS_reg[2][38]  ( .D(n7333), .CK(CLK), .QN(n62184) );
  DFF_X1 \REGISTERS_reg[2][37]  ( .D(n7332), .CK(CLK), .QN(n62185) );
  DFF_X1 \REGISTERS_reg[2][36]  ( .D(n7331), .CK(CLK), .QN(n62186) );
  DFF_X1 \REGISTERS_reg[2][35]  ( .D(n7330), .CK(CLK), .QN(n62187) );
  DFF_X1 \REGISTERS_reg[2][34]  ( .D(n7329), .CK(CLK), .QN(n62188) );
  DFF_X1 \REGISTERS_reg[2][33]  ( .D(n7328), .CK(CLK), .QN(n62189) );
  DFF_X1 \REGISTERS_reg[2][32]  ( .D(n7327), .CK(CLK), .QN(n62190) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n7326), .CK(CLK), .QN(n62191) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n7325), .CK(CLK), .QN(n62192) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n7324), .CK(CLK), .QN(n62193) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n7323), .CK(CLK), .QN(n62194) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n7322), .CK(CLK), .QN(n62195) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n7321), .CK(CLK), .QN(n62196) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n7320), .CK(CLK), .QN(n62197) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n7319), .CK(CLK), .QN(n62198) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n7318), .CK(CLK), .QN(n62199) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n7317), .CK(CLK), .QN(n62200) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n7316), .CK(CLK), .QN(n62201) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n7315), .CK(CLK), .QN(n62202) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n7314), .CK(CLK), .QN(n62203) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n7313), .CK(CLK), .QN(n62204) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n7312), .CK(CLK), .QN(n62205) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n7311), .CK(CLK), .QN(n62206) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n7310), .CK(CLK), .QN(n62207) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n7309), .CK(CLK), .QN(n62208) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n7308), .CK(CLK), .QN(n62209) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n7307), .CK(CLK), .QN(n62210) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n7306), .CK(CLK), .QN(n62211) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n7305), .CK(CLK), .QN(n62212) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n7304), .CK(CLK), .QN(n62213) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n7303), .CK(CLK), .QN(n62214) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n7302), .CK(CLK), .QN(n62215) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n7301), .CK(CLK), .QN(n62216) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n7300), .CK(CLK), .QN(n62217) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n7299), .CK(CLK), .QN(n62218) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n7298), .CK(CLK), .QN(n62219) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n7297), .CK(CLK), .QN(n62220) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n7296), .CK(CLK), .QN(n62221) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n7295), .CK(CLK), .QN(n62222) );
  DFF_X1 \REGISTERS_reg[6][59]  ( .D(n7098), .CK(CLK), .QN(n62429) );
  DFF_X1 \REGISTERS_reg[6][58]  ( .D(n7097), .CK(CLK), .QN(n62430) );
  DFF_X1 \REGISTERS_reg[6][57]  ( .D(n7096), .CK(CLK), .QN(n62431) );
  DFF_X1 \REGISTERS_reg[6][56]  ( .D(n7095), .CK(CLK), .QN(n62432) );
  DFF_X1 \REGISTERS_reg[6][55]  ( .D(n7094), .CK(CLK), .QN(n62433) );
  DFF_X1 \REGISTERS_reg[6][54]  ( .D(n7093), .CK(CLK), .QN(n62434) );
  DFF_X1 \REGISTERS_reg[6][53]  ( .D(n7092), .CK(CLK), .QN(n62435) );
  DFF_X1 \REGISTERS_reg[6][52]  ( .D(n7091), .CK(CLK), .QN(n62436) );
  DFF_X1 \REGISTERS_reg[6][51]  ( .D(n7090), .CK(CLK), .QN(n62437) );
  DFF_X1 \REGISTERS_reg[6][50]  ( .D(n7089), .CK(CLK), .QN(n62438) );
  DFF_X1 \REGISTERS_reg[6][49]  ( .D(n7088), .CK(CLK), .QN(n62439) );
  DFF_X1 \REGISTERS_reg[6][48]  ( .D(n7087), .CK(CLK), .QN(n62440) );
  DFF_X1 \REGISTERS_reg[6][47]  ( .D(n7086), .CK(CLK), .QN(n62441) );
  DFF_X1 \REGISTERS_reg[6][46]  ( .D(n7085), .CK(CLK), .QN(n62442) );
  DFF_X1 \REGISTERS_reg[6][45]  ( .D(n7084), .CK(CLK), .QN(n62443) );
  DFF_X1 \REGISTERS_reg[6][44]  ( .D(n7083), .CK(CLK), .QN(n62444) );
  DFF_X1 \REGISTERS_reg[6][43]  ( .D(n7082), .CK(CLK), .QN(n62445) );
  DFF_X1 \REGISTERS_reg[6][42]  ( .D(n7081), .CK(CLK), .QN(n62446) );
  DFF_X1 \REGISTERS_reg[6][41]  ( .D(n7080), .CK(CLK), .QN(n62447) );
  DFF_X1 \REGISTERS_reg[6][40]  ( .D(n7079), .CK(CLK), .QN(n62448) );
  DFF_X1 \REGISTERS_reg[6][39]  ( .D(n7078), .CK(CLK), .QN(n62449) );
  DFF_X1 \REGISTERS_reg[6][38]  ( .D(n7077), .CK(CLK), .QN(n62450) );
  DFF_X1 \REGISTERS_reg[6][37]  ( .D(n7076), .CK(CLK), .QN(n62451) );
  DFF_X1 \REGISTERS_reg[6][36]  ( .D(n7075), .CK(CLK), .QN(n62452) );
  DFF_X1 \REGISTERS_reg[6][35]  ( .D(n7074), .CK(CLK), .QN(n62453) );
  DFF_X1 \REGISTERS_reg[6][34]  ( .D(n7073), .CK(CLK), .QN(n62454) );
  DFF_X1 \REGISTERS_reg[6][33]  ( .D(n7072), .CK(CLK), .QN(n62455) );
  DFF_X1 \REGISTERS_reg[6][32]  ( .D(n7071), .CK(CLK), .QN(n62456) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n7070), .CK(CLK), .QN(n62457) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n7069), .CK(CLK), .QN(n62458) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n7068), .CK(CLK), .QN(n62459) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n7067), .CK(CLK), .QN(n62460) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n7066), .CK(CLK), .QN(n62461) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n7065), .CK(CLK), .QN(n62462) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n7064), .CK(CLK), .QN(n62463) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n7063), .CK(CLK), .QN(n62464) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n7062), .CK(CLK), .QN(n62465) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n7061), .CK(CLK), .QN(n62466) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n7060), .CK(CLK), .QN(n62467) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n7059), .CK(CLK), .QN(n62468) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n7058), .CK(CLK), .QN(n62469) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n7057), .CK(CLK), .QN(n62470) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n7056), .CK(CLK), .QN(n62471) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n7055), .CK(CLK), .QN(n62472) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n7054), .CK(CLK), .QN(n62473) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n7053), .CK(CLK), .QN(n62474) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n7052), .CK(CLK), .QN(n62475) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n7051), .CK(CLK), .QN(n62476) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n7050), .CK(CLK), .QN(n62477) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n7049), .CK(CLK), .QN(n62478) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n7048), .CK(CLK), .QN(n62479) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n7047), .CK(CLK), .QN(n62480) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n7046), .CK(CLK), .QN(n62481) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n7045), .CK(CLK), .QN(n62482) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n7044), .CK(CLK), .QN(n62483) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n7043), .CK(CLK), .QN(n62484) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n7042), .CK(CLK), .QN(n62485) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n7041), .CK(CLK), .QN(n62486) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n7040), .CK(CLK), .QN(n62487) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n7039), .CK(CLK), .QN(n62488) );
  DFF_X1 \REGISTERS_reg[4][59]  ( .D(n7226), .CK(CLK), .Q(n59088), .QN(n62296)
         );
  DFF_X1 \REGISTERS_reg[4][58]  ( .D(n7225), .CK(CLK), .Q(n59087), .QN(n62297)
         );
  DFF_X1 \REGISTERS_reg[4][57]  ( .D(n7224), .CK(CLK), .Q(n59086), .QN(n62298)
         );
  DFF_X1 \REGISTERS_reg[4][56]  ( .D(n7223), .CK(CLK), .Q(n59085), .QN(n62299)
         );
  DFF_X1 \REGISTERS_reg[4][55]  ( .D(n7222), .CK(CLK), .Q(n59084), .QN(n62300)
         );
  DFF_X1 \REGISTERS_reg[4][54]  ( .D(n7221), .CK(CLK), .Q(n59083), .QN(n62301)
         );
  DFF_X1 \REGISTERS_reg[4][53]  ( .D(n7220), .CK(CLK), .Q(n59082), .QN(n62302)
         );
  DFF_X1 \REGISTERS_reg[4][52]  ( .D(n7219), .CK(CLK), .Q(n59081), .QN(n62303)
         );
  DFF_X1 \REGISTERS_reg[4][51]  ( .D(n7218), .CK(CLK), .Q(n59080), .QN(n62304)
         );
  DFF_X1 \REGISTERS_reg[4][50]  ( .D(n7217), .CK(CLK), .Q(n59079), .QN(n62305)
         );
  DFF_X1 \REGISTERS_reg[4][49]  ( .D(n7216), .CK(CLK), .Q(n59078), .QN(n62306)
         );
  DFF_X1 \REGISTERS_reg[4][48]  ( .D(n7215), .CK(CLK), .Q(n59077), .QN(n62307)
         );
  DFF_X1 \REGISTERS_reg[4][47]  ( .D(n7214), .CK(CLK), .Q(n59076), .QN(n62308)
         );
  DFF_X1 \REGISTERS_reg[4][46]  ( .D(n7213), .CK(CLK), .Q(n59075), .QN(n62309)
         );
  DFF_X1 \REGISTERS_reg[4][45]  ( .D(n7212), .CK(CLK), .Q(n59074), .QN(n62310)
         );
  DFF_X1 \REGISTERS_reg[4][44]  ( .D(n7211), .CK(CLK), .Q(n59073), .QN(n62311)
         );
  DFF_X1 \REGISTERS_reg[4][43]  ( .D(n7210), .CK(CLK), .Q(n59072), .QN(n62312)
         );
  DFF_X1 \REGISTERS_reg[4][42]  ( .D(n7209), .CK(CLK), .Q(n59071), .QN(n62313)
         );
  DFF_X1 \REGISTERS_reg[4][41]  ( .D(n7208), .CK(CLK), .Q(n59070), .QN(n62314)
         );
  DFF_X1 \REGISTERS_reg[4][40]  ( .D(n7207), .CK(CLK), .Q(n59069), .QN(n62315)
         );
  DFF_X1 \REGISTERS_reg[4][39]  ( .D(n7206), .CK(CLK), .Q(n59068), .QN(n62316)
         );
  DFF_X1 \REGISTERS_reg[4][38]  ( .D(n7205), .CK(CLK), .Q(n59067), .QN(n62317)
         );
  DFF_X1 \REGISTERS_reg[4][37]  ( .D(n7204), .CK(CLK), .Q(n59066), .QN(n62318)
         );
  DFF_X1 \REGISTERS_reg[4][36]  ( .D(n7203), .CK(CLK), .Q(n59065), .QN(n62319)
         );
  DFF_X1 \REGISTERS_reg[4][35]  ( .D(n7202), .CK(CLK), .Q(n59064), .QN(n62320)
         );
  DFF_X1 \REGISTERS_reg[4][34]  ( .D(n7201), .CK(CLK), .Q(n59063), .QN(n62321)
         );
  DFF_X1 \REGISTERS_reg[4][33]  ( .D(n7200), .CK(CLK), .Q(n59062), .QN(n62322)
         );
  DFF_X1 \REGISTERS_reg[4][32]  ( .D(n7199), .CK(CLK), .Q(n59061), .QN(n62323)
         );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n7198), .CK(CLK), .Q(n59060), .QN(n62324)
         );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n7197), .CK(CLK), .Q(n59059), .QN(n62325)
         );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n7196), .CK(CLK), .Q(n59058), .QN(n62326)
         );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n7195), .CK(CLK), .Q(n59057), .QN(n62327)
         );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n7194), .CK(CLK), .Q(n59056), .QN(n62328)
         );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n7193), .CK(CLK), .Q(n59055), .QN(n62329)
         );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n7192), .CK(CLK), .Q(n59054), .QN(n62330)
         );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n7191), .CK(CLK), .Q(n59053), .QN(n62331)
         );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n7190), .CK(CLK), .Q(n59052), .QN(n62332)
         );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n7189), .CK(CLK), .Q(n59051), .QN(n62333)
         );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n7188), .CK(CLK), .Q(n59050), .QN(n62334)
         );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n7187), .CK(CLK), .Q(n59049), .QN(n62335)
         );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n7186), .CK(CLK), .Q(n59048), .QN(n62336)
         );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n7185), .CK(CLK), .Q(n59047), .QN(n62337)
         );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n7184), .CK(CLK), .Q(n59046), .QN(n62338)
         );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n7183), .CK(CLK), .Q(n59045), .QN(n62339)
         );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n7182), .CK(CLK), .Q(n59044), .QN(n62340)
         );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n7181), .CK(CLK), .Q(n59043), .QN(n62341)
         );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n7180), .CK(CLK), .Q(n59042), .QN(n62342)
         );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n7179), .CK(CLK), .Q(n59041), .QN(n62343)
         );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n7178), .CK(CLK), .Q(n59040), .QN(n62344)
         );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n7177), .CK(CLK), .Q(n59039), .QN(n62345)
         );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n7176), .CK(CLK), .Q(n59038), .QN(n62346)
         );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n7175), .CK(CLK), .Q(n59037), .QN(n62347)
         );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n7174), .CK(CLK), .Q(n59036), .QN(n62348)
         );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n7173), .CK(CLK), .Q(n59035), .QN(n62349)
         );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n7172), .CK(CLK), .Q(n59034), .QN(n62350)
         );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n7171), .CK(CLK), .Q(n59033), .QN(n62351)
         );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n7170), .CK(CLK), .Q(n59032), .QN(n62352)
         );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n7169), .CK(CLK), .Q(n59031), .QN(n62353)
         );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n7168), .CK(CLK), .Q(n59030), .QN(n62354)
         );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n7167), .CK(CLK), .Q(n59029), .QN(n62355)
         );
  DFF_X1 \REGISTERS_reg[1][59]  ( .D(n7418), .CK(CLK), .QN(n62096) );
  DFF_X1 \REGISTERS_reg[1][58]  ( .D(n7417), .CK(CLK), .QN(n62097) );
  DFF_X1 \REGISTERS_reg[1][57]  ( .D(n7416), .CK(CLK), .QN(n62098) );
  DFF_X1 \REGISTERS_reg[1][56]  ( .D(n7415), .CK(CLK), .QN(n62099) );
  DFF_X1 \REGISTERS_reg[1][55]  ( .D(n7414), .CK(CLK), .QN(n62100) );
  DFF_X1 \REGISTERS_reg[1][54]  ( .D(n7413), .CK(CLK), .QN(n62101) );
  DFF_X1 \REGISTERS_reg[1][53]  ( .D(n7412), .CK(CLK), .QN(n62102) );
  DFF_X1 \REGISTERS_reg[1][52]  ( .D(n7411), .CK(CLK), .QN(n62103) );
  DFF_X1 \REGISTERS_reg[1][51]  ( .D(n7410), .CK(CLK), .QN(n62104) );
  DFF_X1 \REGISTERS_reg[1][50]  ( .D(n7409), .CK(CLK), .QN(n62105) );
  DFF_X1 \REGISTERS_reg[1][49]  ( .D(n7408), .CK(CLK), .QN(n62106) );
  DFF_X1 \REGISTERS_reg[1][48]  ( .D(n7407), .CK(CLK), .QN(n62107) );
  DFF_X1 \REGISTERS_reg[1][47]  ( .D(n7406), .CK(CLK), .QN(n62108) );
  DFF_X1 \REGISTERS_reg[1][46]  ( .D(n7405), .CK(CLK), .QN(n62109) );
  DFF_X1 \REGISTERS_reg[1][45]  ( .D(n7404), .CK(CLK), .QN(n62110) );
  DFF_X1 \REGISTERS_reg[1][44]  ( .D(n7403), .CK(CLK), .QN(n62111) );
  DFF_X1 \REGISTERS_reg[1][43]  ( .D(n7402), .CK(CLK), .QN(n62112) );
  DFF_X1 \REGISTERS_reg[1][42]  ( .D(n7401), .CK(CLK), .QN(n62113) );
  DFF_X1 \REGISTERS_reg[1][41]  ( .D(n7400), .CK(CLK), .QN(n62114) );
  DFF_X1 \REGISTERS_reg[1][40]  ( .D(n7399), .CK(CLK), .QN(n62115) );
  DFF_X1 \REGISTERS_reg[1][39]  ( .D(n7398), .CK(CLK), .QN(n62116) );
  DFF_X1 \REGISTERS_reg[1][38]  ( .D(n7397), .CK(CLK), .QN(n62117) );
  DFF_X1 \REGISTERS_reg[1][37]  ( .D(n7396), .CK(CLK), .QN(n62118) );
  DFF_X1 \REGISTERS_reg[1][36]  ( .D(n7395), .CK(CLK), .QN(n62119) );
  DFF_X1 \REGISTERS_reg[1][35]  ( .D(n7394), .CK(CLK), .QN(n62120) );
  DFF_X1 \REGISTERS_reg[1][34]  ( .D(n7393), .CK(CLK), .QN(n62121) );
  DFF_X1 \REGISTERS_reg[1][33]  ( .D(n7392), .CK(CLK), .QN(n62122) );
  DFF_X1 \REGISTERS_reg[1][32]  ( .D(n7391), .CK(CLK), .QN(n62123) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n7390), .CK(CLK), .QN(n62124) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n7389), .CK(CLK), .QN(n62125) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n7388), .CK(CLK), .QN(n62126) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n7387), .CK(CLK), .QN(n62127) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n7386), .CK(CLK), .QN(n62128) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n7385), .CK(CLK), .QN(n62129) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n7384), .CK(CLK), .QN(n62130) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n7383), .CK(CLK), .QN(n62131) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n7382), .CK(CLK), .QN(n62132) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n7381), .CK(CLK), .QN(n62133) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n7380), .CK(CLK), .QN(n62134) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n7379), .CK(CLK), .QN(n62135) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n7378), .CK(CLK), .QN(n62136) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n7377), .CK(CLK), .QN(n62137) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n7376), .CK(CLK), .QN(n62138) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n7375), .CK(CLK), .QN(n62139) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n7374), .CK(CLK), .QN(n62140) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n7373), .CK(CLK), .QN(n62141) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n7372), .CK(CLK), .QN(n62142) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n7371), .CK(CLK), .QN(n62143) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n7370), .CK(CLK), .QN(n62144) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n7369), .CK(CLK), .QN(n62145) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n7368), .CK(CLK), .QN(n62146) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n7367), .CK(CLK), .QN(n62147) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n7366), .CK(CLK), .QN(n62148) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n7365), .CK(CLK), .QN(n62149) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n7364), .CK(CLK), .QN(n62150) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n7363), .CK(CLK), .QN(n62151) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n7362), .CK(CLK), .QN(n62152) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n7361), .CK(CLK), .QN(n62153) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n7360), .CK(CLK), .QN(n62154) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n7359), .CK(CLK), .QN(n62155) );
  DFF_X1 \REGISTERS_reg[8][59]  ( .D(n6970), .CK(CLK), .Q(n58366), .QN(n62565)
         );
  DFF_X1 \REGISTERS_reg[8][58]  ( .D(n6969), .CK(CLK), .Q(n58365), .QN(n62566)
         );
  DFF_X1 \REGISTERS_reg[8][57]  ( .D(n6968), .CK(CLK), .Q(n58364), .QN(n62567)
         );
  DFF_X1 \REGISTERS_reg[8][56]  ( .D(n6967), .CK(CLK), .Q(n58363), .QN(n62568)
         );
  DFF_X1 \REGISTERS_reg[8][55]  ( .D(n6966), .CK(CLK), .Q(n58362), .QN(n62569)
         );
  DFF_X1 \REGISTERS_reg[8][54]  ( .D(n6965), .CK(CLK), .Q(n58361), .QN(n62570)
         );
  DFF_X1 \REGISTERS_reg[8][53]  ( .D(n6964), .CK(CLK), .Q(n58360), .QN(n62571)
         );
  DFF_X1 \REGISTERS_reg[8][52]  ( .D(n6963), .CK(CLK), .Q(n58359), .QN(n62572)
         );
  DFF_X1 \REGISTERS_reg[8][51]  ( .D(n6962), .CK(CLK), .Q(n58358), .QN(n62573)
         );
  DFF_X1 \REGISTERS_reg[8][50]  ( .D(n6961), .CK(CLK), .Q(n58357), .QN(n62574)
         );
  DFF_X1 \REGISTERS_reg[8][49]  ( .D(n6960), .CK(CLK), .Q(n58356), .QN(n62575)
         );
  DFF_X1 \REGISTERS_reg[8][48]  ( .D(n6959), .CK(CLK), .Q(n58355), .QN(n62576)
         );
  DFF_X1 \REGISTERS_reg[8][47]  ( .D(n6958), .CK(CLK), .Q(n58354), .QN(n62577)
         );
  DFF_X1 \REGISTERS_reg[8][46]  ( .D(n6957), .CK(CLK), .Q(n58353), .QN(n62578)
         );
  DFF_X1 \REGISTERS_reg[8][45]  ( .D(n6956), .CK(CLK), .Q(n58352), .QN(n62579)
         );
  DFF_X1 \REGISTERS_reg[8][44]  ( .D(n6955), .CK(CLK), .Q(n58351), .QN(n62580)
         );
  DFF_X1 \REGISTERS_reg[8][43]  ( .D(n6954), .CK(CLK), .Q(n58350), .QN(n62581)
         );
  DFF_X1 \REGISTERS_reg[8][42]  ( .D(n6953), .CK(CLK), .Q(n58349), .QN(n62582)
         );
  DFF_X1 \REGISTERS_reg[8][41]  ( .D(n6952), .CK(CLK), .Q(n58348), .QN(n62583)
         );
  DFF_X1 \REGISTERS_reg[8][40]  ( .D(n6951), .CK(CLK), .Q(n58347), .QN(n62584)
         );
  DFF_X1 \REGISTERS_reg[8][39]  ( .D(n6950), .CK(CLK), .Q(n58346), .QN(n62585)
         );
  DFF_X1 \REGISTERS_reg[8][38]  ( .D(n6949), .CK(CLK), .Q(n58345), .QN(n62586)
         );
  DFF_X1 \REGISTERS_reg[8][37]  ( .D(n6948), .CK(CLK), .Q(n58344), .QN(n62587)
         );
  DFF_X1 \REGISTERS_reg[8][36]  ( .D(n6947), .CK(CLK), .Q(n58343), .QN(n62588)
         );
  DFF_X1 \REGISTERS_reg[8][35]  ( .D(n6946), .CK(CLK), .Q(n58342), .QN(n62589)
         );
  DFF_X1 \REGISTERS_reg[8][34]  ( .D(n6945), .CK(CLK), .Q(n58341), .QN(n62590)
         );
  DFF_X1 \REGISTERS_reg[8][33]  ( .D(n6944), .CK(CLK), .Q(n58340), .QN(n62591)
         );
  DFF_X1 \REGISTERS_reg[8][32]  ( .D(n6943), .CK(CLK), .Q(n58339), .QN(n62592)
         );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n6942), .CK(CLK), .Q(n58338), .QN(n62593)
         );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n6941), .CK(CLK), .Q(n58337), .QN(n62594)
         );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n6940), .CK(CLK), .Q(n58336), .QN(n62595)
         );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n6939), .CK(CLK), .Q(n58335), .QN(n62596)
         );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n6938), .CK(CLK), .Q(n58334), .QN(n62597)
         );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n6937), .CK(CLK), .Q(n58333), .QN(n62598)
         );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n6936), .CK(CLK), .Q(n58332), .QN(n62599)
         );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n6935), .CK(CLK), .Q(n58331), .QN(n62600)
         );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n6934), .CK(CLK), .Q(n58330), .QN(n62601)
         );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n6933), .CK(CLK), .Q(n58329), .QN(n62602)
         );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n6932), .CK(CLK), .Q(n58328), .QN(n62603)
         );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n6931), .CK(CLK), .Q(n58327), .QN(n62604)
         );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n6930), .CK(CLK), .Q(n58326), .QN(n62605)
         );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n6929), .CK(CLK), .Q(n58325), .QN(n62606)
         );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n6928), .CK(CLK), .Q(n58324), .QN(n62607)
         );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n6927), .CK(CLK), .Q(n58323), .QN(n62608)
         );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n6926), .CK(CLK), .Q(n58322), .QN(n62609)
         );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n6925), .CK(CLK), .Q(n58321), .QN(n62610)
         );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n6924), .CK(CLK), .Q(n58320), .QN(n62611)
         );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n6923), .CK(CLK), .Q(n58319), .QN(n62612)
         );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n6922), .CK(CLK), .Q(n58318), .QN(n62613)
         );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n6921), .CK(CLK), .Q(n58317), .QN(n62614)
         );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n6920), .CK(CLK), .Q(n58316), .QN(n62615)
         );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n6919), .CK(CLK), .Q(n58315), .QN(n62616)
         );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n6918), .CK(CLK), .Q(n58314), .QN(n62617)
         );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n6917), .CK(CLK), .Q(n58313), .QN(n62618)
         );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n6916), .CK(CLK), .Q(n58312), .QN(n62619)
         );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n6915), .CK(CLK), .Q(n58311), .QN(n62620)
         );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n6914), .CK(CLK), .Q(n58310), .QN(n62621)
         );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n6913), .CK(CLK), .Q(n58309), .QN(n62622)
         );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n6912), .CK(CLK), .Q(n58308), .QN(n62623)
         );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n6911), .CK(CLK), .Q(n58307), .QN(n62624)
         );
  DFF_X1 \REGISTERS_reg[14][59]  ( .D(n6586), .CK(CLK), .Q(n56597), .QN(n62832) );
  DFF_X1 \REGISTERS_reg[14][58]  ( .D(n6585), .CK(CLK), .Q(n56621), .QN(n62833) );
  DFF_X1 \REGISTERS_reg[14][57]  ( .D(n6584), .CK(CLK), .Q(n56645), .QN(n62834) );
  DFF_X1 \REGISTERS_reg[14][56]  ( .D(n6583), .CK(CLK), .Q(n56669), .QN(n62835) );
  DFF_X1 \REGISTERS_reg[14][55]  ( .D(n6582), .CK(CLK), .Q(n56693), .QN(n62836) );
  DFF_X1 \REGISTERS_reg[14][54]  ( .D(n6581), .CK(CLK), .Q(n56717), .QN(n62837) );
  DFF_X1 \REGISTERS_reg[14][53]  ( .D(n6580), .CK(CLK), .Q(n56741), .QN(n62838) );
  DFF_X1 \REGISTERS_reg[14][52]  ( .D(n6579), .CK(CLK), .Q(n56765), .QN(n62839) );
  DFF_X1 \REGISTERS_reg[14][51]  ( .D(n6578), .CK(CLK), .Q(n56789), .QN(n62840) );
  DFF_X1 \REGISTERS_reg[14][50]  ( .D(n6577), .CK(CLK), .Q(n56813), .QN(n62841) );
  DFF_X1 \REGISTERS_reg[14][49]  ( .D(n6576), .CK(CLK), .Q(n56837), .QN(n62842) );
  DFF_X1 \REGISTERS_reg[14][48]  ( .D(n6575), .CK(CLK), .Q(n56861), .QN(n62843) );
  DFF_X1 \REGISTERS_reg[14][47]  ( .D(n6574), .CK(CLK), .Q(n56885), .QN(n62844) );
  DFF_X1 \REGISTERS_reg[14][46]  ( .D(n6573), .CK(CLK), .Q(n56909), .QN(n62845) );
  DFF_X1 \REGISTERS_reg[14][45]  ( .D(n6572), .CK(CLK), .Q(n56933), .QN(n62846) );
  DFF_X1 \REGISTERS_reg[14][44]  ( .D(n6571), .CK(CLK), .Q(n56957), .QN(n62847) );
  DFF_X1 \REGISTERS_reg[14][43]  ( .D(n6570), .CK(CLK), .Q(n56981), .QN(n62848) );
  DFF_X1 \REGISTERS_reg[14][42]  ( .D(n6569), .CK(CLK), .Q(n57005), .QN(n62849) );
  DFF_X1 \REGISTERS_reg[14][41]  ( .D(n6568), .CK(CLK), .Q(n57029), .QN(n62850) );
  DFF_X1 \REGISTERS_reg[14][40]  ( .D(n6567), .CK(CLK), .Q(n57053), .QN(n62851) );
  DFF_X1 \REGISTERS_reg[14][39]  ( .D(n6566), .CK(CLK), .Q(n57077), .QN(n62852) );
  DFF_X1 \REGISTERS_reg[14][38]  ( .D(n6565), .CK(CLK), .Q(n57101), .QN(n62853) );
  DFF_X1 \REGISTERS_reg[14][37]  ( .D(n6564), .CK(CLK), .Q(n57125), .QN(n62854) );
  DFF_X1 \REGISTERS_reg[14][36]  ( .D(n6563), .CK(CLK), .Q(n57149), .QN(n62855) );
  DFF_X1 \REGISTERS_reg[14][35]  ( .D(n6562), .CK(CLK), .Q(n57173), .QN(n62856) );
  DFF_X1 \REGISTERS_reg[14][34]  ( .D(n6561), .CK(CLK), .Q(n57197), .QN(n62857) );
  DFF_X1 \REGISTERS_reg[14][33]  ( .D(n6560), .CK(CLK), .Q(n57221), .QN(n62858) );
  DFF_X1 \REGISTERS_reg[14][32]  ( .D(n6559), .CK(CLK), .Q(n57245), .QN(n62859) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n6558), .CK(CLK), .Q(n57269), .QN(n62860) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n6557), .CK(CLK), .Q(n57293), .QN(n62861) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n6556), .CK(CLK), .Q(n57317), .QN(n62862) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n6555), .CK(CLK), .Q(n57341), .QN(n62863) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n6554), .CK(CLK), .Q(n57365), .QN(n62864) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n6553), .CK(CLK), .Q(n57389), .QN(n62865) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n6552), .CK(CLK), .Q(n57413), .QN(n62866) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n6551), .CK(CLK), .Q(n57437), .QN(n62867) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n6550), .CK(CLK), .Q(n57461), .QN(n62868) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n6549), .CK(CLK), .Q(n57485), .QN(n62869) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n6548), .CK(CLK), .Q(n57509), .QN(n62870) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n6547), .CK(CLK), .Q(n57533), .QN(n62871) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n6546), .CK(CLK), .Q(n57557), .QN(n62872) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n6545), .CK(CLK), .Q(n57581), .QN(n62873) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n6544), .CK(CLK), .Q(n57605), .QN(n62874) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n6543), .CK(CLK), .Q(n57629), .QN(n62875) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n6542), .CK(CLK), .Q(n57653), .QN(n62876) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n6541), .CK(CLK), .Q(n57677), .QN(n62877) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n6540), .CK(CLK), .Q(n57701), .QN(n62878) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n6539), .CK(CLK), .Q(n57725), .QN(n62879) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n6538), .CK(CLK), .Q(n57749), .QN(n62880) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n6537), .CK(CLK), .Q(n57773), .QN(n62881) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n6536), .CK(CLK), .Q(n57797), .QN(n62882)
         );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n6535), .CK(CLK), .Q(n57821), .QN(n62883)
         );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n6534), .CK(CLK), .Q(n57845), .QN(n62884)
         );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n6533), .CK(CLK), .Q(n57869), .QN(n62885)
         );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n6532), .CK(CLK), .Q(n57893), .QN(n62886)
         );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n6531), .CK(CLK), .Q(n57917), .QN(n62887)
         );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n6530), .CK(CLK), .Q(n57941), .QN(n62888)
         );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n6529), .CK(CLK), .Q(n57965), .QN(n62889)
         );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n6528), .CK(CLK), .Q(n57989), .QN(n62890)
         );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n6527), .CK(CLK), .Q(n58013), .QN(n62891)
         );
  DFF_X1 \REGISTERS_reg[13][59]  ( .D(n6650), .CK(CLK), .Q(n56609), .QN(n62766) );
  DFF_X1 \REGISTERS_reg[13][58]  ( .D(n6649), .CK(CLK), .Q(n56633), .QN(n62767) );
  DFF_X1 \REGISTERS_reg[13][57]  ( .D(n6648), .CK(CLK), .Q(n56657), .QN(n62768) );
  DFF_X1 \REGISTERS_reg[13][56]  ( .D(n6647), .CK(CLK), .Q(n56681), .QN(n62769) );
  DFF_X1 \REGISTERS_reg[13][55]  ( .D(n6646), .CK(CLK), .Q(n56705), .QN(n62770) );
  DFF_X1 \REGISTERS_reg[13][54]  ( .D(n6645), .CK(CLK), .Q(n56729), .QN(n62771) );
  DFF_X1 \REGISTERS_reg[13][53]  ( .D(n6644), .CK(CLK), .Q(n56753), .QN(n62772) );
  DFF_X1 \REGISTERS_reg[13][52]  ( .D(n6643), .CK(CLK), .Q(n56777), .QN(n62773) );
  DFF_X1 \REGISTERS_reg[13][51]  ( .D(n6642), .CK(CLK), .Q(n56801), .QN(n62774) );
  DFF_X1 \REGISTERS_reg[13][50]  ( .D(n6641), .CK(CLK), .Q(n56825), .QN(n62775) );
  DFF_X1 \REGISTERS_reg[13][49]  ( .D(n6640), .CK(CLK), .Q(n56849), .QN(n62776) );
  DFF_X1 \REGISTERS_reg[13][48]  ( .D(n6639), .CK(CLK), .Q(n56873), .QN(n62777) );
  DFF_X1 \REGISTERS_reg[13][47]  ( .D(n6638), .CK(CLK), .Q(n56897), .QN(n62778) );
  DFF_X1 \REGISTERS_reg[13][46]  ( .D(n6637), .CK(CLK), .Q(n56921), .QN(n62779) );
  DFF_X1 \REGISTERS_reg[13][45]  ( .D(n6636), .CK(CLK), .Q(n56945), .QN(n62780) );
  DFF_X1 \REGISTERS_reg[13][44]  ( .D(n6635), .CK(CLK), .Q(n56969), .QN(n62781) );
  DFF_X1 \REGISTERS_reg[13][43]  ( .D(n6634), .CK(CLK), .Q(n56993), .QN(n62782) );
  DFF_X1 \REGISTERS_reg[13][42]  ( .D(n6633), .CK(CLK), .Q(n57017), .QN(n62783) );
  DFF_X1 \REGISTERS_reg[13][41]  ( .D(n6632), .CK(CLK), .Q(n57041), .QN(n62784) );
  DFF_X1 \REGISTERS_reg[13][40]  ( .D(n6631), .CK(CLK), .Q(n57065), .QN(n62785) );
  DFF_X1 \REGISTERS_reg[13][39]  ( .D(n6630), .CK(CLK), .Q(n57089), .QN(n62786) );
  DFF_X1 \REGISTERS_reg[13][38]  ( .D(n6629), .CK(CLK), .Q(n57113), .QN(n62787) );
  DFF_X1 \REGISTERS_reg[13][37]  ( .D(n6628), .CK(CLK), .Q(n57137), .QN(n62788) );
  DFF_X1 \REGISTERS_reg[13][36]  ( .D(n6627), .CK(CLK), .Q(n57161), .QN(n62789) );
  DFF_X1 \REGISTERS_reg[13][35]  ( .D(n6626), .CK(CLK), .Q(n57185), .QN(n62790) );
  DFF_X1 \REGISTERS_reg[13][34]  ( .D(n6625), .CK(CLK), .Q(n57209), .QN(n62791) );
  DFF_X1 \REGISTERS_reg[13][33]  ( .D(n6624), .CK(CLK), .Q(n57233), .QN(n62792) );
  DFF_X1 \REGISTERS_reg[13][32]  ( .D(n6623), .CK(CLK), .Q(n57257), .QN(n62793) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n6622), .CK(CLK), .Q(n57281), .QN(n62794) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n6621), .CK(CLK), .Q(n57305), .QN(n62795) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n6620), .CK(CLK), .Q(n57329), .QN(n62796) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n6619), .CK(CLK), .Q(n57353), .QN(n62797) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n6618), .CK(CLK), .Q(n57377), .QN(n62798) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n6617), .CK(CLK), .Q(n57401), .QN(n62799) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n6616), .CK(CLK), .Q(n57425), .QN(n62800) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n6615), .CK(CLK), .Q(n57449), .QN(n62801) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n6614), .CK(CLK), .Q(n57473), .QN(n62802) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n6613), .CK(CLK), .Q(n57497), .QN(n62803) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n6612), .CK(CLK), .Q(n57521), .QN(n62804) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n6611), .CK(CLK), .Q(n57545), .QN(n62805) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n6610), .CK(CLK), .Q(n57569), .QN(n62806) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n6609), .CK(CLK), .Q(n57593), .QN(n62807) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n6608), .CK(CLK), .Q(n57617), .QN(n62808) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n6607), .CK(CLK), .Q(n57641), .QN(n62809) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n6606), .CK(CLK), .Q(n57665), .QN(n62810) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n6605), .CK(CLK), .Q(n57689), .QN(n62811) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n6604), .CK(CLK), .Q(n57713), .QN(n62812) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n6603), .CK(CLK), .Q(n57737), .QN(n62813) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n6602), .CK(CLK), .Q(n57761), .QN(n62814) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n6601), .CK(CLK), .Q(n57785), .QN(n62815) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n6600), .CK(CLK), .Q(n57809), .QN(n62816)
         );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n6599), .CK(CLK), .Q(n57833), .QN(n62817)
         );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n6598), .CK(CLK), .Q(n57857), .QN(n62818)
         );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n6597), .CK(CLK), .Q(n57881), .QN(n62819)
         );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n6596), .CK(CLK), .Q(n57905), .QN(n62820)
         );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n6595), .CK(CLK), .Q(n57929), .QN(n62821)
         );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n6594), .CK(CLK), .Q(n57953), .QN(n62822)
         );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n6593), .CK(CLK), .Q(n57977), .QN(n62823)
         );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n6592), .CK(CLK), .Q(n58001), .QN(n62824)
         );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n6591), .CK(CLK), .Q(n58036), .QN(n62825)
         );
  DFF_X1 \REGISTERS_reg[11][59]  ( .D(n6778), .CK(CLK), .QN(n62702) );
  DFF_X1 \REGISTERS_reg[11][58]  ( .D(n6777), .CK(CLK), .QN(n62703) );
  DFF_X1 \REGISTERS_reg[11][57]  ( .D(n6776), .CK(CLK), .QN(n62704) );
  DFF_X1 \REGISTERS_reg[11][56]  ( .D(n6775), .CK(CLK), .QN(n62705) );
  DFF_X1 \REGISTERS_reg[11][55]  ( .D(n6774), .CK(CLK), .QN(n62706) );
  DFF_X1 \REGISTERS_reg[11][54]  ( .D(n6773), .CK(CLK), .QN(n62707) );
  DFF_X1 \REGISTERS_reg[11][53]  ( .D(n6772), .CK(CLK), .QN(n62708) );
  DFF_X1 \REGISTERS_reg[11][52]  ( .D(n6771), .CK(CLK), .QN(n62709) );
  DFF_X1 \REGISTERS_reg[11][51]  ( .D(n6770), .CK(CLK), .QN(n62710) );
  DFF_X1 \REGISTERS_reg[11][50]  ( .D(n6769), .CK(CLK), .QN(n62711) );
  DFF_X1 \REGISTERS_reg[11][49]  ( .D(n6768), .CK(CLK), .QN(n62712) );
  DFF_X1 \REGISTERS_reg[11][48]  ( .D(n6767), .CK(CLK), .QN(n62713) );
  DFF_X1 \REGISTERS_reg[11][47]  ( .D(n6766), .CK(CLK), .QN(n62714) );
  DFF_X1 \REGISTERS_reg[11][46]  ( .D(n6765), .CK(CLK), .QN(n62715) );
  DFF_X1 \REGISTERS_reg[11][45]  ( .D(n6764), .CK(CLK), .QN(n62716) );
  DFF_X1 \REGISTERS_reg[11][44]  ( .D(n6763), .CK(CLK), .QN(n62717) );
  DFF_X1 \REGISTERS_reg[11][43]  ( .D(n6762), .CK(CLK), .QN(n62718) );
  DFF_X1 \REGISTERS_reg[11][42]  ( .D(n6761), .CK(CLK), .QN(n62719) );
  DFF_X1 \REGISTERS_reg[11][41]  ( .D(n6760), .CK(CLK), .QN(n62720) );
  DFF_X1 \REGISTERS_reg[11][40]  ( .D(n6759), .CK(CLK), .QN(n62721) );
  DFF_X1 \REGISTERS_reg[11][39]  ( .D(n6758), .CK(CLK), .QN(n62722) );
  DFF_X1 \REGISTERS_reg[11][38]  ( .D(n6757), .CK(CLK), .QN(n62723) );
  DFF_X1 \REGISTERS_reg[11][37]  ( .D(n6756), .CK(CLK), .QN(n62724) );
  DFF_X1 \REGISTERS_reg[11][36]  ( .D(n6755), .CK(CLK), .QN(n62725) );
  DFF_X1 \REGISTERS_reg[11][35]  ( .D(n6754), .CK(CLK), .QN(n62726) );
  DFF_X1 \REGISTERS_reg[11][34]  ( .D(n6753), .CK(CLK), .QN(n62727) );
  DFF_X1 \REGISTERS_reg[11][33]  ( .D(n6752), .CK(CLK), .QN(n62728) );
  DFF_X1 \REGISTERS_reg[11][32]  ( .D(n6751), .CK(CLK), .QN(n62729) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n6750), .CK(CLK), .QN(n62730) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n6749), .CK(CLK), .QN(n62731) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n6748), .CK(CLK), .QN(n62732) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n6747), .CK(CLK), .QN(n62733) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n6746), .CK(CLK), .QN(n62734) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n6745), .CK(CLK), .QN(n62735) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n6744), .CK(CLK), .QN(n62736) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n6743), .CK(CLK), .QN(n62737) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n6742), .CK(CLK), .QN(n62738) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n6741), .CK(CLK), .QN(n62739) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n6740), .CK(CLK), .QN(n62740) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n6739), .CK(CLK), .QN(n62741) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n6738), .CK(CLK), .QN(n62742) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n6737), .CK(CLK), .QN(n62743) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n6736), .CK(CLK), .QN(n62744) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n6735), .CK(CLK), .QN(n62745) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n6734), .CK(CLK), .QN(n62746) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n6733), .CK(CLK), .QN(n62747) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n6732), .CK(CLK), .QN(n62748) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n6731), .CK(CLK), .QN(n62749) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n6730), .CK(CLK), .QN(n62750) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n6729), .CK(CLK), .QN(n62751) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n6728), .CK(CLK), .QN(n62752) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n6727), .CK(CLK), .QN(n62753) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n6726), .CK(CLK), .QN(n62754) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n6725), .CK(CLK), .QN(n62755) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n6724), .CK(CLK), .QN(n62756) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n6723), .CK(CLK), .QN(n62757) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n6722), .CK(CLK), .QN(n62758) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n6721), .CK(CLK), .QN(n62759) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n6720), .CK(CLK), .QN(n62760) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n6719), .CK(CLK), .QN(n62761) );
  DFF_X1 \REGISTERS_reg[9][59]  ( .D(n6906), .CK(CLK), .Q(n8899), .QN(n62632)
         );
  DFF_X1 \REGISTERS_reg[9][58]  ( .D(n6905), .CK(CLK), .Q(n8900), .QN(n62633)
         );
  DFF_X1 \REGISTERS_reg[9][57]  ( .D(n6904), .CK(CLK), .Q(n8901), .QN(n62634)
         );
  DFF_X1 \REGISTERS_reg[9][56]  ( .D(n6903), .CK(CLK), .Q(n8902), .QN(n62635)
         );
  DFF_X1 \REGISTERS_reg[9][55]  ( .D(n6902), .CK(CLK), .Q(n8903), .QN(n62636)
         );
  DFF_X1 \REGISTERS_reg[9][54]  ( .D(n6901), .CK(CLK), .Q(n8904), .QN(n62637)
         );
  DFF_X1 \REGISTERS_reg[9][53]  ( .D(n6900), .CK(CLK), .Q(n8905), .QN(n62638)
         );
  DFF_X1 \REGISTERS_reg[9][52]  ( .D(n6899), .CK(CLK), .Q(n8906), .QN(n62639)
         );
  DFF_X1 \REGISTERS_reg[9][51]  ( .D(n6898), .CK(CLK), .Q(n8907), .QN(n62640)
         );
  DFF_X1 \REGISTERS_reg[9][50]  ( .D(n6897), .CK(CLK), .Q(n8908), .QN(n62641)
         );
  DFF_X1 \REGISTERS_reg[9][49]  ( .D(n6896), .CK(CLK), .Q(n8909), .QN(n62642)
         );
  DFF_X1 \REGISTERS_reg[9][48]  ( .D(n6895), .CK(CLK), .Q(n8910), .QN(n62643)
         );
  DFF_X1 \REGISTERS_reg[9][47]  ( .D(n6894), .CK(CLK), .Q(n8911), .QN(n62644)
         );
  DFF_X1 \REGISTERS_reg[9][46]  ( .D(n6893), .CK(CLK), .Q(n8912), .QN(n62645)
         );
  DFF_X1 \REGISTERS_reg[9][45]  ( .D(n6892), .CK(CLK), .Q(n8913), .QN(n62646)
         );
  DFF_X1 \REGISTERS_reg[9][44]  ( .D(n6891), .CK(CLK), .Q(n8914), .QN(n62647)
         );
  DFF_X1 \REGISTERS_reg[9][43]  ( .D(n6890), .CK(CLK), .Q(n8915), .QN(n62648)
         );
  DFF_X1 \REGISTERS_reg[9][42]  ( .D(n6889), .CK(CLK), .Q(n8916), .QN(n62649)
         );
  DFF_X1 \REGISTERS_reg[9][41]  ( .D(n6888), .CK(CLK), .Q(n8917), .QN(n62650)
         );
  DFF_X1 \REGISTERS_reg[9][40]  ( .D(n6887), .CK(CLK), .Q(n8918), .QN(n62651)
         );
  DFF_X1 \REGISTERS_reg[9][39]  ( .D(n6886), .CK(CLK), .Q(n8919), .QN(n62652)
         );
  DFF_X1 \REGISTERS_reg[9][38]  ( .D(n6885), .CK(CLK), .Q(n8920), .QN(n62653)
         );
  DFF_X1 \REGISTERS_reg[9][37]  ( .D(n6884), .CK(CLK), .Q(n8921), .QN(n62654)
         );
  DFF_X1 \REGISTERS_reg[9][36]  ( .D(n6883), .CK(CLK), .Q(n8922), .QN(n62655)
         );
  DFF_X1 \REGISTERS_reg[9][35]  ( .D(n6882), .CK(CLK), .Q(n8923), .QN(n62656)
         );
  DFF_X1 \REGISTERS_reg[9][34]  ( .D(n6881), .CK(CLK), .Q(n8924), .QN(n62657)
         );
  DFF_X1 \REGISTERS_reg[9][33]  ( .D(n6880), .CK(CLK), .Q(n8925), .QN(n62658)
         );
  DFF_X1 \REGISTERS_reg[9][32]  ( .D(n6879), .CK(CLK), .Q(n8926), .QN(n62659)
         );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n6878), .CK(CLK), .Q(n8927), .QN(n62660)
         );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n6877), .CK(CLK), .Q(n8928), .QN(n62661)
         );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n6876), .CK(CLK), .Q(n8929), .QN(n62662)
         );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n6875), .CK(CLK), .Q(n8930), .QN(n62663)
         );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n6874), .CK(CLK), .Q(n8931), .QN(n62664)
         );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n6873), .CK(CLK), .Q(n8932), .QN(n62665)
         );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n6872), .CK(CLK), .Q(n8933), .QN(n62666)
         );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n6871), .CK(CLK), .Q(n8934), .QN(n62667)
         );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n6870), .CK(CLK), .Q(n8935), .QN(n62668)
         );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n6869), .CK(CLK), .Q(n8936), .QN(n62669)
         );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n6868), .CK(CLK), .Q(n8937), .QN(n62670)
         );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n6867), .CK(CLK), .Q(n8938), .QN(n62671)
         );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n6866), .CK(CLK), .Q(n8939), .QN(n62672)
         );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n6865), .CK(CLK), .Q(n8940), .QN(n62673)
         );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n6864), .CK(CLK), .Q(n8941), .QN(n62674)
         );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n6863), .CK(CLK), .Q(n8942), .QN(n62675)
         );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n6862), .CK(CLK), .Q(n8943), .QN(n62676)
         );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n6861), .CK(CLK), .Q(n8944), .QN(n62677)
         );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n6860), .CK(CLK), .Q(n8945), .QN(n62678)
         );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n6859), .CK(CLK), .Q(n8946), .QN(n62679)
         );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n6858), .CK(CLK), .Q(n8947), .QN(n62680)
         );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n6857), .CK(CLK), .Q(n8948), .QN(n62681)
         );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n6856), .CK(CLK), .Q(n8949), .QN(n62682)
         );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n6855), .CK(CLK), .Q(n8950), .QN(n62683)
         );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n6854), .CK(CLK), .Q(n8951), .QN(n62684)
         );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n6853), .CK(CLK), .Q(n8952), .QN(n62685)
         );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n6852), .CK(CLK), .Q(n8953), .QN(n62686)
         );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n6851), .CK(CLK), .Q(n8954), .QN(n62687)
         );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n6850), .CK(CLK), .Q(n8955), .QN(n62688)
         );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n6849), .CK(CLK), .Q(n8956), .QN(n62689)
         );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n6848), .CK(CLK), .Q(n8957), .QN(n62690)
         );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n6847), .CK(CLK), .Q(n8958), .QN(n62691)
         );
  DFF_X1 \REGISTERS_reg[15][59]  ( .D(n6522), .CK(CLK), .Q(n58650), .QN(n62898) );
  DFF_X1 \REGISTERS_reg[15][58]  ( .D(n6521), .CK(CLK), .Q(n58649), .QN(n62899) );
  DFF_X1 \REGISTERS_reg[15][57]  ( .D(n6520), .CK(CLK), .Q(n58648), .QN(n62900) );
  DFF_X1 \REGISTERS_reg[15][56]  ( .D(n6519), .CK(CLK), .Q(n58647), .QN(n62901) );
  DFF_X1 \REGISTERS_reg[15][55]  ( .D(n6518), .CK(CLK), .Q(n58646), .QN(n62902) );
  DFF_X1 \REGISTERS_reg[15][54]  ( .D(n6517), .CK(CLK), .Q(n58645), .QN(n62903) );
  DFF_X1 \REGISTERS_reg[15][53]  ( .D(n6516), .CK(CLK), .Q(n58644), .QN(n62904) );
  DFF_X1 \REGISTERS_reg[15][52]  ( .D(n6515), .CK(CLK), .Q(n58643), .QN(n62905) );
  DFF_X1 \REGISTERS_reg[15][51]  ( .D(n6514), .CK(CLK), .Q(n56791), .QN(n62906) );
  DFF_X1 \REGISTERS_reg[15][50]  ( .D(n6513), .CK(CLK), .Q(n56815), .QN(n62907) );
  DFF_X1 \REGISTERS_reg[15][49]  ( .D(n6512), .CK(CLK), .Q(n56839), .QN(n62908) );
  DFF_X1 \REGISTERS_reg[15][48]  ( .D(n6511), .CK(CLK), .Q(n56863), .QN(n62909) );
  DFF_X1 \REGISTERS_reg[15][47]  ( .D(n6510), .CK(CLK), .Q(n56887), .QN(n62910) );
  DFF_X1 \REGISTERS_reg[15][46]  ( .D(n6509), .CK(CLK), .Q(n56911), .QN(n62911) );
  DFF_X1 \REGISTERS_reg[15][45]  ( .D(n6508), .CK(CLK), .Q(n56935), .QN(n62912) );
  DFF_X1 \REGISTERS_reg[15][44]  ( .D(n6507), .CK(CLK), .Q(n56959), .QN(n62913) );
  DFF_X1 \REGISTERS_reg[15][43]  ( .D(n6506), .CK(CLK), .Q(n56983), .QN(n62914) );
  DFF_X1 \REGISTERS_reg[15][42]  ( .D(n6505), .CK(CLK), .Q(n57007), .QN(n62915) );
  DFF_X1 \REGISTERS_reg[15][41]  ( .D(n6504), .CK(CLK), .Q(n57031), .QN(n62916) );
  DFF_X1 \REGISTERS_reg[15][40]  ( .D(n6503), .CK(CLK), .Q(n57055), .QN(n62917) );
  DFF_X1 \REGISTERS_reg[15][39]  ( .D(n6502), .CK(CLK), .Q(n57079), .QN(n62918) );
  DFF_X1 \REGISTERS_reg[15][38]  ( .D(n6501), .CK(CLK), .Q(n57103), .QN(n62919) );
  DFF_X1 \REGISTERS_reg[15][37]  ( .D(n6500), .CK(CLK), .Q(n57127), .QN(n62920) );
  DFF_X1 \REGISTERS_reg[15][36]  ( .D(n6499), .CK(CLK), .Q(n57151), .QN(n62921) );
  DFF_X1 \REGISTERS_reg[15][35]  ( .D(n6498), .CK(CLK), .Q(n57175), .QN(n62922) );
  DFF_X1 \REGISTERS_reg[15][34]  ( .D(n6497), .CK(CLK), .Q(n57199), .QN(n62923) );
  DFF_X1 \REGISTERS_reg[15][33]  ( .D(n6496), .CK(CLK), .Q(n57223), .QN(n62924) );
  DFF_X1 \REGISTERS_reg[15][32]  ( .D(n6495), .CK(CLK), .Q(n57247), .QN(n62925) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n6494), .CK(CLK), .Q(n57271), .QN(n62926) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n6493), .CK(CLK), .Q(n57295), .QN(n62927) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n6492), .CK(CLK), .Q(n57319), .QN(n62928) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n6491), .CK(CLK), .Q(n57343), .QN(n62929) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n6490), .CK(CLK), .Q(n57367), .QN(n62930) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n6489), .CK(CLK), .Q(n57391), .QN(n62931) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n6488), .CK(CLK), .Q(n57415), .QN(n62932) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n6487), .CK(CLK), .Q(n57439), .QN(n62933) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n6486), .CK(CLK), .Q(n57463), .QN(n62934) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n6485), .CK(CLK), .Q(n57487), .QN(n62935) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n6484), .CK(CLK), .Q(n57511), .QN(n62936) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n6483), .CK(CLK), .Q(n57535), .QN(n62937) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n6482), .CK(CLK), .Q(n57559), .QN(n62938) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n6481), .CK(CLK), .Q(n57583), .QN(n62939) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n6480), .CK(CLK), .Q(n57607), .QN(n62940) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n6479), .CK(CLK), .Q(n57631), .QN(n62941) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n6478), .CK(CLK), .Q(n58642), .QN(n62942) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n6477), .CK(CLK), .Q(n58641), .QN(n62943) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n6476), .CK(CLK), .Q(n58640), .QN(n62944) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n6475), .CK(CLK), .Q(n58639), .QN(n62945) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n6474), .CK(CLK), .Q(n58638), .QN(n62946) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n6473), .CK(CLK), .Q(n58637), .QN(n62947) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n6472), .CK(CLK), .Q(n58636), .QN(n62948)
         );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n6471), .CK(CLK), .Q(n58635), .QN(n62949)
         );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n6470), .CK(CLK), .Q(n58634), .QN(n62950)
         );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n6469), .CK(CLK), .Q(n58633), .QN(n62951)
         );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n6468), .CK(CLK), .Q(n58632), .QN(n62952)
         );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n6467), .CK(CLK), .Q(n58631), .QN(n62953)
         );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n6466), .CK(CLK), .Q(n58630), .QN(n62954)
         );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n6465), .CK(CLK), .Q(n58629), .QN(n62955)
         );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n6464), .CK(CLK), .Q(n58628), .QN(n62956)
         );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n6463), .CK(CLK), .Q(n58627), .QN(n62957)
         );
  DFF_X1 \OUT1_reg[63]  ( .D(n5501), .CK(CLK), .Q(OUT1[63]) );
  DFF_X1 \OUT1_reg[62]  ( .D(n5499), .CK(CLK), .Q(OUT1[62]) );
  DFF_X1 \OUT1_reg[61]  ( .D(n5497), .CK(CLK), .Q(OUT1[61]) );
  DFF_X1 \OUT1_reg[60]  ( .D(n5495), .CK(CLK), .Q(OUT1[60]) );
  NOR3_X1 U45462 ( .A1(n67434), .A2(ADD_RD2[1]), .A3(n66299), .ZN(n66278) );
  NOR3_X1 U45463 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n67434), .ZN(n66281)
         );
  NOR3_X1 U45464 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n67632), .ZN(n65078)
         );
  NOR3_X1 U45465 ( .A1(n67632), .A2(ADD_RD1[1]), .A3(n65099), .ZN(n65086) );
  AND3_X1 U45466 ( .A1(ENABLE), .A2(n68057), .A3(RD1), .ZN(n66494) );
  BUF_X1 U45467 ( .A(n67852), .Z(n67854) );
  BUF_X1 U45468 ( .A(n68256), .Z(n68258) );
  BUF_X1 U45469 ( .A(n67852), .Z(n67855) );
  BUF_X1 U45470 ( .A(n67852), .Z(n67856) );
  BUF_X1 U45471 ( .A(n67853), .Z(n67857) );
  BUF_X1 U45472 ( .A(n67853), .Z(n67858) );
  BUF_X1 U45473 ( .A(n68256), .Z(n68259) );
  BUF_X1 U45474 ( .A(n68256), .Z(n68260) );
  BUF_X1 U45475 ( .A(n68257), .Z(n68261) );
  BUF_X1 U45476 ( .A(n68257), .Z(n68262) );
  BUF_X1 U45477 ( .A(n61959), .Z(n68251) );
  BUF_X1 U45478 ( .A(n61959), .Z(n68252) );
  BUF_X1 U45479 ( .A(n61959), .Z(n68253) );
  BUF_X1 U45480 ( .A(n61959), .Z(n68254) );
  BUF_X1 U45481 ( .A(n65111), .Z(n67440) );
  BUF_X1 U45482 ( .A(n65111), .Z(n67441) );
  BUF_X1 U45483 ( .A(n65111), .Z(n67442) );
  BUF_X1 U45484 ( .A(n65111), .Z(n67443) );
  BUF_X1 U45485 ( .A(n65111), .Z(n67444) );
  BUF_X1 U45486 ( .A(n67891), .Z(n67893) );
  BUF_X1 U45487 ( .A(n67941), .Z(n67943) );
  BUF_X1 U45488 ( .A(n67954), .Z(n67956) );
  BUF_X1 U45489 ( .A(n68045), .Z(n68047) );
  BUF_X1 U45490 ( .A(n68006), .Z(n68008) );
  BUF_X1 U45491 ( .A(n67967), .Z(n67969) );
  BUF_X1 U45492 ( .A(n67801), .Z(n67803) );
  BUF_X1 U45493 ( .A(n67839), .Z(n67841) );
  BUF_X1 U45494 ( .A(n67750), .Z(n67752) );
  BUF_X1 U45495 ( .A(n67737), .Z(n67739) );
  BUF_X1 U45496 ( .A(n67660), .Z(n67662) );
  BUF_X1 U45497 ( .A(n67878), .Z(n67880) );
  BUF_X1 U45498 ( .A(n68032), .Z(n68034) );
  BUF_X1 U45499 ( .A(n68019), .Z(n68021) );
  BUF_X1 U45500 ( .A(n67993), .Z(n67995) );
  BUF_X1 U45501 ( .A(n67814), .Z(n67816) );
  BUF_X1 U45502 ( .A(n67686), .Z(n67688) );
  BUF_X1 U45503 ( .A(n67673), .Z(n67675) );
  BUF_X1 U45504 ( .A(n67980), .Z(n67982) );
  BUF_X1 U45505 ( .A(n67776), .Z(n67778) );
  BUF_X1 U45506 ( .A(n67763), .Z(n67765) );
  BUF_X1 U45507 ( .A(n67712), .Z(n67714) );
  BUF_X1 U45508 ( .A(n67699), .Z(n67701) );
  BUF_X1 U45509 ( .A(n67865), .Z(n67867) );
  BUF_X1 U45510 ( .A(n67916), .Z(n67918) );
  BUF_X1 U45511 ( .A(n67941), .Z(n67944) );
  BUF_X1 U45512 ( .A(n67941), .Z(n67945) );
  BUF_X1 U45513 ( .A(n67942), .Z(n67946) );
  BUF_X1 U45514 ( .A(n67954), .Z(n67957) );
  BUF_X1 U45515 ( .A(n67954), .Z(n67958) );
  BUF_X1 U45516 ( .A(n67955), .Z(n67959) );
  BUF_X1 U45517 ( .A(n68045), .Z(n68048) );
  BUF_X1 U45518 ( .A(n68045), .Z(n68049) );
  BUF_X1 U45519 ( .A(n68046), .Z(n68050) );
  BUF_X1 U45520 ( .A(n68006), .Z(n68009) );
  BUF_X1 U45521 ( .A(n68006), .Z(n68010) );
  BUF_X1 U45522 ( .A(n68007), .Z(n68011) );
  BUF_X1 U45523 ( .A(n67967), .Z(n67970) );
  BUF_X1 U45524 ( .A(n67967), .Z(n67971) );
  BUF_X1 U45525 ( .A(n67968), .Z(n67972) );
  BUF_X1 U45526 ( .A(n67942), .Z(n67947) );
  BUF_X1 U45527 ( .A(n67801), .Z(n67804) );
  BUF_X1 U45528 ( .A(n67801), .Z(n67805) );
  BUF_X1 U45529 ( .A(n67802), .Z(n67806) );
  BUF_X1 U45530 ( .A(n67839), .Z(n67842) );
  BUF_X1 U45531 ( .A(n67839), .Z(n67843) );
  BUF_X1 U45532 ( .A(n67840), .Z(n67844) );
  BUF_X1 U45533 ( .A(n67750), .Z(n67753) );
  BUF_X1 U45534 ( .A(n67750), .Z(n67754) );
  BUF_X1 U45535 ( .A(n67751), .Z(n67755) );
  BUF_X1 U45536 ( .A(n67737), .Z(n67740) );
  BUF_X1 U45537 ( .A(n67737), .Z(n67741) );
  BUF_X1 U45538 ( .A(n67738), .Z(n67742) );
  BUF_X1 U45539 ( .A(n67955), .Z(n67960) );
  BUF_X1 U45540 ( .A(n68046), .Z(n68051) );
  BUF_X1 U45541 ( .A(n68007), .Z(n68012) );
  BUF_X1 U45542 ( .A(n67660), .Z(n67663) );
  BUF_X1 U45543 ( .A(n67660), .Z(n67664) );
  BUF_X1 U45544 ( .A(n67661), .Z(n67665) );
  BUF_X1 U45545 ( .A(n67968), .Z(n67973) );
  BUF_X1 U45546 ( .A(n67802), .Z(n67807) );
  BUF_X1 U45547 ( .A(n67840), .Z(n67845) );
  BUF_X1 U45548 ( .A(n67751), .Z(n67756) );
  BUF_X1 U45549 ( .A(n67738), .Z(n67743) );
  BUF_X1 U45550 ( .A(n67661), .Z(n67666) );
  BUF_X1 U45551 ( .A(n67878), .Z(n67881) );
  BUF_X1 U45552 ( .A(n67878), .Z(n67882) );
  BUF_X1 U45553 ( .A(n67879), .Z(n67883) );
  BUF_X1 U45554 ( .A(n68032), .Z(n68035) );
  BUF_X1 U45555 ( .A(n68032), .Z(n68036) );
  BUF_X1 U45556 ( .A(n68033), .Z(n68037) );
  BUF_X1 U45557 ( .A(n68019), .Z(n68022) );
  BUF_X1 U45558 ( .A(n68019), .Z(n68023) );
  BUF_X1 U45559 ( .A(n68020), .Z(n68024) );
  BUF_X1 U45560 ( .A(n67993), .Z(n67996) );
  BUF_X1 U45561 ( .A(n67993), .Z(n67997) );
  BUF_X1 U45562 ( .A(n67994), .Z(n67998) );
  BUF_X1 U45563 ( .A(n67814), .Z(n67817) );
  BUF_X1 U45564 ( .A(n67814), .Z(n67818) );
  BUF_X1 U45565 ( .A(n67815), .Z(n67819) );
  BUF_X1 U45566 ( .A(n67686), .Z(n67689) );
  BUF_X1 U45567 ( .A(n67686), .Z(n67690) );
  BUF_X1 U45568 ( .A(n67687), .Z(n67691) );
  BUF_X1 U45569 ( .A(n67673), .Z(n67676) );
  BUF_X1 U45570 ( .A(n67673), .Z(n67677) );
  BUF_X1 U45571 ( .A(n67674), .Z(n67678) );
  BUF_X1 U45572 ( .A(n67879), .Z(n67884) );
  BUF_X1 U45573 ( .A(n68033), .Z(n68038) );
  BUF_X1 U45574 ( .A(n68020), .Z(n68025) );
  BUF_X1 U45575 ( .A(n67994), .Z(n67999) );
  BUF_X1 U45576 ( .A(n67815), .Z(n67820) );
  BUF_X1 U45577 ( .A(n67687), .Z(n67692) );
  BUF_X1 U45578 ( .A(n67674), .Z(n67679) );
  BUF_X1 U45579 ( .A(n67980), .Z(n67983) );
  BUF_X1 U45580 ( .A(n67980), .Z(n67984) );
  BUF_X1 U45581 ( .A(n67981), .Z(n67985) );
  BUF_X1 U45582 ( .A(n67776), .Z(n67779) );
  BUF_X1 U45583 ( .A(n67776), .Z(n67780) );
  BUF_X1 U45584 ( .A(n67777), .Z(n67781) );
  BUF_X1 U45585 ( .A(n67763), .Z(n67766) );
  BUF_X1 U45586 ( .A(n67763), .Z(n67767) );
  BUF_X1 U45587 ( .A(n67764), .Z(n67768) );
  BUF_X1 U45588 ( .A(n67712), .Z(n67715) );
  BUF_X1 U45589 ( .A(n67712), .Z(n67716) );
  BUF_X1 U45590 ( .A(n67713), .Z(n67717) );
  BUF_X1 U45591 ( .A(n67699), .Z(n67702) );
  BUF_X1 U45592 ( .A(n67699), .Z(n67703) );
  BUF_X1 U45593 ( .A(n67700), .Z(n67704) );
  BUF_X1 U45594 ( .A(n67981), .Z(n67986) );
  BUF_X1 U45595 ( .A(n67777), .Z(n67782) );
  BUF_X1 U45596 ( .A(n67764), .Z(n67769) );
  BUF_X1 U45597 ( .A(n67713), .Z(n67718) );
  BUF_X1 U45598 ( .A(n67700), .Z(n67705) );
  BUF_X1 U45599 ( .A(n67865), .Z(n67868) );
  BUF_X1 U45600 ( .A(n67865), .Z(n67869) );
  BUF_X1 U45601 ( .A(n67866), .Z(n67870) );
  BUF_X1 U45602 ( .A(n67866), .Z(n67871) );
  BUF_X1 U45603 ( .A(n67892), .Z(n67897) );
  BUF_X1 U45604 ( .A(n67892), .Z(n67896) );
  BUF_X1 U45605 ( .A(n67891), .Z(n67895) );
  BUF_X1 U45606 ( .A(n67891), .Z(n67894) );
  BUF_X1 U45607 ( .A(n67916), .Z(n67919) );
  BUF_X1 U45608 ( .A(n67916), .Z(n67920) );
  BUF_X1 U45609 ( .A(n67917), .Z(n67921) );
  BUF_X1 U45610 ( .A(n67917), .Z(n67922) );
  BUF_X1 U45611 ( .A(n62092), .Z(n68039) );
  BUF_X1 U45612 ( .A(n62092), .Z(n68040) );
  BUF_X1 U45613 ( .A(n62092), .Z(n68041) );
  BUF_X1 U45614 ( .A(n62092), .Z(n68042) );
  BUF_X1 U45615 ( .A(n62092), .Z(n68043) );
  BUF_X1 U45616 ( .A(n63766), .Z(n67654) );
  BUF_X1 U45617 ( .A(n63766), .Z(n67655) );
  BUF_X1 U45618 ( .A(n63766), .Z(n67656) );
  BUF_X1 U45619 ( .A(n63766), .Z(n67657) );
  BUF_X1 U45620 ( .A(n63766), .Z(n67658) );
  BUF_X1 U45621 ( .A(n62159), .Z(n68026) );
  BUF_X1 U45622 ( .A(n62159), .Z(n68027) );
  BUF_X1 U45623 ( .A(n62159), .Z(n68028) );
  BUF_X1 U45624 ( .A(n62159), .Z(n68029) );
  BUF_X1 U45625 ( .A(n62159), .Z(n68030) );
  BUF_X1 U45626 ( .A(n62628), .Z(n67935) );
  BUF_X1 U45627 ( .A(n62628), .Z(n67936) );
  BUF_X1 U45628 ( .A(n62628), .Z(n67937) );
  BUF_X1 U45629 ( .A(n62628), .Z(n67938) );
  BUF_X1 U45630 ( .A(n62628), .Z(n67939) );
  BUF_X1 U45631 ( .A(n62561), .Z(n67948) );
  BUF_X1 U45632 ( .A(n62561), .Z(n67949) );
  BUF_X1 U45633 ( .A(n62561), .Z(n67950) );
  BUF_X1 U45634 ( .A(n62561), .Z(n67951) );
  BUF_X1 U45635 ( .A(n62561), .Z(n67952) );
  BUF_X1 U45636 ( .A(n62695), .Z(n67923) );
  BUF_X1 U45637 ( .A(n62695), .Z(n67924) );
  BUF_X1 U45638 ( .A(n62695), .Z(n67925) );
  BUF_X1 U45639 ( .A(n62695), .Z(n67926) );
  BUF_X1 U45640 ( .A(n62695), .Z(n67927) );
  BUF_X1 U45641 ( .A(n62292), .Z(n68000) );
  BUF_X1 U45642 ( .A(n62292), .Z(n68001) );
  BUF_X1 U45643 ( .A(n62292), .Z(n68002) );
  BUF_X1 U45644 ( .A(n62292), .Z(n68003) );
  BUF_X1 U45645 ( .A(n62292), .Z(n68004) );
  BUF_X1 U45646 ( .A(n62495), .Z(n67961) );
  BUF_X1 U45647 ( .A(n62495), .Z(n67962) );
  BUF_X1 U45648 ( .A(n62495), .Z(n67963) );
  BUF_X1 U45649 ( .A(n62495), .Z(n67964) );
  BUF_X1 U45650 ( .A(n62495), .Z(n67965) );
  BUF_X1 U45651 ( .A(n63163), .Z(n67795) );
  BUF_X1 U45652 ( .A(n63163), .Z(n67796) );
  BUF_X1 U45653 ( .A(n63163), .Z(n67797) );
  BUF_X1 U45654 ( .A(n63163), .Z(n67798) );
  BUF_X1 U45655 ( .A(n63163), .Z(n67799) );
  BUF_X1 U45656 ( .A(n62961), .Z(n67846) );
  BUF_X1 U45657 ( .A(n62961), .Z(n67847) );
  BUF_X1 U45658 ( .A(n62961), .Z(n67848) );
  BUF_X1 U45659 ( .A(n62961), .Z(n67849) );
  BUF_X1 U45660 ( .A(n62961), .Z(n67850) );
  BUF_X1 U45661 ( .A(n63028), .Z(n67833) );
  BUF_X1 U45662 ( .A(n63028), .Z(n67834) );
  BUF_X1 U45663 ( .A(n63028), .Z(n67835) );
  BUF_X1 U45664 ( .A(n63028), .Z(n67836) );
  BUF_X1 U45665 ( .A(n63028), .Z(n67837) );
  BUF_X1 U45666 ( .A(n63364), .Z(n67744) );
  BUF_X1 U45667 ( .A(n63364), .Z(n67745) );
  BUF_X1 U45668 ( .A(n63364), .Z(n67746) );
  BUF_X1 U45669 ( .A(n63364), .Z(n67747) );
  BUF_X1 U45670 ( .A(n63364), .Z(n67748) );
  BUF_X1 U45671 ( .A(n63431), .Z(n67731) );
  BUF_X1 U45672 ( .A(n63431), .Z(n67732) );
  BUF_X1 U45673 ( .A(n63431), .Z(n67733) );
  BUF_X1 U45674 ( .A(n63431), .Z(n67734) );
  BUF_X1 U45675 ( .A(n63431), .Z(n67735) );
  BUF_X1 U45676 ( .A(n63499), .Z(n67719) );
  BUF_X1 U45677 ( .A(n63499), .Z(n67720) );
  BUF_X1 U45678 ( .A(n63499), .Z(n67721) );
  BUF_X1 U45679 ( .A(n63499), .Z(n67722) );
  BUF_X1 U45680 ( .A(n63499), .Z(n67723) );
  BUF_X1 U45681 ( .A(n62763), .Z(n67898) );
  BUF_X1 U45682 ( .A(n62763), .Z(n67899) );
  BUF_X1 U45683 ( .A(n62763), .Z(n67900) );
  BUF_X1 U45684 ( .A(n62763), .Z(n67901) );
  BUF_X1 U45685 ( .A(n62763), .Z(n67902) );
  BUF_X1 U45686 ( .A(n62828), .Z(n67872) );
  BUF_X1 U45687 ( .A(n62828), .Z(n67873) );
  BUF_X1 U45688 ( .A(n62828), .Z(n67874) );
  BUF_X1 U45689 ( .A(n62828), .Z(n67875) );
  BUF_X1 U45690 ( .A(n62828), .Z(n67876) );
  BUF_X1 U45691 ( .A(n62226), .Z(n68013) );
  BUF_X1 U45692 ( .A(n62226), .Z(n68014) );
  BUF_X1 U45693 ( .A(n62226), .Z(n68015) );
  BUF_X1 U45694 ( .A(n62226), .Z(n68016) );
  BUF_X1 U45695 ( .A(n62226), .Z(n68017) );
  BUF_X1 U45696 ( .A(n62359), .Z(n67987) );
  BUF_X1 U45697 ( .A(n62359), .Z(n67988) );
  BUF_X1 U45698 ( .A(n62359), .Z(n67989) );
  BUF_X1 U45699 ( .A(n62359), .Z(n67990) );
  BUF_X1 U45700 ( .A(n62359), .Z(n67991) );
  BUF_X1 U45701 ( .A(n63097), .Z(n67808) );
  BUF_X1 U45702 ( .A(n63097), .Z(n67809) );
  BUF_X1 U45703 ( .A(n63097), .Z(n67810) );
  BUF_X1 U45704 ( .A(n63097), .Z(n67811) );
  BUF_X1 U45705 ( .A(n63097), .Z(n67812) );
  BUF_X1 U45706 ( .A(n63634), .Z(n67680) );
  BUF_X1 U45707 ( .A(n63634), .Z(n67681) );
  BUF_X1 U45708 ( .A(n63634), .Z(n67682) );
  BUF_X1 U45709 ( .A(n63634), .Z(n67683) );
  BUF_X1 U45710 ( .A(n63634), .Z(n67684) );
  BUF_X1 U45711 ( .A(n63700), .Z(n67667) );
  BUF_X1 U45712 ( .A(n63700), .Z(n67668) );
  BUF_X1 U45713 ( .A(n63700), .Z(n67669) );
  BUF_X1 U45714 ( .A(n63700), .Z(n67670) );
  BUF_X1 U45715 ( .A(n63700), .Z(n67671) );
  BUF_X1 U45716 ( .A(n62425), .Z(n67974) );
  BUF_X1 U45717 ( .A(n62425), .Z(n67975) );
  BUF_X1 U45718 ( .A(n62425), .Z(n67976) );
  BUF_X1 U45719 ( .A(n62425), .Z(n67977) );
  BUF_X1 U45720 ( .A(n62425), .Z(n67978) );
  BUF_X1 U45721 ( .A(n63094), .Z(n67821) );
  BUF_X1 U45722 ( .A(n63094), .Z(n67822) );
  BUF_X1 U45723 ( .A(n63094), .Z(n67823) );
  BUF_X1 U45724 ( .A(n63094), .Z(n67824) );
  BUF_X1 U45725 ( .A(n63094), .Z(n67825) );
  BUF_X1 U45726 ( .A(n63231), .Z(n67770) );
  BUF_X1 U45727 ( .A(n63231), .Z(n67771) );
  BUF_X1 U45728 ( .A(n63231), .Z(n67772) );
  BUF_X1 U45729 ( .A(n63231), .Z(n67773) );
  BUF_X1 U45730 ( .A(n63231), .Z(n67774) );
  BUF_X1 U45731 ( .A(n63228), .Z(n67783) );
  BUF_X1 U45732 ( .A(n63228), .Z(n67784) );
  BUF_X1 U45733 ( .A(n63228), .Z(n67785) );
  BUF_X1 U45734 ( .A(n63228), .Z(n67786) );
  BUF_X1 U45735 ( .A(n63228), .Z(n67787) );
  BUF_X1 U45736 ( .A(n63298), .Z(n67757) );
  BUF_X1 U45737 ( .A(n63298), .Z(n67758) );
  BUF_X1 U45738 ( .A(n63298), .Z(n67759) );
  BUF_X1 U45739 ( .A(n63298), .Z(n67760) );
  BUF_X1 U45740 ( .A(n63298), .Z(n67761) );
  BUF_X1 U45741 ( .A(n63502), .Z(n67706) );
  BUF_X1 U45742 ( .A(n63502), .Z(n67707) );
  BUF_X1 U45743 ( .A(n63502), .Z(n67708) );
  BUF_X1 U45744 ( .A(n63502), .Z(n67709) );
  BUF_X1 U45745 ( .A(n63502), .Z(n67710) );
  BUF_X1 U45746 ( .A(n63568), .Z(n67693) );
  BUF_X1 U45747 ( .A(n63568), .Z(n67694) );
  BUF_X1 U45748 ( .A(n63568), .Z(n67695) );
  BUF_X1 U45749 ( .A(n63568), .Z(n67696) );
  BUF_X1 U45750 ( .A(n63568), .Z(n67697) );
  BUF_X1 U45751 ( .A(n62894), .Z(n67859) );
  BUF_X1 U45752 ( .A(n62894), .Z(n67860) );
  BUF_X1 U45753 ( .A(n62894), .Z(n67861) );
  BUF_X1 U45754 ( .A(n62894), .Z(n67862) );
  BUF_X1 U45755 ( .A(n62894), .Z(n67863) );
  BUF_X1 U45756 ( .A(n62765), .Z(n67885) );
  BUF_X1 U45757 ( .A(n62765), .Z(n67886) );
  BUF_X1 U45758 ( .A(n62765), .Z(n67887) );
  BUF_X1 U45759 ( .A(n62765), .Z(n67888) );
  BUF_X1 U45760 ( .A(n62765), .Z(n67889) );
  BUF_X1 U45761 ( .A(n62698), .Z(n67910) );
  BUF_X1 U45762 ( .A(n62698), .Z(n67911) );
  BUF_X1 U45763 ( .A(n62698), .Z(n67912) );
  BUF_X1 U45764 ( .A(n62698), .Z(n67913) );
  BUF_X1 U45765 ( .A(n62698), .Z(n67914) );
  BUF_X1 U45766 ( .A(n61959), .Z(n68250) );
  BUF_X1 U45767 ( .A(n61957), .Z(n68256) );
  BUF_X1 U45768 ( .A(n62959), .Z(n67852) );
  BUF_X1 U45769 ( .A(n61957), .Z(n68257) );
  BUF_X1 U45770 ( .A(n62959), .Z(n67853) );
  INV_X1 U45771 ( .A(n66494), .ZN(n67632) );
  INV_X1 U45772 ( .A(n66494), .ZN(n67633) );
  INV_X1 U45773 ( .A(n66494), .ZN(n67634) );
  INV_X1 U45774 ( .A(n66494), .ZN(n67635) );
  BUF_X1 U45775 ( .A(n63790), .Z(n67588) );
  BUF_X1 U45776 ( .A(n65146), .Z(n67278) );
  BUF_X1 U45777 ( .A(n65146), .Z(n67279) );
  BUF_X1 U45778 ( .A(n65146), .Z(n67280) );
  BUF_X1 U45779 ( .A(n65146), .Z(n67281) );
  BUF_X1 U45780 ( .A(n65146), .Z(n67282) );
  BUF_X1 U45781 ( .A(n65141), .Z(n67302) );
  BUF_X1 U45782 ( .A(n65141), .Z(n67303) );
  BUF_X1 U45783 ( .A(n65141), .Z(n67304) );
  BUF_X1 U45784 ( .A(n65141), .Z(n67305) );
  BUF_X1 U45785 ( .A(n65141), .Z(n67306) );
  BUF_X1 U45786 ( .A(n63815), .Z(n67476) );
  BUF_X1 U45787 ( .A(n63815), .Z(n67477) );
  BUF_X1 U45788 ( .A(n63815), .Z(n67478) );
  BUF_X1 U45789 ( .A(n63815), .Z(n67479) );
  BUF_X1 U45790 ( .A(n63815), .Z(n67480) );
  BUF_X1 U45791 ( .A(n63810), .Z(n67500) );
  BUF_X1 U45792 ( .A(n63810), .Z(n67501) );
  BUF_X1 U45793 ( .A(n63810), .Z(n67502) );
  BUF_X1 U45794 ( .A(n63810), .Z(n67503) );
  BUF_X1 U45795 ( .A(n63810), .Z(n67504) );
  BUF_X1 U45796 ( .A(n65116), .Z(n67416) );
  BUF_X1 U45797 ( .A(n65121), .Z(n67392) );
  BUF_X1 U45798 ( .A(n65126), .Z(n67368) );
  BUF_X1 U45799 ( .A(n65116), .Z(n67417) );
  BUF_X1 U45800 ( .A(n65121), .Z(n67393) );
  BUF_X1 U45801 ( .A(n65126), .Z(n67369) );
  BUF_X1 U45802 ( .A(n65116), .Z(n67418) );
  BUF_X1 U45803 ( .A(n65121), .Z(n67394) );
  BUF_X1 U45804 ( .A(n65126), .Z(n67370) );
  BUF_X1 U45805 ( .A(n65116), .Z(n67419) );
  BUF_X1 U45806 ( .A(n65121), .Z(n67395) );
  BUF_X1 U45807 ( .A(n65126), .Z(n67371) );
  BUF_X1 U45808 ( .A(n65116), .Z(n67420) );
  BUF_X1 U45809 ( .A(n65121), .Z(n67396) );
  BUF_X1 U45810 ( .A(n65126), .Z(n67372) );
  BUF_X1 U45811 ( .A(n63794), .Z(n67566) );
  BUF_X1 U45812 ( .A(n63788), .Z(n67590) );
  BUF_X1 U45813 ( .A(n63794), .Z(n67567) );
  BUF_X1 U45814 ( .A(n63788), .Z(n67591) );
  BUF_X1 U45815 ( .A(n63794), .Z(n67568) );
  BUF_X1 U45816 ( .A(n63788), .Z(n67592) );
  BUF_X1 U45817 ( .A(n63794), .Z(n67569) );
  BUF_X1 U45818 ( .A(n63788), .Z(n67593) );
  BUF_X1 U45819 ( .A(n63794), .Z(n67570) );
  BUF_X1 U45820 ( .A(n63788), .Z(n67594) );
  BUF_X1 U45821 ( .A(n63778), .Z(n67636) );
  BUF_X1 U45822 ( .A(n63783), .Z(n67614) );
  BUF_X1 U45823 ( .A(n63778), .Z(n67637) );
  BUF_X1 U45824 ( .A(n63783), .Z(n67615) );
  BUF_X1 U45825 ( .A(n63778), .Z(n67638) );
  BUF_X1 U45826 ( .A(n63783), .Z(n67616) );
  BUF_X1 U45827 ( .A(n63778), .Z(n67639) );
  BUF_X1 U45828 ( .A(n63783), .Z(n67617) );
  BUF_X1 U45829 ( .A(n63778), .Z(n67640) );
  BUF_X1 U45830 ( .A(n63783), .Z(n67618) );
  BUF_X1 U45831 ( .A(n65142), .Z(n67296) );
  BUF_X1 U45832 ( .A(n65147), .Z(n67272) );
  BUF_X1 U45833 ( .A(n65142), .Z(n67297) );
  BUF_X1 U45834 ( .A(n65147), .Z(n67273) );
  BUF_X1 U45835 ( .A(n65142), .Z(n67298) );
  BUF_X1 U45836 ( .A(n65147), .Z(n67274) );
  BUF_X1 U45837 ( .A(n65142), .Z(n67299) );
  BUF_X1 U45838 ( .A(n65147), .Z(n67275) );
  BUF_X1 U45839 ( .A(n65142), .Z(n67300) );
  BUF_X1 U45840 ( .A(n65147), .Z(n67276) );
  BUF_X1 U45841 ( .A(n63811), .Z(n67494) );
  BUF_X1 U45842 ( .A(n63816), .Z(n67470) );
  BUF_X1 U45843 ( .A(n63811), .Z(n67495) );
  BUF_X1 U45844 ( .A(n63816), .Z(n67471) );
  BUF_X1 U45845 ( .A(n63811), .Z(n67496) );
  BUF_X1 U45846 ( .A(n63816), .Z(n67472) );
  BUF_X1 U45847 ( .A(n63811), .Z(n67497) );
  BUF_X1 U45848 ( .A(n63816), .Z(n67473) );
  BUF_X1 U45849 ( .A(n63811), .Z(n67498) );
  BUF_X1 U45850 ( .A(n63816), .Z(n67474) );
  BUF_X1 U45851 ( .A(n65113), .Z(n67429) );
  BUF_X1 U45852 ( .A(n65113), .Z(n67430) );
  BUF_X1 U45853 ( .A(n65113), .Z(n67431) );
  BUF_X1 U45854 ( .A(n65113), .Z(n67432) );
  BUF_X1 U45855 ( .A(n65108), .Z(n67453) );
  BUF_X1 U45856 ( .A(n65118), .Z(n67405) );
  BUF_X1 U45857 ( .A(n65123), .Z(n67381) );
  BUF_X1 U45858 ( .A(n65108), .Z(n67454) );
  BUF_X1 U45859 ( .A(n65118), .Z(n67406) );
  BUF_X1 U45860 ( .A(n65123), .Z(n67382) );
  BUF_X1 U45861 ( .A(n65108), .Z(n67455) );
  BUF_X1 U45862 ( .A(n65118), .Z(n67407) );
  BUF_X1 U45863 ( .A(n65123), .Z(n67383) );
  BUF_X1 U45864 ( .A(n65108), .Z(n67456) );
  BUF_X1 U45865 ( .A(n65118), .Z(n67408) );
  BUF_X1 U45866 ( .A(n65123), .Z(n67384) );
  BUF_X1 U45867 ( .A(n63775), .Z(n67649) );
  BUF_X1 U45868 ( .A(n63775), .Z(n67650) );
  BUF_X1 U45869 ( .A(n63775), .Z(n67651) );
  BUF_X1 U45870 ( .A(n63775), .Z(n67652) );
  BUF_X1 U45871 ( .A(n63791), .Z(n67579) );
  BUF_X1 U45872 ( .A(n63785), .Z(n67603) );
  BUF_X1 U45873 ( .A(n63780), .Z(n67627) );
  BUF_X1 U45874 ( .A(n63791), .Z(n67580) );
  BUF_X1 U45875 ( .A(n63785), .Z(n67604) );
  BUF_X1 U45876 ( .A(n63780), .Z(n67628) );
  BUF_X1 U45877 ( .A(n63791), .Z(n67581) );
  BUF_X1 U45878 ( .A(n63785), .Z(n67605) );
  BUF_X1 U45879 ( .A(n63780), .Z(n67629) );
  BUF_X1 U45880 ( .A(n63791), .Z(n67582) );
  BUF_X1 U45881 ( .A(n63785), .Z(n67606) );
  BUF_X1 U45882 ( .A(n63780), .Z(n67630) );
  BUF_X1 U45883 ( .A(n65140), .Z(n67308) );
  BUF_X1 U45884 ( .A(n65140), .Z(n67309) );
  BUF_X1 U45885 ( .A(n65140), .Z(n67310) );
  BUF_X1 U45886 ( .A(n65140), .Z(n67311) );
  BUF_X1 U45887 ( .A(n65140), .Z(n67312) );
  BUF_X1 U45888 ( .A(n63809), .Z(n67506) );
  BUF_X1 U45889 ( .A(n63809), .Z(n67507) );
  BUF_X1 U45890 ( .A(n63809), .Z(n67508) );
  BUF_X1 U45891 ( .A(n63809), .Z(n67509) );
  BUF_X1 U45892 ( .A(n63809), .Z(n67510) );
  BUF_X1 U45893 ( .A(n63807), .Z(n67518) );
  BUF_X1 U45894 ( .A(n63807), .Z(n67519) );
  BUF_X1 U45895 ( .A(n63807), .Z(n67520) );
  BUF_X1 U45896 ( .A(n63807), .Z(n67521) );
  BUF_X1 U45897 ( .A(n63807), .Z(n67522) );
  BUF_X1 U45898 ( .A(n65138), .Z(n67320) );
  BUF_X1 U45899 ( .A(n65138), .Z(n67321) );
  BUF_X1 U45900 ( .A(n65138), .Z(n67322) );
  BUF_X1 U45901 ( .A(n65138), .Z(n67323) );
  BUF_X1 U45902 ( .A(n65138), .Z(n67324) );
  BUF_X1 U45903 ( .A(n65139), .Z(n67314) );
  BUF_X1 U45904 ( .A(n65139), .Z(n67315) );
  BUF_X1 U45905 ( .A(n65139), .Z(n67316) );
  BUF_X1 U45906 ( .A(n65139), .Z(n67317) );
  BUF_X1 U45907 ( .A(n65139), .Z(n67318) );
  BUF_X1 U45908 ( .A(n63808), .Z(n67512) );
  BUF_X1 U45909 ( .A(n63808), .Z(n67513) );
  BUF_X1 U45910 ( .A(n63808), .Z(n67514) );
  BUF_X1 U45911 ( .A(n63808), .Z(n67515) );
  BUF_X1 U45912 ( .A(n63808), .Z(n67516) );
  BUF_X1 U45913 ( .A(n65117), .Z(n67410) );
  BUF_X1 U45914 ( .A(n65117), .Z(n67411) );
  BUF_X1 U45915 ( .A(n65117), .Z(n67412) );
  BUF_X1 U45916 ( .A(n65117), .Z(n67413) );
  BUF_X1 U45917 ( .A(n65117), .Z(n67414) );
  BUF_X1 U45918 ( .A(n65122), .Z(n67386) );
  BUF_X1 U45919 ( .A(n65127), .Z(n67362) );
  BUF_X1 U45920 ( .A(n65122), .Z(n67387) );
  BUF_X1 U45921 ( .A(n65127), .Z(n67363) );
  BUF_X1 U45922 ( .A(n65122), .Z(n67388) );
  BUF_X1 U45923 ( .A(n65127), .Z(n67364) );
  BUF_X1 U45924 ( .A(n65122), .Z(n67389) );
  BUF_X1 U45925 ( .A(n65127), .Z(n67365) );
  BUF_X1 U45926 ( .A(n65122), .Z(n67390) );
  BUF_X1 U45927 ( .A(n65127), .Z(n67366) );
  BUF_X1 U45928 ( .A(n63795), .Z(n67560) );
  BUF_X1 U45929 ( .A(n63795), .Z(n67561) );
  BUF_X1 U45930 ( .A(n63795), .Z(n67562) );
  BUF_X1 U45931 ( .A(n63795), .Z(n67563) );
  BUF_X1 U45932 ( .A(n63795), .Z(n67564) );
  BUF_X1 U45933 ( .A(n63784), .Z(n67608) );
  BUF_X1 U45934 ( .A(n63784), .Z(n67609) );
  BUF_X1 U45935 ( .A(n63784), .Z(n67610) );
  BUF_X1 U45936 ( .A(n63784), .Z(n67611) );
  BUF_X1 U45937 ( .A(n63784), .Z(n67612) );
  NAND2_X1 U45938 ( .A1(n68057), .A2(n68047), .ZN(n62092) );
  NAND2_X1 U45939 ( .A1(n68057), .A2(n67662), .ZN(n63766) );
  NAND2_X1 U45940 ( .A1(n68057), .A2(n68034), .ZN(n62159) );
  BUF_X1 U45941 ( .A(n63790), .Z(n67584) );
  BUF_X1 U45942 ( .A(n63790), .Z(n67585) );
  BUF_X1 U45943 ( .A(n63790), .Z(n67586) );
  BUF_X1 U45944 ( .A(n63790), .Z(n67587) );
  BUF_X1 U45945 ( .A(n62693), .Z(n67929) );
  BUF_X1 U45946 ( .A(n63498), .Z(n67725) );
  BUF_X1 U45947 ( .A(n62762), .Z(n67904) );
  BUF_X1 U45948 ( .A(n63093), .Z(n67827) );
  BUF_X1 U45949 ( .A(n63227), .Z(n67789) );
  BUF_X1 U45950 ( .A(n62693), .Z(n67930) );
  BUF_X1 U45951 ( .A(n62693), .Z(n67931) );
  BUF_X1 U45952 ( .A(n62693), .Z(n67932) );
  BUF_X1 U45953 ( .A(n62693), .Z(n67933) );
  BUF_X1 U45954 ( .A(n63498), .Z(n67726) );
  BUF_X1 U45955 ( .A(n63498), .Z(n67727) );
  BUF_X1 U45956 ( .A(n63498), .Z(n67728) );
  BUF_X1 U45957 ( .A(n63498), .Z(n67729) );
  BUF_X1 U45958 ( .A(n62762), .Z(n67905) );
  BUF_X1 U45959 ( .A(n62762), .Z(n67906) );
  BUF_X1 U45960 ( .A(n62762), .Z(n67907) );
  BUF_X1 U45961 ( .A(n62762), .Z(n67908) );
  BUF_X1 U45962 ( .A(n63093), .Z(n67828) );
  BUF_X1 U45963 ( .A(n63093), .Z(n67829) );
  BUF_X1 U45964 ( .A(n63093), .Z(n67830) );
  BUF_X1 U45965 ( .A(n63093), .Z(n67831) );
  BUF_X1 U45966 ( .A(n63227), .Z(n67790) );
  BUF_X1 U45967 ( .A(n63227), .Z(n67791) );
  BUF_X1 U45968 ( .A(n63227), .Z(n67792) );
  BUF_X1 U45969 ( .A(n63227), .Z(n67793) );
  BUF_X1 U45970 ( .A(n65132), .Z(n67356) );
  BUF_X1 U45971 ( .A(n65134), .Z(n67344) );
  BUF_X1 U45972 ( .A(n65132), .Z(n67357) );
  BUF_X1 U45973 ( .A(n65134), .Z(n67345) );
  BUF_X1 U45974 ( .A(n65132), .Z(n67358) );
  BUF_X1 U45975 ( .A(n65134), .Z(n67346) );
  BUF_X1 U45976 ( .A(n65132), .Z(n67359) );
  BUF_X1 U45977 ( .A(n65134), .Z(n67347) );
  BUF_X1 U45978 ( .A(n65132), .Z(n67360) );
  BUF_X1 U45979 ( .A(n65134), .Z(n67348) );
  BUF_X1 U45980 ( .A(n65144), .Z(n67290) );
  BUF_X1 U45981 ( .A(n65149), .Z(n67266) );
  BUF_X1 U45982 ( .A(n65144), .Z(n67291) );
  BUF_X1 U45983 ( .A(n65149), .Z(n67267) );
  BUF_X1 U45984 ( .A(n65144), .Z(n67292) );
  BUF_X1 U45985 ( .A(n65149), .Z(n67268) );
  BUF_X1 U45986 ( .A(n65144), .Z(n67293) );
  BUF_X1 U45987 ( .A(n65149), .Z(n67269) );
  BUF_X1 U45988 ( .A(n65144), .Z(n67294) );
  BUF_X1 U45989 ( .A(n65149), .Z(n67270) );
  BUF_X1 U45990 ( .A(n63805), .Z(n67530) );
  BUF_X1 U45991 ( .A(n63801), .Z(n67554) );
  BUF_X1 U45992 ( .A(n63803), .Z(n67542) );
  BUF_X1 U45993 ( .A(n63805), .Z(n67531) );
  BUF_X1 U45994 ( .A(n63801), .Z(n67555) );
  BUF_X1 U45995 ( .A(n63803), .Z(n67543) );
  BUF_X1 U45996 ( .A(n63805), .Z(n67532) );
  BUF_X1 U45997 ( .A(n63801), .Z(n67556) );
  BUF_X1 U45998 ( .A(n63803), .Z(n67544) );
  BUF_X1 U45999 ( .A(n63805), .Z(n67533) );
  BUF_X1 U46000 ( .A(n63801), .Z(n67557) );
  BUF_X1 U46001 ( .A(n63803), .Z(n67545) );
  BUF_X1 U46002 ( .A(n63805), .Z(n67534) );
  BUF_X1 U46003 ( .A(n63801), .Z(n67558) );
  BUF_X1 U46004 ( .A(n63803), .Z(n67546) );
  BUF_X1 U46005 ( .A(n63818), .Z(n67464) );
  BUF_X1 U46006 ( .A(n63818), .Z(n67465) );
  BUF_X1 U46007 ( .A(n63818), .Z(n67466) );
  BUF_X1 U46008 ( .A(n63818), .Z(n67467) );
  BUF_X1 U46009 ( .A(n63818), .Z(n67468) );
  BUF_X1 U46010 ( .A(n65136), .Z(n67332) );
  BUF_X1 U46011 ( .A(n65136), .Z(n67333) );
  BUF_X1 U46012 ( .A(n65136), .Z(n67334) );
  BUF_X1 U46013 ( .A(n65136), .Z(n67335) );
  BUF_X1 U46014 ( .A(n65136), .Z(n67336) );
  BUF_X1 U46015 ( .A(n63813), .Z(n67488) );
  BUF_X1 U46016 ( .A(n63813), .Z(n67489) );
  BUF_X1 U46017 ( .A(n63813), .Z(n67490) );
  BUF_X1 U46018 ( .A(n63813), .Z(n67491) );
  BUF_X1 U46019 ( .A(n63813), .Z(n67492) );
  NAND2_X1 U46020 ( .A1(n68054), .A2(n67803), .ZN(n63163) );
  NAND2_X1 U46021 ( .A1(n68054), .A2(n67827), .ZN(n63094) );
  NAND2_X1 U46022 ( .A1(n68054), .A2(n67778), .ZN(n63231) );
  NAND2_X1 U46023 ( .A1(n68054), .A2(n67789), .ZN(n63228) );
  NAND2_X1 U46024 ( .A1(n68056), .A2(n67943), .ZN(n62628) );
  NAND2_X1 U46025 ( .A1(n68056), .A2(n67956), .ZN(n62561) );
  NAND2_X1 U46026 ( .A1(n68056), .A2(n68008), .ZN(n62292) );
  NAND2_X1 U46027 ( .A1(n68056), .A2(n67969), .ZN(n62495) );
  NAND2_X1 U46028 ( .A1(n68055), .A2(n67854), .ZN(n62961) );
  NAND2_X1 U46029 ( .A1(n68055), .A2(n67841), .ZN(n63028) );
  NAND2_X1 U46030 ( .A1(n68055), .A2(n67752), .ZN(n63364) );
  NAND2_X1 U46031 ( .A1(n68056), .A2(n67739), .ZN(n63431) );
  NAND2_X1 U46032 ( .A1(n68055), .A2(n67725), .ZN(n63499) );
  NAND2_X1 U46033 ( .A1(n68055), .A2(n67904), .ZN(n62763) );
  NAND2_X1 U46034 ( .A1(n68055), .A2(n67880), .ZN(n62828) );
  NAND2_X1 U46035 ( .A1(n68056), .A2(n68021), .ZN(n62226) );
  NAND2_X1 U46036 ( .A1(n68056), .A2(n67995), .ZN(n62359) );
  NAND2_X1 U46037 ( .A1(n68055), .A2(n67816), .ZN(n63097) );
  NAND2_X1 U46038 ( .A1(n68056), .A2(n67688), .ZN(n63634) );
  NAND2_X1 U46039 ( .A1(n68056), .A2(n67675), .ZN(n63700) );
  NAND2_X1 U46040 ( .A1(n68055), .A2(n67929), .ZN(n62695) );
  NAND2_X1 U46041 ( .A1(n68056), .A2(n67982), .ZN(n62425) );
  NAND2_X1 U46042 ( .A1(n68055), .A2(n67765), .ZN(n63298) );
  NAND2_X1 U46043 ( .A1(n68056), .A2(n67714), .ZN(n63502) );
  NAND2_X1 U46044 ( .A1(n68056), .A2(n67701), .ZN(n63568) );
  NAND2_X1 U46045 ( .A1(n68055), .A2(n67867), .ZN(n62894) );
  NAND2_X1 U46046 ( .A1(n68055), .A2(n67893), .ZN(n62765) );
  NAND2_X1 U46047 ( .A1(n68055), .A2(n67918), .ZN(n62698) );
  BUF_X1 U46048 ( .A(n65145), .Z(n67284) );
  BUF_X1 U46049 ( .A(n65133), .Z(n67350) );
  BUF_X1 U46050 ( .A(n65150), .Z(n67260) );
  BUF_X1 U46051 ( .A(n65145), .Z(n67285) );
  BUF_X1 U46052 ( .A(n65133), .Z(n67351) );
  BUF_X1 U46053 ( .A(n65150), .Z(n67261) );
  BUF_X1 U46054 ( .A(n65145), .Z(n67286) );
  BUF_X1 U46055 ( .A(n65133), .Z(n67352) );
  BUF_X1 U46056 ( .A(n65150), .Z(n67262) );
  BUF_X1 U46057 ( .A(n65145), .Z(n67287) );
  BUF_X1 U46058 ( .A(n65133), .Z(n67353) );
  BUF_X1 U46059 ( .A(n65150), .Z(n67263) );
  BUF_X1 U46060 ( .A(n65145), .Z(n67288) );
  BUF_X1 U46061 ( .A(n65133), .Z(n67354) );
  BUF_X1 U46062 ( .A(n65150), .Z(n67264) );
  BUF_X1 U46063 ( .A(n65135), .Z(n67338) );
  BUF_X1 U46064 ( .A(n65135), .Z(n67339) );
  BUF_X1 U46065 ( .A(n65135), .Z(n67340) );
  BUF_X1 U46066 ( .A(n65135), .Z(n67341) );
  BUF_X1 U46067 ( .A(n65135), .Z(n67342) );
  BUF_X1 U46068 ( .A(n63806), .Z(n67524) );
  BUF_X1 U46069 ( .A(n63814), .Z(n67482) );
  BUF_X1 U46070 ( .A(n63806), .Z(n67525) );
  BUF_X1 U46071 ( .A(n63814), .Z(n67483) );
  BUF_X1 U46072 ( .A(n63806), .Z(n67526) );
  BUF_X1 U46073 ( .A(n63814), .Z(n67484) );
  BUF_X1 U46074 ( .A(n63806), .Z(n67527) );
  BUF_X1 U46075 ( .A(n63814), .Z(n67485) );
  BUF_X1 U46076 ( .A(n63806), .Z(n67528) );
  BUF_X1 U46077 ( .A(n63814), .Z(n67486) );
  BUF_X1 U46078 ( .A(n63819), .Z(n67458) );
  BUF_X1 U46079 ( .A(n63819), .Z(n67459) );
  BUF_X1 U46080 ( .A(n63819), .Z(n67460) );
  BUF_X1 U46081 ( .A(n63819), .Z(n67461) );
  BUF_X1 U46082 ( .A(n63819), .Z(n67462) );
  BUF_X1 U46083 ( .A(n65137), .Z(n67326) );
  BUF_X1 U46084 ( .A(n65137), .Z(n67327) );
  BUF_X1 U46085 ( .A(n65137), .Z(n67328) );
  BUF_X1 U46086 ( .A(n65137), .Z(n67329) );
  BUF_X1 U46087 ( .A(n65137), .Z(n67330) );
  BUF_X1 U46088 ( .A(n63802), .Z(n67548) );
  BUF_X1 U46089 ( .A(n63804), .Z(n67536) );
  BUF_X1 U46090 ( .A(n63802), .Z(n67549) );
  BUF_X1 U46091 ( .A(n63804), .Z(n67537) );
  BUF_X1 U46092 ( .A(n63802), .Z(n67550) );
  BUF_X1 U46093 ( .A(n63804), .Z(n67538) );
  BUF_X1 U46094 ( .A(n63802), .Z(n67551) );
  BUF_X1 U46095 ( .A(n63804), .Z(n67539) );
  BUF_X1 U46096 ( .A(n63802), .Z(n67552) );
  BUF_X1 U46097 ( .A(n63804), .Z(n67540) );
  BUF_X1 U46098 ( .A(n65114), .Z(n67422) );
  BUF_X1 U46099 ( .A(n65114), .Z(n67423) );
  BUF_X1 U46100 ( .A(n65114), .Z(n67424) );
  BUF_X1 U46101 ( .A(n65114), .Z(n67425) );
  BUF_X1 U46102 ( .A(n65114), .Z(n67426) );
  BUF_X1 U46103 ( .A(n65119), .Z(n67398) );
  BUF_X1 U46104 ( .A(n65119), .Z(n67399) );
  BUF_X1 U46105 ( .A(n65119), .Z(n67400) );
  BUF_X1 U46106 ( .A(n65119), .Z(n67401) );
  BUF_X1 U46107 ( .A(n65119), .Z(n67402) );
  BUF_X1 U46108 ( .A(n63792), .Z(n67572) );
  BUF_X1 U46109 ( .A(n63792), .Z(n67573) );
  BUF_X1 U46110 ( .A(n63792), .Z(n67574) );
  BUF_X1 U46111 ( .A(n63792), .Z(n67575) );
  BUF_X1 U46112 ( .A(n63792), .Z(n67576) );
  BUF_X1 U46113 ( .A(n63786), .Z(n67596) );
  BUF_X1 U46114 ( .A(n63786), .Z(n67597) );
  BUF_X1 U46115 ( .A(n63786), .Z(n67598) );
  BUF_X1 U46116 ( .A(n63786), .Z(n67599) );
  BUF_X1 U46117 ( .A(n63786), .Z(n67600) );
  BUF_X1 U46118 ( .A(n65109), .Z(n67446) );
  BUF_X1 U46119 ( .A(n65124), .Z(n67374) );
  BUF_X1 U46120 ( .A(n65109), .Z(n67447) );
  BUF_X1 U46121 ( .A(n65124), .Z(n67375) );
  BUF_X1 U46122 ( .A(n65109), .Z(n67448) );
  BUF_X1 U46123 ( .A(n65124), .Z(n67376) );
  BUF_X1 U46124 ( .A(n65109), .Z(n67449) );
  BUF_X1 U46125 ( .A(n65124), .Z(n67377) );
  BUF_X1 U46126 ( .A(n65109), .Z(n67450) );
  BUF_X1 U46127 ( .A(n65124), .Z(n67378) );
  BUF_X1 U46128 ( .A(n63776), .Z(n67642) );
  BUF_X1 U46129 ( .A(n63781), .Z(n67620) );
  BUF_X1 U46130 ( .A(n63776), .Z(n67643) );
  BUF_X1 U46131 ( .A(n63781), .Z(n67621) );
  BUF_X1 U46132 ( .A(n63776), .Z(n67644) );
  BUF_X1 U46133 ( .A(n63781), .Z(n67622) );
  BUF_X1 U46134 ( .A(n63776), .Z(n67645) );
  BUF_X1 U46135 ( .A(n63781), .Z(n67623) );
  BUF_X1 U46136 ( .A(n63776), .Z(n67646) );
  BUF_X1 U46137 ( .A(n63781), .Z(n67624) );
  BUF_X1 U46138 ( .A(n65113), .Z(n67428) );
  BUF_X1 U46139 ( .A(n65108), .Z(n67452) );
  BUF_X1 U46140 ( .A(n63775), .Z(n67648) );
  BUF_X1 U46141 ( .A(n65118), .Z(n67404) );
  BUF_X1 U46142 ( .A(n65123), .Z(n67380) );
  BUF_X1 U46143 ( .A(n63791), .Z(n67578) );
  BUF_X1 U46144 ( .A(n63785), .Z(n67602) );
  BUF_X1 U46145 ( .A(n63780), .Z(n67626) );
  NAND2_X1 U46146 ( .A1(n68057), .A2(n68258), .ZN(n61959) );
  OAI21_X1 U46147 ( .B1(n62088), .B2(n62089), .A(n68052), .ZN(n61957) );
  OAI21_X1 U46148 ( .B1(n62089), .B2(n63025), .A(n68053), .ZN(n62959) );
  AND2_X1 U46149 ( .A1(n66276), .A2(n66277), .ZN(n65111) );
  BUF_X1 U46150 ( .A(n62493), .Z(n67967) );
  BUF_X1 U46151 ( .A(n62224), .Z(n68019) );
  BUF_X1 U46152 ( .A(n62357), .Z(n67993) );
  BUF_X1 U46153 ( .A(n62290), .Z(n68006) );
  BUF_X1 U46154 ( .A(n62157), .Z(n68032) );
  BUF_X1 U46155 ( .A(n62423), .Z(n67980) );
  BUF_X1 U46156 ( .A(n62626), .Z(n67941) );
  BUF_X1 U46157 ( .A(n62559), .Z(n67954) );
  BUF_X1 U46158 ( .A(n63161), .Z(n67801) );
  BUF_X1 U46159 ( .A(n63026), .Z(n67839) );
  BUF_X1 U46160 ( .A(n63362), .Z(n67750) );
  BUF_X1 U46161 ( .A(n63429), .Z(n67737) );
  BUF_X1 U46162 ( .A(n63764), .Z(n67660) );
  BUF_X1 U46163 ( .A(n62826), .Z(n67878) );
  BUF_X1 U46164 ( .A(n63095), .Z(n67814) );
  BUF_X1 U46165 ( .A(n63632), .Z(n67686) );
  BUF_X1 U46166 ( .A(n63698), .Z(n67673) );
  BUF_X1 U46167 ( .A(n63229), .Z(n67776) );
  BUF_X1 U46168 ( .A(n63296), .Z(n67763) );
  BUF_X1 U46169 ( .A(n63500), .Z(n67712) );
  BUF_X1 U46170 ( .A(n63566), .Z(n67699) );
  BUF_X1 U46171 ( .A(n62892), .Z(n67865) );
  BUF_X1 U46172 ( .A(n62764), .Z(n67891) );
  BUF_X1 U46173 ( .A(n62696), .Z(n67916) );
  BUF_X1 U46174 ( .A(n62090), .Z(n68045) );
  BUF_X1 U46175 ( .A(n62493), .Z(n67968) );
  BUF_X1 U46176 ( .A(n62224), .Z(n68020) );
  BUF_X1 U46177 ( .A(n62357), .Z(n67994) );
  BUF_X1 U46178 ( .A(n62290), .Z(n68007) );
  BUF_X1 U46179 ( .A(n62157), .Z(n68033) );
  BUF_X1 U46180 ( .A(n62423), .Z(n67981) );
  BUF_X1 U46181 ( .A(n62626), .Z(n67942) );
  BUF_X1 U46182 ( .A(n62559), .Z(n67955) );
  BUF_X1 U46183 ( .A(n63161), .Z(n67802) );
  BUF_X1 U46184 ( .A(n63026), .Z(n67840) );
  BUF_X1 U46185 ( .A(n63362), .Z(n67751) );
  BUF_X1 U46186 ( .A(n63429), .Z(n67738) );
  BUF_X1 U46187 ( .A(n63764), .Z(n67661) );
  BUF_X1 U46188 ( .A(n62826), .Z(n67879) );
  BUF_X1 U46189 ( .A(n63095), .Z(n67815) );
  BUF_X1 U46190 ( .A(n63632), .Z(n67687) );
  BUF_X1 U46191 ( .A(n63698), .Z(n67674) );
  BUF_X1 U46192 ( .A(n63229), .Z(n67777) );
  BUF_X1 U46193 ( .A(n63296), .Z(n67764) );
  BUF_X1 U46194 ( .A(n63500), .Z(n67713) );
  BUF_X1 U46195 ( .A(n63566), .Z(n67700) );
  BUF_X1 U46196 ( .A(n62892), .Z(n67866) );
  BUF_X1 U46197 ( .A(n62764), .Z(n67892) );
  BUF_X1 U46198 ( .A(n62696), .Z(n67917) );
  BUF_X1 U46199 ( .A(n62090), .Z(n68046) );
  NOR3_X1 U46200 ( .A1(n66301), .A2(n67434), .A3(n66299), .ZN(n66277) );
  NOR3_X1 U46201 ( .A1(n66291), .A2(n66297), .A3(n66292), .ZN(n66276) );
  OAI21_X1 U46202 ( .B1(n62223), .B2(n63428), .A(n68054), .ZN(n63498) );
  OAI21_X1 U46203 ( .B1(n62356), .B2(n62625), .A(n68053), .ZN(n62762) );
  OAI21_X1 U46204 ( .B1(n62223), .B2(n62625), .A(n68052), .ZN(n62693) );
  OAI21_X1 U46205 ( .B1(n62223), .B2(n63025), .A(n68053), .ZN(n63093) );
  OAI21_X1 U46206 ( .B1(n62356), .B2(n63092), .A(n68053), .ZN(n63227) );
  BUF_X1 U46207 ( .A(n65112), .Z(n67434) );
  BUF_X1 U46208 ( .A(n65112), .Z(n67435) );
  BUF_X1 U46209 ( .A(n65112), .Z(n67436) );
  BUF_X1 U46210 ( .A(n65112), .Z(n67437) );
  NOR3_X1 U46211 ( .A1(n65095), .A2(n65094), .A3(n65093), .ZN(n65085) );
  OAI222_X1 U46212 ( .A1(n62891), .A2(n67320), .B1(n63160), .B2(n67314), .C1(
        n62355), .C2(n67308), .ZN(n66293) );
  OAI222_X1 U46213 ( .A1(n62890), .A2(n67320), .B1(n63159), .B2(n67314), .C1(
        n62354), .C2(n67308), .ZN(n66261) );
  OAI222_X1 U46214 ( .A1(n62889), .A2(n67320), .B1(n63158), .B2(n67314), .C1(
        n62353), .C2(n67308), .ZN(n66243) );
  OAI222_X1 U46215 ( .A1(n62888), .A2(n67320), .B1(n63157), .B2(n67314), .C1(
        n62352), .C2(n67308), .ZN(n66225) );
  OAI222_X1 U46216 ( .A1(n62887), .A2(n67320), .B1(n63156), .B2(n67314), .C1(
        n62351), .C2(n67308), .ZN(n66207) );
  OAI222_X1 U46217 ( .A1(n62886), .A2(n67320), .B1(n63155), .B2(n67314), .C1(
        n62350), .C2(n67308), .ZN(n66189) );
  OAI222_X1 U46218 ( .A1(n62885), .A2(n67320), .B1(n63154), .B2(n67314), .C1(
        n62349), .C2(n67308), .ZN(n66171) );
  OAI222_X1 U46219 ( .A1(n62884), .A2(n67320), .B1(n63153), .B2(n67314), .C1(
        n62348), .C2(n67308), .ZN(n66153) );
  OAI222_X1 U46220 ( .A1(n62883), .A2(n67320), .B1(n63152), .B2(n67314), .C1(
        n62347), .C2(n67308), .ZN(n66135) );
  OAI222_X1 U46221 ( .A1(n62882), .A2(n67320), .B1(n63151), .B2(n67314), .C1(
        n62346), .C2(n67308), .ZN(n66117) );
  OAI222_X1 U46222 ( .A1(n62881), .A2(n67320), .B1(n63150), .B2(n67314), .C1(
        n62345), .C2(n67308), .ZN(n66099) );
  OAI222_X1 U46223 ( .A1(n62880), .A2(n67320), .B1(n63149), .B2(n67314), .C1(
        n62344), .C2(n67308), .ZN(n66081) );
  OAI222_X1 U46224 ( .A1(n62879), .A2(n67321), .B1(n63148), .B2(n67315), .C1(
        n62343), .C2(n67309), .ZN(n66063) );
  OAI222_X1 U46225 ( .A1(n62878), .A2(n67321), .B1(n63147), .B2(n67315), .C1(
        n62342), .C2(n67309), .ZN(n66045) );
  OAI222_X1 U46226 ( .A1(n62877), .A2(n67321), .B1(n63146), .B2(n67315), .C1(
        n62341), .C2(n67309), .ZN(n66027) );
  OAI222_X1 U46227 ( .A1(n62876), .A2(n67321), .B1(n63145), .B2(n67315), .C1(
        n62340), .C2(n67309), .ZN(n66009) );
  OAI222_X1 U46228 ( .A1(n62875), .A2(n67321), .B1(n63144), .B2(n67315), .C1(
        n62339), .C2(n67309), .ZN(n65991) );
  OAI222_X1 U46229 ( .A1(n62874), .A2(n67321), .B1(n63143), .B2(n67315), .C1(
        n62338), .C2(n67309), .ZN(n65973) );
  OAI222_X1 U46230 ( .A1(n62873), .A2(n67321), .B1(n63142), .B2(n67315), .C1(
        n62337), .C2(n67309), .ZN(n65955) );
  OAI222_X1 U46231 ( .A1(n62872), .A2(n67321), .B1(n63141), .B2(n67315), .C1(
        n62336), .C2(n67309), .ZN(n65937) );
  OAI222_X1 U46232 ( .A1(n62871), .A2(n67321), .B1(n63140), .B2(n67315), .C1(
        n62335), .C2(n67309), .ZN(n65919) );
  OAI222_X1 U46233 ( .A1(n62870), .A2(n67321), .B1(n63139), .B2(n67315), .C1(
        n62334), .C2(n67309), .ZN(n65901) );
  OAI222_X1 U46234 ( .A1(n62869), .A2(n67321), .B1(n63138), .B2(n67315), .C1(
        n62333), .C2(n67309), .ZN(n65883) );
  OAI222_X1 U46235 ( .A1(n62868), .A2(n67321), .B1(n63137), .B2(n67315), .C1(
        n62332), .C2(n67309), .ZN(n65865) );
  OAI222_X1 U46236 ( .A1(n62867), .A2(n67322), .B1(n63136), .B2(n67316), .C1(
        n62331), .C2(n67310), .ZN(n65847) );
  OAI222_X1 U46237 ( .A1(n62866), .A2(n67322), .B1(n63135), .B2(n67316), .C1(
        n62330), .C2(n67310), .ZN(n65829) );
  OAI222_X1 U46238 ( .A1(n62865), .A2(n67322), .B1(n63134), .B2(n67316), .C1(
        n62329), .C2(n67310), .ZN(n65811) );
  OAI222_X1 U46239 ( .A1(n62864), .A2(n67322), .B1(n63133), .B2(n67316), .C1(
        n62328), .C2(n67310), .ZN(n65793) );
  OAI222_X1 U46240 ( .A1(n62863), .A2(n67322), .B1(n63132), .B2(n67316), .C1(
        n62327), .C2(n67310), .ZN(n65775) );
  OAI222_X1 U46241 ( .A1(n62862), .A2(n67322), .B1(n63131), .B2(n67316), .C1(
        n62326), .C2(n67310), .ZN(n65757) );
  OAI222_X1 U46242 ( .A1(n62861), .A2(n67322), .B1(n63130), .B2(n67316), .C1(
        n62325), .C2(n67310), .ZN(n65739) );
  OAI222_X1 U46243 ( .A1(n62860), .A2(n67322), .B1(n63129), .B2(n67316), .C1(
        n62324), .C2(n67310), .ZN(n65721) );
  OAI222_X1 U46244 ( .A1(n62859), .A2(n67322), .B1(n63128), .B2(n67316), .C1(
        n62323), .C2(n67310), .ZN(n65703) );
  OAI222_X1 U46245 ( .A1(n62858), .A2(n67322), .B1(n63127), .B2(n67316), .C1(
        n62322), .C2(n67310), .ZN(n65685) );
  OAI222_X1 U46246 ( .A1(n62857), .A2(n67322), .B1(n63126), .B2(n67316), .C1(
        n62321), .C2(n67310), .ZN(n65667) );
  OAI222_X1 U46247 ( .A1(n62856), .A2(n67322), .B1(n63125), .B2(n67316), .C1(
        n62320), .C2(n67310), .ZN(n65649) );
  OAI222_X1 U46248 ( .A1(n62855), .A2(n67323), .B1(n63124), .B2(n67317), .C1(
        n62319), .C2(n67311), .ZN(n65631) );
  OAI222_X1 U46249 ( .A1(n62854), .A2(n67323), .B1(n63123), .B2(n67317), .C1(
        n62318), .C2(n67311), .ZN(n65613) );
  OAI222_X1 U46250 ( .A1(n62853), .A2(n67323), .B1(n63122), .B2(n67317), .C1(
        n62317), .C2(n67311), .ZN(n65595) );
  OAI222_X1 U46251 ( .A1(n62852), .A2(n67323), .B1(n63121), .B2(n67317), .C1(
        n62316), .C2(n67311), .ZN(n65577) );
  OAI222_X1 U46252 ( .A1(n62851), .A2(n67323), .B1(n63120), .B2(n67317), .C1(
        n62315), .C2(n67311), .ZN(n65559) );
  OAI222_X1 U46253 ( .A1(n62850), .A2(n67323), .B1(n63119), .B2(n67317), .C1(
        n62314), .C2(n67311), .ZN(n65541) );
  OAI222_X1 U46254 ( .A1(n62849), .A2(n67323), .B1(n63118), .B2(n67317), .C1(
        n62313), .C2(n67311), .ZN(n65523) );
  OAI222_X1 U46255 ( .A1(n62848), .A2(n67323), .B1(n63117), .B2(n67317), .C1(
        n62312), .C2(n67311), .ZN(n65505) );
  OAI222_X1 U46256 ( .A1(n62847), .A2(n67323), .B1(n63116), .B2(n67317), .C1(
        n62311), .C2(n67311), .ZN(n65487) );
  OAI222_X1 U46257 ( .A1(n62846), .A2(n67323), .B1(n63115), .B2(n67317), .C1(
        n62310), .C2(n67311), .ZN(n65469) );
  OAI222_X1 U46258 ( .A1(n62845), .A2(n67323), .B1(n63114), .B2(n67317), .C1(
        n62309), .C2(n67311), .ZN(n65451) );
  OAI222_X1 U46259 ( .A1(n62844), .A2(n67323), .B1(n63113), .B2(n67317), .C1(
        n62308), .C2(n67311), .ZN(n65433) );
  OAI222_X1 U46260 ( .A1(n62843), .A2(n67324), .B1(n63112), .B2(n67318), .C1(
        n62307), .C2(n67312), .ZN(n65415) );
  OAI222_X1 U46261 ( .A1(n62842), .A2(n67324), .B1(n63111), .B2(n67318), .C1(
        n62306), .C2(n67312), .ZN(n65397) );
  OAI222_X1 U46262 ( .A1(n62841), .A2(n67324), .B1(n63110), .B2(n67318), .C1(
        n62305), .C2(n67312), .ZN(n65379) );
  OAI222_X1 U46263 ( .A1(n62840), .A2(n67324), .B1(n63109), .B2(n67318), .C1(
        n62304), .C2(n67312), .ZN(n65361) );
  OAI222_X1 U46264 ( .A1(n62839), .A2(n67324), .B1(n63108), .B2(n67318), .C1(
        n62303), .C2(n67312), .ZN(n65343) );
  OAI222_X1 U46265 ( .A1(n62838), .A2(n67324), .B1(n63107), .B2(n67318), .C1(
        n62302), .C2(n67312), .ZN(n65325) );
  OAI222_X1 U46266 ( .A1(n62837), .A2(n67324), .B1(n63106), .B2(n67318), .C1(
        n62301), .C2(n67312), .ZN(n65307) );
  OAI222_X1 U46267 ( .A1(n62836), .A2(n67324), .B1(n63105), .B2(n67318), .C1(
        n62300), .C2(n67312), .ZN(n65289) );
  OAI222_X1 U46268 ( .A1(n62835), .A2(n67324), .B1(n63104), .B2(n67318), .C1(
        n62299), .C2(n67312), .ZN(n65271) );
  OAI222_X1 U46269 ( .A1(n62834), .A2(n67324), .B1(n63103), .B2(n67318), .C1(
        n62298), .C2(n67312), .ZN(n65253) );
  OAI222_X1 U46270 ( .A1(n62833), .A2(n67324), .B1(n63102), .B2(n67318), .C1(
        n62297), .C2(n67312), .ZN(n65235) );
  OAI222_X1 U46271 ( .A1(n62832), .A2(n67324), .B1(n63101), .B2(n67318), .C1(
        n62296), .C2(n67312), .ZN(n65217) );
  OAI222_X1 U46272 ( .A1(n63226), .A2(n67518), .B1(n62155), .B2(n67512), .C1(
        n62558), .C2(n67506), .ZN(n65089) );
  OAI222_X1 U46273 ( .A1(n63225), .A2(n67518), .B1(n62154), .B2(n67512), .C1(
        n62557), .C2(n67506), .ZN(n65057) );
  OAI222_X1 U46274 ( .A1(n63224), .A2(n67518), .B1(n62153), .B2(n67512), .C1(
        n62556), .C2(n67506), .ZN(n65037) );
  OAI222_X1 U46275 ( .A1(n63223), .A2(n67518), .B1(n62152), .B2(n67512), .C1(
        n62555), .C2(n67506), .ZN(n65017) );
  OAI222_X1 U46276 ( .A1(n63222), .A2(n67518), .B1(n62151), .B2(n67512), .C1(
        n62554), .C2(n67506), .ZN(n64997) );
  OAI222_X1 U46277 ( .A1(n63221), .A2(n67518), .B1(n62150), .B2(n67512), .C1(
        n62553), .C2(n67506), .ZN(n64977) );
  OAI222_X1 U46278 ( .A1(n63220), .A2(n67518), .B1(n62149), .B2(n67512), .C1(
        n62552), .C2(n67506), .ZN(n64957) );
  OAI222_X1 U46279 ( .A1(n63219), .A2(n67518), .B1(n62148), .B2(n67512), .C1(
        n62551), .C2(n67506), .ZN(n64937) );
  OAI222_X1 U46280 ( .A1(n63218), .A2(n67518), .B1(n62147), .B2(n67512), .C1(
        n62550), .C2(n67506), .ZN(n64917) );
  OAI222_X1 U46281 ( .A1(n63217), .A2(n67518), .B1(n62146), .B2(n67512), .C1(
        n62549), .C2(n67506), .ZN(n64897) );
  OAI222_X1 U46282 ( .A1(n63216), .A2(n67518), .B1(n62145), .B2(n67512), .C1(
        n62548), .C2(n67506), .ZN(n64877) );
  OAI222_X1 U46283 ( .A1(n63215), .A2(n67518), .B1(n62144), .B2(n67512), .C1(
        n62547), .C2(n67506), .ZN(n64857) );
  OAI222_X1 U46284 ( .A1(n63214), .A2(n67519), .B1(n62143), .B2(n67513), .C1(
        n62546), .C2(n67507), .ZN(n64837) );
  OAI222_X1 U46285 ( .A1(n63213), .A2(n67519), .B1(n62142), .B2(n67513), .C1(
        n62545), .C2(n67507), .ZN(n64817) );
  OAI222_X1 U46286 ( .A1(n63212), .A2(n67519), .B1(n62141), .B2(n67513), .C1(
        n62544), .C2(n67507), .ZN(n64797) );
  OAI222_X1 U46287 ( .A1(n63211), .A2(n67519), .B1(n62140), .B2(n67513), .C1(
        n62543), .C2(n67507), .ZN(n64777) );
  OAI222_X1 U46288 ( .A1(n63210), .A2(n67519), .B1(n62139), .B2(n67513), .C1(
        n62542), .C2(n67507), .ZN(n64757) );
  OAI222_X1 U46289 ( .A1(n63209), .A2(n67519), .B1(n62138), .B2(n67513), .C1(
        n62541), .C2(n67507), .ZN(n64737) );
  OAI222_X1 U46290 ( .A1(n63208), .A2(n67519), .B1(n62137), .B2(n67513), .C1(
        n62540), .C2(n67507), .ZN(n64717) );
  OAI222_X1 U46291 ( .A1(n63207), .A2(n67519), .B1(n62136), .B2(n67513), .C1(
        n62539), .C2(n67507), .ZN(n64697) );
  OAI222_X1 U46292 ( .A1(n63206), .A2(n67519), .B1(n62135), .B2(n67513), .C1(
        n62538), .C2(n67507), .ZN(n64677) );
  OAI222_X1 U46293 ( .A1(n63205), .A2(n67519), .B1(n62134), .B2(n67513), .C1(
        n62537), .C2(n67507), .ZN(n64657) );
  OAI222_X1 U46294 ( .A1(n63204), .A2(n67519), .B1(n62133), .B2(n67513), .C1(
        n62536), .C2(n67507), .ZN(n64637) );
  OAI222_X1 U46295 ( .A1(n63203), .A2(n67519), .B1(n62132), .B2(n67513), .C1(
        n62535), .C2(n67507), .ZN(n64617) );
  OAI222_X1 U46296 ( .A1(n63202), .A2(n67520), .B1(n62131), .B2(n67514), .C1(
        n62534), .C2(n67508), .ZN(n64597) );
  OAI222_X1 U46297 ( .A1(n63201), .A2(n67520), .B1(n62130), .B2(n67514), .C1(
        n62533), .C2(n67508), .ZN(n64577) );
  OAI222_X1 U46298 ( .A1(n63200), .A2(n67520), .B1(n62129), .B2(n67514), .C1(
        n62532), .C2(n67508), .ZN(n64557) );
  OAI222_X1 U46299 ( .A1(n63199), .A2(n67520), .B1(n62128), .B2(n67514), .C1(
        n62531), .C2(n67508), .ZN(n64537) );
  OAI222_X1 U46300 ( .A1(n63198), .A2(n67520), .B1(n62127), .B2(n67514), .C1(
        n62530), .C2(n67508), .ZN(n64517) );
  OAI222_X1 U46301 ( .A1(n63197), .A2(n67520), .B1(n62126), .B2(n67514), .C1(
        n62529), .C2(n67508), .ZN(n64497) );
  OAI222_X1 U46302 ( .A1(n63196), .A2(n67520), .B1(n62125), .B2(n67514), .C1(
        n62528), .C2(n67508), .ZN(n64477) );
  OAI222_X1 U46303 ( .A1(n63195), .A2(n67520), .B1(n62124), .B2(n67514), .C1(
        n62527), .C2(n67508), .ZN(n64457) );
  OAI222_X1 U46304 ( .A1(n63194), .A2(n67520), .B1(n62123), .B2(n67514), .C1(
        n62526), .C2(n67508), .ZN(n64437) );
  OAI222_X1 U46305 ( .A1(n63193), .A2(n67520), .B1(n62122), .B2(n67514), .C1(
        n62525), .C2(n67508), .ZN(n64417) );
  OAI222_X1 U46306 ( .A1(n63192), .A2(n67520), .B1(n62121), .B2(n67514), .C1(
        n62524), .C2(n67508), .ZN(n64397) );
  OAI222_X1 U46307 ( .A1(n63191), .A2(n67520), .B1(n62120), .B2(n67514), .C1(
        n62523), .C2(n67508), .ZN(n64377) );
  OAI222_X1 U46308 ( .A1(n63190), .A2(n67521), .B1(n62119), .B2(n67515), .C1(
        n62522), .C2(n67509), .ZN(n64357) );
  OAI222_X1 U46309 ( .A1(n63189), .A2(n67521), .B1(n62118), .B2(n67515), .C1(
        n62521), .C2(n67509), .ZN(n64337) );
  OAI222_X1 U46310 ( .A1(n63188), .A2(n67521), .B1(n62117), .B2(n67515), .C1(
        n62520), .C2(n67509), .ZN(n64317) );
  OAI222_X1 U46311 ( .A1(n63187), .A2(n67521), .B1(n62116), .B2(n67515), .C1(
        n62519), .C2(n67509), .ZN(n64297) );
  OAI222_X1 U46312 ( .A1(n63186), .A2(n67521), .B1(n62115), .B2(n67515), .C1(
        n62518), .C2(n67509), .ZN(n64277) );
  OAI222_X1 U46313 ( .A1(n63185), .A2(n67521), .B1(n62114), .B2(n67515), .C1(
        n62517), .C2(n67509), .ZN(n64257) );
  OAI222_X1 U46314 ( .A1(n63184), .A2(n67521), .B1(n62113), .B2(n67515), .C1(
        n62516), .C2(n67509), .ZN(n64237) );
  OAI222_X1 U46315 ( .A1(n63183), .A2(n67521), .B1(n62112), .B2(n67515), .C1(
        n62515), .C2(n67509), .ZN(n64217) );
  OAI222_X1 U46316 ( .A1(n63182), .A2(n67521), .B1(n62111), .B2(n67515), .C1(
        n62514), .C2(n67509), .ZN(n64197) );
  OAI222_X1 U46317 ( .A1(n63181), .A2(n67521), .B1(n62110), .B2(n67515), .C1(
        n62513), .C2(n67509), .ZN(n64177) );
  OAI222_X1 U46318 ( .A1(n63180), .A2(n67521), .B1(n62109), .B2(n67515), .C1(
        n62512), .C2(n67509), .ZN(n64157) );
  OAI222_X1 U46319 ( .A1(n63179), .A2(n67521), .B1(n62108), .B2(n67515), .C1(
        n62511), .C2(n67509), .ZN(n64137) );
  OAI222_X1 U46320 ( .A1(n63178), .A2(n67522), .B1(n62107), .B2(n67516), .C1(
        n62510), .C2(n67510), .ZN(n64117) );
  OAI222_X1 U46321 ( .A1(n63177), .A2(n67522), .B1(n62106), .B2(n67516), .C1(
        n62509), .C2(n67510), .ZN(n64097) );
  OAI222_X1 U46322 ( .A1(n63176), .A2(n67522), .B1(n62105), .B2(n67516), .C1(
        n62508), .C2(n67510), .ZN(n64077) );
  OAI222_X1 U46323 ( .A1(n63175), .A2(n67522), .B1(n62104), .B2(n67516), .C1(
        n62507), .C2(n67510), .ZN(n64057) );
  OAI222_X1 U46324 ( .A1(n63174), .A2(n67522), .B1(n62103), .B2(n67516), .C1(
        n62506), .C2(n67510), .ZN(n64037) );
  OAI222_X1 U46325 ( .A1(n63173), .A2(n67522), .B1(n62102), .B2(n67516), .C1(
        n62505), .C2(n67510), .ZN(n64017) );
  OAI222_X1 U46326 ( .A1(n63172), .A2(n67522), .B1(n62101), .B2(n67516), .C1(
        n62504), .C2(n67510), .ZN(n63997) );
  OAI222_X1 U46327 ( .A1(n63171), .A2(n67522), .B1(n62100), .B2(n67516), .C1(
        n62503), .C2(n67510), .ZN(n63977) );
  OAI222_X1 U46328 ( .A1(n63170), .A2(n67522), .B1(n62099), .B2(n67516), .C1(
        n62502), .C2(n67510), .ZN(n63957) );
  OAI222_X1 U46329 ( .A1(n63169), .A2(n67522), .B1(n62098), .B2(n67516), .C1(
        n62501), .C2(n67510), .ZN(n63937) );
  OAI222_X1 U46330 ( .A1(n63168), .A2(n67522), .B1(n62097), .B2(n67516), .C1(
        n62500), .C2(n67510), .ZN(n63917) );
  OAI222_X1 U46331 ( .A1(n63167), .A2(n67522), .B1(n62096), .B2(n67516), .C1(
        n62499), .C2(n67510), .ZN(n63897) );
  OAI222_X1 U46332 ( .A1(n62829), .A2(n67325), .B1(n63098), .B2(n67319), .C1(
        n62293), .C2(n67313), .ZN(n65163) );
  OAI222_X1 U46333 ( .A1(n62827), .A2(n67325), .B1(n63096), .B2(n67319), .C1(
        n62291), .C2(n67313), .ZN(n65128) );
  OAI222_X1 U46334 ( .A1(n62831), .A2(n67325), .B1(n63100), .B2(n67319), .C1(
        n62295), .C2(n67313), .ZN(n65199) );
  OAI222_X1 U46335 ( .A1(n62830), .A2(n67325), .B1(n63099), .B2(n67319), .C1(
        n62294), .C2(n67313), .ZN(n65181) );
  NAND2_X1 U46336 ( .A1(n65086), .A2(n65081), .ZN(n63804) );
  NAND2_X1 U46337 ( .A1(n66278), .A2(n66279), .ZN(n65109) );
  NAND2_X1 U46338 ( .A1(n66278), .A2(n66290), .ZN(n65124) );
  NAND2_X1 U46339 ( .A1(n66281), .A2(n66290), .ZN(n65137) );
  NAND2_X1 U46340 ( .A1(n66277), .A2(n66290), .ZN(n65136) );
  NAND2_X1 U46341 ( .A1(n63496), .A2(n63497), .ZN(n62089) );
  BUF_X1 U46342 ( .A(n62087), .Z(n68053) );
  BUF_X1 U46343 ( .A(n62087), .Z(n68052) );
  BUF_X1 U46344 ( .A(n62087), .Z(n68054) );
  BUF_X1 U46345 ( .A(n62087), .Z(n68056) );
  BUF_X1 U46346 ( .A(n62087), .Z(n68055) );
  NAND2_X1 U46347 ( .A1(n66283), .A2(n66290), .ZN(n65139) );
  NAND2_X1 U46348 ( .A1(n66287), .A2(n66283), .ZN(n65145) );
  NAND2_X1 U46349 ( .A1(n66285), .A2(n66283), .ZN(n65133) );
  NAND2_X1 U46350 ( .A1(n66279), .A2(n66283), .ZN(n65132) );
  NAND2_X1 U46351 ( .A1(n66289), .A2(n66283), .ZN(n65134) );
  NAND2_X1 U46352 ( .A1(n66286), .A2(n66283), .ZN(n65150) );
  NAND2_X1 U46353 ( .A1(n66276), .A2(n66283), .ZN(n65114) );
  NAND2_X1 U46354 ( .A1(n65073), .A2(n65078), .ZN(n63806) );
  NAND2_X1 U46355 ( .A1(n65076), .A2(n65078), .ZN(n63805) );
  NAND2_X1 U46356 ( .A1(n65080), .A2(n65078), .ZN(n63801) );
  NAND2_X1 U46357 ( .A1(n65082), .A2(n65086), .ZN(n63803) );
  NAND2_X1 U46358 ( .A1(n65077), .A2(n65086), .ZN(n63792) );
  NAND2_X1 U46359 ( .A1(n65085), .A2(n65086), .ZN(n63814) );
  NAND2_X1 U46360 ( .A1(n66276), .A2(n66278), .ZN(n65119) );
  NAND2_X1 U46361 ( .A1(n65078), .A2(n65081), .ZN(n63808) );
  OAI22_X1 U46362 ( .A1(n62699), .A2(n67349), .B1(n62895), .B2(n67343), .ZN(
        n65165) );
  OAI22_X1 U46363 ( .A1(n62697), .A2(n67349), .B1(n62893), .B2(n67343), .ZN(
        n65130) );
  OAI22_X1 U46364 ( .A1(n62701), .A2(n67349), .B1(n62897), .B2(n67343), .ZN(
        n65201) );
  OAI22_X1 U46365 ( .A1(n62700), .A2(n67349), .B1(n62896), .B2(n67343), .ZN(
        n65183) );
  OAI22_X1 U46366 ( .A1(n63432), .A2(n67271), .B1(n62227), .B2(n67265), .ZN(
        n65168) );
  OAI22_X1 U46367 ( .A1(n63430), .A2(n67271), .B1(n62225), .B2(n67265), .ZN(
        n65148) );
  OAI22_X1 U46368 ( .A1(n63434), .A2(n67271), .B1(n62229), .B2(n67265), .ZN(
        n65204) );
  OAI22_X1 U46369 ( .A1(n63433), .A2(n67271), .B1(n62228), .B2(n67265), .ZN(
        n65186) );
  OAI22_X1 U46370 ( .A1(n63301), .A2(n67493), .B1(n63637), .B2(n67487), .ZN(
        n63881) );
  OAI22_X1 U46371 ( .A1(n62701), .A2(n67469), .B1(n62162), .B2(n67463), .ZN(
        n63882) );
  OAI22_X1 U46372 ( .A1(n63300), .A2(n67493), .B1(n63636), .B2(n67487), .ZN(
        n63860) );
  OAI22_X1 U46373 ( .A1(n62700), .A2(n67469), .B1(n62161), .B2(n67463), .ZN(
        n63861) );
  OAI22_X1 U46374 ( .A1(n63299), .A2(n67493), .B1(n63635), .B2(n67487), .ZN(
        n63839) );
  OAI22_X1 U46375 ( .A1(n62699), .A2(n67469), .B1(n62160), .B2(n67463), .ZN(
        n63840) );
  OAI22_X1 U46376 ( .A1(n63297), .A2(n67493), .B1(n63633), .B2(n67487), .ZN(
        n63812) );
  OAI22_X1 U46377 ( .A1(n62697), .A2(n67469), .B1(n62158), .B2(n67463), .ZN(
        n63817) );
  OAI22_X1 U46378 ( .A1(n63299), .A2(n67337), .B1(n63029), .B2(n67331), .ZN(
        n65164) );
  OAI22_X1 U46379 ( .A1(n63297), .A2(n67337), .B1(n63027), .B2(n67331), .ZN(
        n65129) );
  OAI22_X1 U46380 ( .A1(n63301), .A2(n67337), .B1(n63031), .B2(n67331), .ZN(
        n65200) );
  OAI22_X1 U46381 ( .A1(n63300), .A2(n67337), .B1(n63030), .B2(n67331), .ZN(
        n65182) );
  OAI22_X1 U46382 ( .A1(n62964), .A2(n67535), .B1(n62564), .B2(n67529), .ZN(
        n63878) );
  OAI22_X1 U46383 ( .A1(n62963), .A2(n67535), .B1(n62563), .B2(n67529), .ZN(
        n63857) );
  OAI22_X1 U46384 ( .A1(n62962), .A2(n67535), .B1(n62562), .B2(n67529), .ZN(
        n63836) );
  OAI22_X1 U46385 ( .A1(n62960), .A2(n67535), .B1(n62560), .B2(n67529), .ZN(
        n63798) );
  NAND2_X1 U46386 ( .A1(n66286), .A2(n66281), .ZN(n65144) );
  NAND2_X1 U46387 ( .A1(n66276), .A2(n66281), .ZN(n65149) );
  NAND2_X1 U46388 ( .A1(n66278), .A2(n66287), .ZN(n65140) );
  NAND2_X1 U46389 ( .A1(n66289), .A2(n66277), .ZN(n65135) );
  OAI22_X1 U46390 ( .A1(n62761), .A2(n67344), .B1(n62957), .B2(n67338), .ZN(
        n66295) );
  OAI22_X1 U46391 ( .A1(n62760), .A2(n67344), .B1(n62956), .B2(n67338), .ZN(
        n66263) );
  OAI22_X1 U46392 ( .A1(n62759), .A2(n67344), .B1(n62955), .B2(n67338), .ZN(
        n66245) );
  OAI22_X1 U46393 ( .A1(n62758), .A2(n67344), .B1(n62954), .B2(n67338), .ZN(
        n66227) );
  OAI22_X1 U46394 ( .A1(n62757), .A2(n67344), .B1(n62953), .B2(n67338), .ZN(
        n66209) );
  OAI22_X1 U46395 ( .A1(n62756), .A2(n67344), .B1(n62952), .B2(n67338), .ZN(
        n66191) );
  OAI22_X1 U46396 ( .A1(n62755), .A2(n67344), .B1(n62951), .B2(n67338), .ZN(
        n66173) );
  OAI22_X1 U46397 ( .A1(n62754), .A2(n67344), .B1(n62950), .B2(n67338), .ZN(
        n66155) );
  OAI22_X1 U46398 ( .A1(n62753), .A2(n67344), .B1(n62949), .B2(n67338), .ZN(
        n66137) );
  OAI22_X1 U46399 ( .A1(n62752), .A2(n67344), .B1(n62948), .B2(n67338), .ZN(
        n66119) );
  OAI22_X1 U46400 ( .A1(n62751), .A2(n67344), .B1(n62947), .B2(n67338), .ZN(
        n66101) );
  OAI22_X1 U46401 ( .A1(n62750), .A2(n67344), .B1(n62946), .B2(n67338), .ZN(
        n66083) );
  OAI22_X1 U46402 ( .A1(n62749), .A2(n67345), .B1(n62945), .B2(n67339), .ZN(
        n66065) );
  OAI22_X1 U46403 ( .A1(n62748), .A2(n67345), .B1(n62944), .B2(n67339), .ZN(
        n66047) );
  OAI22_X1 U46404 ( .A1(n62747), .A2(n67345), .B1(n62943), .B2(n67339), .ZN(
        n66029) );
  OAI22_X1 U46405 ( .A1(n62746), .A2(n67345), .B1(n62942), .B2(n67339), .ZN(
        n66011) );
  OAI22_X1 U46406 ( .A1(n62745), .A2(n67345), .B1(n62941), .B2(n67339), .ZN(
        n65993) );
  OAI22_X1 U46407 ( .A1(n62744), .A2(n67345), .B1(n62940), .B2(n67339), .ZN(
        n65975) );
  OAI22_X1 U46408 ( .A1(n62743), .A2(n67345), .B1(n62939), .B2(n67339), .ZN(
        n65957) );
  OAI22_X1 U46409 ( .A1(n62742), .A2(n67345), .B1(n62938), .B2(n67339), .ZN(
        n65939) );
  OAI22_X1 U46410 ( .A1(n62741), .A2(n67345), .B1(n62937), .B2(n67339), .ZN(
        n65921) );
  OAI22_X1 U46411 ( .A1(n62740), .A2(n67345), .B1(n62936), .B2(n67339), .ZN(
        n65903) );
  OAI22_X1 U46412 ( .A1(n62739), .A2(n67345), .B1(n62935), .B2(n67339), .ZN(
        n65885) );
  OAI22_X1 U46413 ( .A1(n62738), .A2(n67345), .B1(n62934), .B2(n67339), .ZN(
        n65867) );
  OAI22_X1 U46414 ( .A1(n62737), .A2(n67346), .B1(n62933), .B2(n67340), .ZN(
        n65849) );
  OAI22_X1 U46415 ( .A1(n62736), .A2(n67346), .B1(n62932), .B2(n67340), .ZN(
        n65831) );
  OAI22_X1 U46416 ( .A1(n62735), .A2(n67346), .B1(n62931), .B2(n67340), .ZN(
        n65813) );
  OAI22_X1 U46417 ( .A1(n62734), .A2(n67346), .B1(n62930), .B2(n67340), .ZN(
        n65795) );
  OAI22_X1 U46418 ( .A1(n62733), .A2(n67346), .B1(n62929), .B2(n67340), .ZN(
        n65777) );
  OAI22_X1 U46419 ( .A1(n62732), .A2(n67346), .B1(n62928), .B2(n67340), .ZN(
        n65759) );
  OAI22_X1 U46420 ( .A1(n62731), .A2(n67346), .B1(n62927), .B2(n67340), .ZN(
        n65741) );
  OAI22_X1 U46421 ( .A1(n62730), .A2(n67346), .B1(n62926), .B2(n67340), .ZN(
        n65723) );
  OAI22_X1 U46422 ( .A1(n62729), .A2(n67346), .B1(n62925), .B2(n67340), .ZN(
        n65705) );
  OAI22_X1 U46423 ( .A1(n62728), .A2(n67346), .B1(n62924), .B2(n67340), .ZN(
        n65687) );
  OAI22_X1 U46424 ( .A1(n62727), .A2(n67346), .B1(n62923), .B2(n67340), .ZN(
        n65669) );
  OAI22_X1 U46425 ( .A1(n62726), .A2(n67346), .B1(n62922), .B2(n67340), .ZN(
        n65651) );
  OAI22_X1 U46426 ( .A1(n62725), .A2(n67347), .B1(n62921), .B2(n67341), .ZN(
        n65633) );
  OAI22_X1 U46427 ( .A1(n62724), .A2(n67347), .B1(n62920), .B2(n67341), .ZN(
        n65615) );
  OAI22_X1 U46428 ( .A1(n62723), .A2(n67347), .B1(n62919), .B2(n67341), .ZN(
        n65597) );
  OAI22_X1 U46429 ( .A1(n62722), .A2(n67347), .B1(n62918), .B2(n67341), .ZN(
        n65579) );
  OAI22_X1 U46430 ( .A1(n62721), .A2(n67347), .B1(n62917), .B2(n67341), .ZN(
        n65561) );
  OAI22_X1 U46431 ( .A1(n62720), .A2(n67347), .B1(n62916), .B2(n67341), .ZN(
        n65543) );
  OAI22_X1 U46432 ( .A1(n62719), .A2(n67347), .B1(n62915), .B2(n67341), .ZN(
        n65525) );
  OAI22_X1 U46433 ( .A1(n62718), .A2(n67347), .B1(n62914), .B2(n67341), .ZN(
        n65507) );
  OAI22_X1 U46434 ( .A1(n62717), .A2(n67347), .B1(n62913), .B2(n67341), .ZN(
        n65489) );
  OAI22_X1 U46435 ( .A1(n62716), .A2(n67347), .B1(n62912), .B2(n67341), .ZN(
        n65471) );
  OAI22_X1 U46436 ( .A1(n62715), .A2(n67347), .B1(n62911), .B2(n67341), .ZN(
        n65453) );
  OAI22_X1 U46437 ( .A1(n62714), .A2(n67347), .B1(n62910), .B2(n67341), .ZN(
        n65435) );
  OAI22_X1 U46438 ( .A1(n62713), .A2(n67348), .B1(n62909), .B2(n67342), .ZN(
        n65417) );
  OAI22_X1 U46439 ( .A1(n62712), .A2(n67348), .B1(n62908), .B2(n67342), .ZN(
        n65399) );
  OAI22_X1 U46440 ( .A1(n62711), .A2(n67348), .B1(n62907), .B2(n67342), .ZN(
        n65381) );
  OAI22_X1 U46441 ( .A1(n62710), .A2(n67348), .B1(n62906), .B2(n67342), .ZN(
        n65363) );
  OAI22_X1 U46442 ( .A1(n62709), .A2(n67348), .B1(n62905), .B2(n67342), .ZN(
        n65345) );
  OAI22_X1 U46443 ( .A1(n62708), .A2(n67348), .B1(n62904), .B2(n67342), .ZN(
        n65327) );
  OAI22_X1 U46444 ( .A1(n62707), .A2(n67348), .B1(n62903), .B2(n67342), .ZN(
        n65309) );
  OAI22_X1 U46445 ( .A1(n62706), .A2(n67348), .B1(n62902), .B2(n67342), .ZN(
        n65291) );
  OAI22_X1 U46446 ( .A1(n62705), .A2(n67348), .B1(n62901), .B2(n67342), .ZN(
        n65273) );
  OAI22_X1 U46447 ( .A1(n62704), .A2(n67348), .B1(n62900), .B2(n67342), .ZN(
        n65255) );
  OAI22_X1 U46448 ( .A1(n62703), .A2(n67348), .B1(n62899), .B2(n67342), .ZN(
        n65237) );
  OAI22_X1 U46449 ( .A1(n62702), .A2(n67348), .B1(n62898), .B2(n67342), .ZN(
        n65219) );
  OAI22_X1 U46450 ( .A1(n62155), .A2(n67290), .B1(n62222), .B2(n67284), .ZN(
        n66298) );
  OAI22_X1 U46451 ( .A1(n63494), .A2(n67266), .B1(n62289), .B2(n67260), .ZN(
        n66300) );
  OAI22_X1 U46452 ( .A1(n62154), .A2(n67290), .B1(n62221), .B2(n67284), .ZN(
        n66265) );
  OAI22_X1 U46453 ( .A1(n63493), .A2(n67266), .B1(n62288), .B2(n67260), .ZN(
        n66266) );
  OAI22_X1 U46454 ( .A1(n62153), .A2(n67290), .B1(n62220), .B2(n67284), .ZN(
        n66247) );
  OAI22_X1 U46455 ( .A1(n63492), .A2(n67266), .B1(n62287), .B2(n67260), .ZN(
        n66248) );
  OAI22_X1 U46456 ( .A1(n62152), .A2(n67290), .B1(n62219), .B2(n67284), .ZN(
        n66229) );
  OAI22_X1 U46457 ( .A1(n63491), .A2(n67266), .B1(n62286), .B2(n67260), .ZN(
        n66230) );
  OAI22_X1 U46458 ( .A1(n62151), .A2(n67290), .B1(n62218), .B2(n67284), .ZN(
        n66211) );
  OAI22_X1 U46459 ( .A1(n63490), .A2(n67266), .B1(n62285), .B2(n67260), .ZN(
        n66212) );
  OAI22_X1 U46460 ( .A1(n62150), .A2(n67290), .B1(n62217), .B2(n67284), .ZN(
        n66193) );
  OAI22_X1 U46461 ( .A1(n63489), .A2(n67266), .B1(n62284), .B2(n67260), .ZN(
        n66194) );
  OAI22_X1 U46462 ( .A1(n62149), .A2(n67290), .B1(n62216), .B2(n67284), .ZN(
        n66175) );
  OAI22_X1 U46463 ( .A1(n63488), .A2(n67266), .B1(n62283), .B2(n67260), .ZN(
        n66176) );
  OAI22_X1 U46464 ( .A1(n62148), .A2(n67290), .B1(n62215), .B2(n67284), .ZN(
        n66157) );
  OAI22_X1 U46465 ( .A1(n63487), .A2(n67266), .B1(n62282), .B2(n67260), .ZN(
        n66158) );
  OAI22_X1 U46466 ( .A1(n62147), .A2(n67290), .B1(n62214), .B2(n67284), .ZN(
        n66139) );
  OAI22_X1 U46467 ( .A1(n63486), .A2(n67266), .B1(n62281), .B2(n67260), .ZN(
        n66140) );
  OAI22_X1 U46468 ( .A1(n62146), .A2(n67290), .B1(n62213), .B2(n67284), .ZN(
        n66121) );
  OAI22_X1 U46469 ( .A1(n63485), .A2(n67266), .B1(n62280), .B2(n67260), .ZN(
        n66122) );
  OAI22_X1 U46470 ( .A1(n62145), .A2(n67290), .B1(n62212), .B2(n67284), .ZN(
        n66103) );
  OAI22_X1 U46471 ( .A1(n63484), .A2(n67266), .B1(n62279), .B2(n67260), .ZN(
        n66104) );
  OAI22_X1 U46472 ( .A1(n62144), .A2(n67290), .B1(n62211), .B2(n67284), .ZN(
        n66085) );
  OAI22_X1 U46473 ( .A1(n63483), .A2(n67266), .B1(n62278), .B2(n67260), .ZN(
        n66086) );
  OAI22_X1 U46474 ( .A1(n62143), .A2(n67291), .B1(n62210), .B2(n67285), .ZN(
        n66067) );
  OAI22_X1 U46475 ( .A1(n63482), .A2(n67267), .B1(n62277), .B2(n67261), .ZN(
        n66068) );
  OAI22_X1 U46476 ( .A1(n62142), .A2(n67291), .B1(n62209), .B2(n67285), .ZN(
        n66049) );
  OAI22_X1 U46477 ( .A1(n63481), .A2(n67267), .B1(n62276), .B2(n67261), .ZN(
        n66050) );
  OAI22_X1 U46478 ( .A1(n62141), .A2(n67291), .B1(n62208), .B2(n67285), .ZN(
        n66031) );
  OAI22_X1 U46479 ( .A1(n63480), .A2(n67267), .B1(n62275), .B2(n67261), .ZN(
        n66032) );
  OAI22_X1 U46480 ( .A1(n62140), .A2(n67291), .B1(n62207), .B2(n67285), .ZN(
        n66013) );
  OAI22_X1 U46481 ( .A1(n63479), .A2(n67267), .B1(n62274), .B2(n67261), .ZN(
        n66014) );
  OAI22_X1 U46482 ( .A1(n62139), .A2(n67291), .B1(n62206), .B2(n67285), .ZN(
        n65995) );
  OAI22_X1 U46483 ( .A1(n63478), .A2(n67267), .B1(n62273), .B2(n67261), .ZN(
        n65996) );
  OAI22_X1 U46484 ( .A1(n62138), .A2(n67291), .B1(n62205), .B2(n67285), .ZN(
        n65977) );
  OAI22_X1 U46485 ( .A1(n63477), .A2(n67267), .B1(n62272), .B2(n67261), .ZN(
        n65978) );
  OAI22_X1 U46486 ( .A1(n62137), .A2(n67291), .B1(n62204), .B2(n67285), .ZN(
        n65959) );
  OAI22_X1 U46487 ( .A1(n63476), .A2(n67267), .B1(n62271), .B2(n67261), .ZN(
        n65960) );
  OAI22_X1 U46488 ( .A1(n62136), .A2(n67291), .B1(n62203), .B2(n67285), .ZN(
        n65941) );
  OAI22_X1 U46489 ( .A1(n63475), .A2(n67267), .B1(n62270), .B2(n67261), .ZN(
        n65942) );
  OAI22_X1 U46490 ( .A1(n62135), .A2(n67291), .B1(n62202), .B2(n67285), .ZN(
        n65923) );
  OAI22_X1 U46491 ( .A1(n63474), .A2(n67267), .B1(n62269), .B2(n67261), .ZN(
        n65924) );
  OAI22_X1 U46492 ( .A1(n62134), .A2(n67291), .B1(n62201), .B2(n67285), .ZN(
        n65905) );
  OAI22_X1 U46493 ( .A1(n63473), .A2(n67267), .B1(n62268), .B2(n67261), .ZN(
        n65906) );
  OAI22_X1 U46494 ( .A1(n62133), .A2(n67291), .B1(n62200), .B2(n67285), .ZN(
        n65887) );
  OAI22_X1 U46495 ( .A1(n63472), .A2(n67267), .B1(n62267), .B2(n67261), .ZN(
        n65888) );
  OAI22_X1 U46496 ( .A1(n62132), .A2(n67291), .B1(n62199), .B2(n67285), .ZN(
        n65869) );
  OAI22_X1 U46497 ( .A1(n63471), .A2(n67267), .B1(n62266), .B2(n67261), .ZN(
        n65870) );
  OAI22_X1 U46498 ( .A1(n62131), .A2(n67292), .B1(n62198), .B2(n67286), .ZN(
        n65851) );
  OAI22_X1 U46499 ( .A1(n63470), .A2(n67268), .B1(n62265), .B2(n67262), .ZN(
        n65852) );
  OAI22_X1 U46500 ( .A1(n62130), .A2(n67292), .B1(n62197), .B2(n67286), .ZN(
        n65833) );
  OAI22_X1 U46501 ( .A1(n63469), .A2(n67268), .B1(n62264), .B2(n67262), .ZN(
        n65834) );
  OAI22_X1 U46502 ( .A1(n62129), .A2(n67292), .B1(n62196), .B2(n67286), .ZN(
        n65815) );
  OAI22_X1 U46503 ( .A1(n63468), .A2(n67268), .B1(n62263), .B2(n67262), .ZN(
        n65816) );
  OAI22_X1 U46504 ( .A1(n62128), .A2(n67292), .B1(n62195), .B2(n67286), .ZN(
        n65797) );
  OAI22_X1 U46505 ( .A1(n63467), .A2(n67268), .B1(n62262), .B2(n67262), .ZN(
        n65798) );
  OAI22_X1 U46506 ( .A1(n62127), .A2(n67292), .B1(n62194), .B2(n67286), .ZN(
        n65779) );
  OAI22_X1 U46507 ( .A1(n63466), .A2(n67268), .B1(n62261), .B2(n67262), .ZN(
        n65780) );
  OAI22_X1 U46508 ( .A1(n62126), .A2(n67292), .B1(n62193), .B2(n67286), .ZN(
        n65761) );
  OAI22_X1 U46509 ( .A1(n63465), .A2(n67268), .B1(n62260), .B2(n67262), .ZN(
        n65762) );
  OAI22_X1 U46510 ( .A1(n62125), .A2(n67292), .B1(n62192), .B2(n67286), .ZN(
        n65743) );
  OAI22_X1 U46511 ( .A1(n63464), .A2(n67268), .B1(n62259), .B2(n67262), .ZN(
        n65744) );
  OAI22_X1 U46512 ( .A1(n62124), .A2(n67292), .B1(n62191), .B2(n67286), .ZN(
        n65725) );
  OAI22_X1 U46513 ( .A1(n63463), .A2(n67268), .B1(n62258), .B2(n67262), .ZN(
        n65726) );
  OAI22_X1 U46514 ( .A1(n62123), .A2(n67292), .B1(n62190), .B2(n67286), .ZN(
        n65707) );
  OAI22_X1 U46515 ( .A1(n63462), .A2(n67268), .B1(n62257), .B2(n67262), .ZN(
        n65708) );
  OAI22_X1 U46516 ( .A1(n62122), .A2(n67292), .B1(n62189), .B2(n67286), .ZN(
        n65689) );
  OAI22_X1 U46517 ( .A1(n63461), .A2(n67268), .B1(n62256), .B2(n67262), .ZN(
        n65690) );
  OAI22_X1 U46518 ( .A1(n62121), .A2(n67292), .B1(n62188), .B2(n67286), .ZN(
        n65671) );
  OAI22_X1 U46519 ( .A1(n63460), .A2(n67268), .B1(n62255), .B2(n67262), .ZN(
        n65672) );
  OAI22_X1 U46520 ( .A1(n62120), .A2(n67292), .B1(n62187), .B2(n67286), .ZN(
        n65653) );
  OAI22_X1 U46521 ( .A1(n63459), .A2(n67268), .B1(n62254), .B2(n67262), .ZN(
        n65654) );
  OAI22_X1 U46522 ( .A1(n62119), .A2(n67293), .B1(n62186), .B2(n67287), .ZN(
        n65635) );
  OAI22_X1 U46523 ( .A1(n63458), .A2(n67269), .B1(n62253), .B2(n67263), .ZN(
        n65636) );
  OAI22_X1 U46524 ( .A1(n62118), .A2(n67293), .B1(n62185), .B2(n67287), .ZN(
        n65617) );
  OAI22_X1 U46525 ( .A1(n63457), .A2(n67269), .B1(n62252), .B2(n67263), .ZN(
        n65618) );
  OAI22_X1 U46526 ( .A1(n62117), .A2(n67293), .B1(n62184), .B2(n67287), .ZN(
        n65599) );
  OAI22_X1 U46527 ( .A1(n63456), .A2(n67269), .B1(n62251), .B2(n67263), .ZN(
        n65600) );
  OAI22_X1 U46528 ( .A1(n62116), .A2(n67293), .B1(n62183), .B2(n67287), .ZN(
        n65581) );
  OAI22_X1 U46529 ( .A1(n63455), .A2(n67269), .B1(n62250), .B2(n67263), .ZN(
        n65582) );
  OAI22_X1 U46530 ( .A1(n62115), .A2(n67293), .B1(n62182), .B2(n67287), .ZN(
        n65563) );
  OAI22_X1 U46531 ( .A1(n63454), .A2(n67269), .B1(n62249), .B2(n67263), .ZN(
        n65564) );
  OAI22_X1 U46532 ( .A1(n62114), .A2(n67293), .B1(n62181), .B2(n67287), .ZN(
        n65545) );
  OAI22_X1 U46533 ( .A1(n63453), .A2(n67269), .B1(n62248), .B2(n67263), .ZN(
        n65546) );
  OAI22_X1 U46534 ( .A1(n62113), .A2(n67293), .B1(n62180), .B2(n67287), .ZN(
        n65527) );
  OAI22_X1 U46535 ( .A1(n63452), .A2(n67269), .B1(n62247), .B2(n67263), .ZN(
        n65528) );
  OAI22_X1 U46536 ( .A1(n62112), .A2(n67293), .B1(n62179), .B2(n67287), .ZN(
        n65509) );
  OAI22_X1 U46537 ( .A1(n63451), .A2(n67269), .B1(n62246), .B2(n67263), .ZN(
        n65510) );
  OAI22_X1 U46538 ( .A1(n62111), .A2(n67293), .B1(n62178), .B2(n67287), .ZN(
        n65491) );
  OAI22_X1 U46539 ( .A1(n63450), .A2(n67269), .B1(n62245), .B2(n67263), .ZN(
        n65492) );
  OAI22_X1 U46540 ( .A1(n62110), .A2(n67293), .B1(n62177), .B2(n67287), .ZN(
        n65473) );
  OAI22_X1 U46541 ( .A1(n63449), .A2(n67269), .B1(n62244), .B2(n67263), .ZN(
        n65474) );
  OAI22_X1 U46542 ( .A1(n62109), .A2(n67293), .B1(n62176), .B2(n67287), .ZN(
        n65455) );
  OAI22_X1 U46543 ( .A1(n63448), .A2(n67269), .B1(n62243), .B2(n67263), .ZN(
        n65456) );
  OAI22_X1 U46544 ( .A1(n62108), .A2(n67293), .B1(n62175), .B2(n67287), .ZN(
        n65437) );
  OAI22_X1 U46545 ( .A1(n63447), .A2(n67269), .B1(n62242), .B2(n67263), .ZN(
        n65438) );
  OAI22_X1 U46546 ( .A1(n62107), .A2(n67294), .B1(n62174), .B2(n67288), .ZN(
        n65419) );
  OAI22_X1 U46547 ( .A1(n63446), .A2(n67270), .B1(n62241), .B2(n67264), .ZN(
        n65420) );
  OAI22_X1 U46548 ( .A1(n62106), .A2(n67294), .B1(n62173), .B2(n67288), .ZN(
        n65401) );
  OAI22_X1 U46549 ( .A1(n63445), .A2(n67270), .B1(n62240), .B2(n67264), .ZN(
        n65402) );
  OAI22_X1 U46550 ( .A1(n62105), .A2(n67294), .B1(n62172), .B2(n67288), .ZN(
        n65383) );
  OAI22_X1 U46551 ( .A1(n63444), .A2(n67270), .B1(n62239), .B2(n67264), .ZN(
        n65384) );
  OAI22_X1 U46552 ( .A1(n62104), .A2(n67294), .B1(n62171), .B2(n67288), .ZN(
        n65365) );
  OAI22_X1 U46553 ( .A1(n63443), .A2(n67270), .B1(n62238), .B2(n67264), .ZN(
        n65366) );
  OAI22_X1 U46554 ( .A1(n62103), .A2(n67294), .B1(n62170), .B2(n67288), .ZN(
        n65347) );
  OAI22_X1 U46555 ( .A1(n63442), .A2(n67270), .B1(n62237), .B2(n67264), .ZN(
        n65348) );
  OAI22_X1 U46556 ( .A1(n62102), .A2(n67294), .B1(n62169), .B2(n67288), .ZN(
        n65329) );
  OAI22_X1 U46557 ( .A1(n63441), .A2(n67270), .B1(n62236), .B2(n67264), .ZN(
        n65330) );
  OAI22_X1 U46558 ( .A1(n62101), .A2(n67294), .B1(n62168), .B2(n67288), .ZN(
        n65311) );
  OAI22_X1 U46559 ( .A1(n63440), .A2(n67270), .B1(n62235), .B2(n67264), .ZN(
        n65312) );
  OAI22_X1 U46560 ( .A1(n62100), .A2(n67294), .B1(n62167), .B2(n67288), .ZN(
        n65293) );
  OAI22_X1 U46561 ( .A1(n63439), .A2(n67270), .B1(n62234), .B2(n67264), .ZN(
        n65294) );
  OAI22_X1 U46562 ( .A1(n62099), .A2(n67294), .B1(n62166), .B2(n67288), .ZN(
        n65275) );
  OAI22_X1 U46563 ( .A1(n63438), .A2(n67270), .B1(n62233), .B2(n67264), .ZN(
        n65276) );
  OAI22_X1 U46564 ( .A1(n62098), .A2(n67294), .B1(n62165), .B2(n67288), .ZN(
        n65257) );
  OAI22_X1 U46565 ( .A1(n63437), .A2(n67270), .B1(n62232), .B2(n67264), .ZN(
        n65258) );
  OAI22_X1 U46566 ( .A1(n62097), .A2(n67294), .B1(n62164), .B2(n67288), .ZN(
        n65239) );
  OAI22_X1 U46567 ( .A1(n63436), .A2(n67270), .B1(n62231), .B2(n67264), .ZN(
        n65240) );
  OAI22_X1 U46568 ( .A1(n62096), .A2(n67294), .B1(n62163), .B2(n67288), .ZN(
        n65221) );
  OAI22_X1 U46569 ( .A1(n63435), .A2(n67270), .B1(n62230), .B2(n67264), .ZN(
        n65222) );
  OAI22_X1 U46570 ( .A1(n63361), .A2(n67488), .B1(n63697), .B2(n67482), .ZN(
        n65096) );
  OAI22_X1 U46571 ( .A1(n62761), .A2(n67464), .B1(n62222), .B2(n67458), .ZN(
        n65098) );
  OAI22_X1 U46572 ( .A1(n63360), .A2(n67488), .B1(n63696), .B2(n67482), .ZN(
        n65061) );
  OAI22_X1 U46573 ( .A1(n62760), .A2(n67464), .B1(n62221), .B2(n67458), .ZN(
        n65062) );
  OAI22_X1 U46574 ( .A1(n63359), .A2(n67488), .B1(n63695), .B2(n67482), .ZN(
        n65041) );
  OAI22_X1 U46575 ( .A1(n62759), .A2(n67464), .B1(n62220), .B2(n67458), .ZN(
        n65042) );
  OAI22_X1 U46576 ( .A1(n63358), .A2(n67488), .B1(n63694), .B2(n67482), .ZN(
        n65021) );
  OAI22_X1 U46577 ( .A1(n62758), .A2(n67464), .B1(n62219), .B2(n67458), .ZN(
        n65022) );
  OAI22_X1 U46578 ( .A1(n63357), .A2(n67488), .B1(n63693), .B2(n67482), .ZN(
        n65001) );
  OAI22_X1 U46579 ( .A1(n62757), .A2(n67464), .B1(n62218), .B2(n67458), .ZN(
        n65002) );
  OAI22_X1 U46580 ( .A1(n63356), .A2(n67488), .B1(n63692), .B2(n67482), .ZN(
        n64981) );
  OAI22_X1 U46581 ( .A1(n62756), .A2(n67464), .B1(n62217), .B2(n67458), .ZN(
        n64982) );
  OAI22_X1 U46582 ( .A1(n63355), .A2(n67488), .B1(n63691), .B2(n67482), .ZN(
        n64961) );
  OAI22_X1 U46583 ( .A1(n62755), .A2(n67464), .B1(n62216), .B2(n67458), .ZN(
        n64962) );
  OAI22_X1 U46584 ( .A1(n63354), .A2(n67488), .B1(n63690), .B2(n67482), .ZN(
        n64941) );
  OAI22_X1 U46585 ( .A1(n62754), .A2(n67464), .B1(n62215), .B2(n67458), .ZN(
        n64942) );
  OAI22_X1 U46586 ( .A1(n63353), .A2(n67488), .B1(n63689), .B2(n67482), .ZN(
        n64921) );
  OAI22_X1 U46587 ( .A1(n62753), .A2(n67464), .B1(n62214), .B2(n67458), .ZN(
        n64922) );
  OAI22_X1 U46588 ( .A1(n63352), .A2(n67488), .B1(n63688), .B2(n67482), .ZN(
        n64901) );
  OAI22_X1 U46589 ( .A1(n62752), .A2(n67464), .B1(n62213), .B2(n67458), .ZN(
        n64902) );
  OAI22_X1 U46590 ( .A1(n63351), .A2(n67488), .B1(n63687), .B2(n67482), .ZN(
        n64881) );
  OAI22_X1 U46591 ( .A1(n62751), .A2(n67464), .B1(n62212), .B2(n67458), .ZN(
        n64882) );
  OAI22_X1 U46592 ( .A1(n63350), .A2(n67488), .B1(n63686), .B2(n67482), .ZN(
        n64861) );
  OAI22_X1 U46593 ( .A1(n62750), .A2(n67464), .B1(n62211), .B2(n67458), .ZN(
        n64862) );
  OAI22_X1 U46594 ( .A1(n63349), .A2(n67489), .B1(n63685), .B2(n67483), .ZN(
        n64841) );
  OAI22_X1 U46595 ( .A1(n62749), .A2(n67465), .B1(n62210), .B2(n67459), .ZN(
        n64842) );
  OAI22_X1 U46596 ( .A1(n63348), .A2(n67489), .B1(n63684), .B2(n67483), .ZN(
        n64821) );
  OAI22_X1 U46597 ( .A1(n62748), .A2(n67465), .B1(n62209), .B2(n67459), .ZN(
        n64822) );
  OAI22_X1 U46598 ( .A1(n63347), .A2(n67489), .B1(n63683), .B2(n67483), .ZN(
        n64801) );
  OAI22_X1 U46599 ( .A1(n62747), .A2(n67465), .B1(n62208), .B2(n67459), .ZN(
        n64802) );
  OAI22_X1 U46600 ( .A1(n63346), .A2(n67489), .B1(n63682), .B2(n67483), .ZN(
        n64781) );
  OAI22_X1 U46601 ( .A1(n62746), .A2(n67465), .B1(n62207), .B2(n67459), .ZN(
        n64782) );
  OAI22_X1 U46602 ( .A1(n63345), .A2(n67489), .B1(n63681), .B2(n67483), .ZN(
        n64761) );
  OAI22_X1 U46603 ( .A1(n62745), .A2(n67465), .B1(n62206), .B2(n67459), .ZN(
        n64762) );
  OAI22_X1 U46604 ( .A1(n63344), .A2(n67489), .B1(n63680), .B2(n67483), .ZN(
        n64741) );
  OAI22_X1 U46605 ( .A1(n62744), .A2(n67465), .B1(n62205), .B2(n67459), .ZN(
        n64742) );
  OAI22_X1 U46606 ( .A1(n63343), .A2(n67489), .B1(n63679), .B2(n67483), .ZN(
        n64721) );
  OAI22_X1 U46607 ( .A1(n62743), .A2(n67465), .B1(n62204), .B2(n67459), .ZN(
        n64722) );
  OAI22_X1 U46608 ( .A1(n63342), .A2(n67489), .B1(n63678), .B2(n67483), .ZN(
        n64701) );
  OAI22_X1 U46609 ( .A1(n62742), .A2(n67465), .B1(n62203), .B2(n67459), .ZN(
        n64702) );
  OAI22_X1 U46610 ( .A1(n63341), .A2(n67489), .B1(n63677), .B2(n67483), .ZN(
        n64681) );
  OAI22_X1 U46611 ( .A1(n62741), .A2(n67465), .B1(n62202), .B2(n67459), .ZN(
        n64682) );
  OAI22_X1 U46612 ( .A1(n63340), .A2(n67489), .B1(n63676), .B2(n67483), .ZN(
        n64661) );
  OAI22_X1 U46613 ( .A1(n62740), .A2(n67465), .B1(n62201), .B2(n67459), .ZN(
        n64662) );
  OAI22_X1 U46614 ( .A1(n63339), .A2(n67489), .B1(n63675), .B2(n67483), .ZN(
        n64641) );
  OAI22_X1 U46615 ( .A1(n62739), .A2(n67465), .B1(n62200), .B2(n67459), .ZN(
        n64642) );
  OAI22_X1 U46616 ( .A1(n63338), .A2(n67489), .B1(n63674), .B2(n67483), .ZN(
        n64621) );
  OAI22_X1 U46617 ( .A1(n62738), .A2(n67465), .B1(n62199), .B2(n67459), .ZN(
        n64622) );
  OAI22_X1 U46618 ( .A1(n63337), .A2(n67490), .B1(n63673), .B2(n67484), .ZN(
        n64601) );
  OAI22_X1 U46619 ( .A1(n62737), .A2(n67466), .B1(n62198), .B2(n67460), .ZN(
        n64602) );
  OAI22_X1 U46620 ( .A1(n63336), .A2(n67490), .B1(n63672), .B2(n67484), .ZN(
        n64581) );
  OAI22_X1 U46621 ( .A1(n62736), .A2(n67466), .B1(n62197), .B2(n67460), .ZN(
        n64582) );
  OAI22_X1 U46622 ( .A1(n63335), .A2(n67490), .B1(n63671), .B2(n67484), .ZN(
        n64561) );
  OAI22_X1 U46623 ( .A1(n62735), .A2(n67466), .B1(n62196), .B2(n67460), .ZN(
        n64562) );
  OAI22_X1 U46624 ( .A1(n63334), .A2(n67490), .B1(n63670), .B2(n67484), .ZN(
        n64541) );
  OAI22_X1 U46625 ( .A1(n62734), .A2(n67466), .B1(n62195), .B2(n67460), .ZN(
        n64542) );
  OAI22_X1 U46626 ( .A1(n63333), .A2(n67490), .B1(n63669), .B2(n67484), .ZN(
        n64521) );
  OAI22_X1 U46627 ( .A1(n62733), .A2(n67466), .B1(n62194), .B2(n67460), .ZN(
        n64522) );
  OAI22_X1 U46628 ( .A1(n63332), .A2(n67490), .B1(n63668), .B2(n67484), .ZN(
        n64501) );
  OAI22_X1 U46629 ( .A1(n62732), .A2(n67466), .B1(n62193), .B2(n67460), .ZN(
        n64502) );
  OAI22_X1 U46630 ( .A1(n63331), .A2(n67490), .B1(n63667), .B2(n67484), .ZN(
        n64481) );
  OAI22_X1 U46631 ( .A1(n62731), .A2(n67466), .B1(n62192), .B2(n67460), .ZN(
        n64482) );
  OAI22_X1 U46632 ( .A1(n63330), .A2(n67490), .B1(n63666), .B2(n67484), .ZN(
        n64461) );
  OAI22_X1 U46633 ( .A1(n62730), .A2(n67466), .B1(n62191), .B2(n67460), .ZN(
        n64462) );
  OAI22_X1 U46634 ( .A1(n63329), .A2(n67490), .B1(n63665), .B2(n67484), .ZN(
        n64441) );
  OAI22_X1 U46635 ( .A1(n62729), .A2(n67466), .B1(n62190), .B2(n67460), .ZN(
        n64442) );
  OAI22_X1 U46636 ( .A1(n63328), .A2(n67490), .B1(n63664), .B2(n67484), .ZN(
        n64421) );
  OAI22_X1 U46637 ( .A1(n62728), .A2(n67466), .B1(n62189), .B2(n67460), .ZN(
        n64422) );
  OAI22_X1 U46638 ( .A1(n63327), .A2(n67490), .B1(n63663), .B2(n67484), .ZN(
        n64401) );
  OAI22_X1 U46639 ( .A1(n62727), .A2(n67466), .B1(n62188), .B2(n67460), .ZN(
        n64402) );
  OAI22_X1 U46640 ( .A1(n63326), .A2(n67490), .B1(n63662), .B2(n67484), .ZN(
        n64381) );
  OAI22_X1 U46641 ( .A1(n62726), .A2(n67466), .B1(n62187), .B2(n67460), .ZN(
        n64382) );
  OAI22_X1 U46642 ( .A1(n63325), .A2(n67491), .B1(n63661), .B2(n67485), .ZN(
        n64361) );
  OAI22_X1 U46643 ( .A1(n62725), .A2(n67467), .B1(n62186), .B2(n67461), .ZN(
        n64362) );
  OAI22_X1 U46644 ( .A1(n63324), .A2(n67491), .B1(n63660), .B2(n67485), .ZN(
        n64341) );
  OAI22_X1 U46645 ( .A1(n62724), .A2(n67467), .B1(n62185), .B2(n67461), .ZN(
        n64342) );
  OAI22_X1 U46646 ( .A1(n63323), .A2(n67491), .B1(n63659), .B2(n67485), .ZN(
        n64321) );
  OAI22_X1 U46647 ( .A1(n62723), .A2(n67467), .B1(n62184), .B2(n67461), .ZN(
        n64322) );
  OAI22_X1 U46648 ( .A1(n63322), .A2(n67491), .B1(n63658), .B2(n67485), .ZN(
        n64301) );
  OAI22_X1 U46649 ( .A1(n62722), .A2(n67467), .B1(n62183), .B2(n67461), .ZN(
        n64302) );
  OAI22_X1 U46650 ( .A1(n63321), .A2(n67491), .B1(n63657), .B2(n67485), .ZN(
        n64281) );
  OAI22_X1 U46651 ( .A1(n62721), .A2(n67467), .B1(n62182), .B2(n67461), .ZN(
        n64282) );
  OAI22_X1 U46652 ( .A1(n63320), .A2(n67491), .B1(n63656), .B2(n67485), .ZN(
        n64261) );
  OAI22_X1 U46653 ( .A1(n62720), .A2(n67467), .B1(n62181), .B2(n67461), .ZN(
        n64262) );
  OAI22_X1 U46654 ( .A1(n63319), .A2(n67491), .B1(n63655), .B2(n67485), .ZN(
        n64241) );
  OAI22_X1 U46655 ( .A1(n62719), .A2(n67467), .B1(n62180), .B2(n67461), .ZN(
        n64242) );
  OAI22_X1 U46656 ( .A1(n63318), .A2(n67491), .B1(n63654), .B2(n67485), .ZN(
        n64221) );
  OAI22_X1 U46657 ( .A1(n62718), .A2(n67467), .B1(n62179), .B2(n67461), .ZN(
        n64222) );
  OAI22_X1 U46658 ( .A1(n63317), .A2(n67491), .B1(n63653), .B2(n67485), .ZN(
        n64201) );
  OAI22_X1 U46659 ( .A1(n62717), .A2(n67467), .B1(n62178), .B2(n67461), .ZN(
        n64202) );
  OAI22_X1 U46660 ( .A1(n63316), .A2(n67491), .B1(n63652), .B2(n67485), .ZN(
        n64181) );
  OAI22_X1 U46661 ( .A1(n62716), .A2(n67467), .B1(n62177), .B2(n67461), .ZN(
        n64182) );
  OAI22_X1 U46662 ( .A1(n63315), .A2(n67491), .B1(n63651), .B2(n67485), .ZN(
        n64161) );
  OAI22_X1 U46663 ( .A1(n62715), .A2(n67467), .B1(n62176), .B2(n67461), .ZN(
        n64162) );
  OAI22_X1 U46664 ( .A1(n63314), .A2(n67491), .B1(n63650), .B2(n67485), .ZN(
        n64141) );
  OAI22_X1 U46665 ( .A1(n62714), .A2(n67467), .B1(n62175), .B2(n67461), .ZN(
        n64142) );
  OAI22_X1 U46666 ( .A1(n63313), .A2(n67492), .B1(n63649), .B2(n67486), .ZN(
        n64121) );
  OAI22_X1 U46667 ( .A1(n62713), .A2(n67468), .B1(n62174), .B2(n67462), .ZN(
        n64122) );
  OAI22_X1 U46668 ( .A1(n63312), .A2(n67492), .B1(n63648), .B2(n67486), .ZN(
        n64101) );
  OAI22_X1 U46669 ( .A1(n62712), .A2(n67468), .B1(n62173), .B2(n67462), .ZN(
        n64102) );
  OAI22_X1 U46670 ( .A1(n63311), .A2(n67492), .B1(n63647), .B2(n67486), .ZN(
        n64081) );
  OAI22_X1 U46671 ( .A1(n62711), .A2(n67468), .B1(n62172), .B2(n67462), .ZN(
        n64082) );
  OAI22_X1 U46672 ( .A1(n63310), .A2(n67492), .B1(n63646), .B2(n67486), .ZN(
        n64061) );
  OAI22_X1 U46673 ( .A1(n62710), .A2(n67468), .B1(n62171), .B2(n67462), .ZN(
        n64062) );
  OAI22_X1 U46674 ( .A1(n63309), .A2(n67492), .B1(n63645), .B2(n67486), .ZN(
        n64041) );
  OAI22_X1 U46675 ( .A1(n62709), .A2(n67468), .B1(n62170), .B2(n67462), .ZN(
        n64042) );
  OAI22_X1 U46676 ( .A1(n63308), .A2(n67492), .B1(n63644), .B2(n67486), .ZN(
        n64021) );
  OAI22_X1 U46677 ( .A1(n62708), .A2(n67468), .B1(n62169), .B2(n67462), .ZN(
        n64022) );
  OAI22_X1 U46678 ( .A1(n63307), .A2(n67492), .B1(n63643), .B2(n67486), .ZN(
        n64001) );
  OAI22_X1 U46679 ( .A1(n62707), .A2(n67468), .B1(n62168), .B2(n67462), .ZN(
        n64002) );
  OAI22_X1 U46680 ( .A1(n63306), .A2(n67492), .B1(n63642), .B2(n67486), .ZN(
        n63981) );
  OAI22_X1 U46681 ( .A1(n62706), .A2(n67468), .B1(n62167), .B2(n67462), .ZN(
        n63982) );
  OAI22_X1 U46682 ( .A1(n63305), .A2(n67492), .B1(n63641), .B2(n67486), .ZN(
        n63961) );
  OAI22_X1 U46683 ( .A1(n62705), .A2(n67468), .B1(n62166), .B2(n67462), .ZN(
        n63962) );
  OAI22_X1 U46684 ( .A1(n63304), .A2(n67492), .B1(n63640), .B2(n67486), .ZN(
        n63941) );
  OAI22_X1 U46685 ( .A1(n62704), .A2(n67468), .B1(n62165), .B2(n67462), .ZN(
        n63942) );
  OAI22_X1 U46686 ( .A1(n63303), .A2(n67492), .B1(n63639), .B2(n67486), .ZN(
        n63921) );
  OAI22_X1 U46687 ( .A1(n62703), .A2(n67468), .B1(n62164), .B2(n67462), .ZN(
        n63922) );
  OAI22_X1 U46688 ( .A1(n63302), .A2(n67492), .B1(n63638), .B2(n67486), .ZN(
        n63901) );
  OAI22_X1 U46689 ( .A1(n62702), .A2(n67468), .B1(n62163), .B2(n67462), .ZN(
        n63902) );
  OAI22_X1 U46690 ( .A1(n63361), .A2(n67332), .B1(n63091), .B2(n67326), .ZN(
        n66294) );
  OAI22_X1 U46691 ( .A1(n63360), .A2(n67332), .B1(n63090), .B2(n67326), .ZN(
        n66262) );
  OAI22_X1 U46692 ( .A1(n63359), .A2(n67332), .B1(n63089), .B2(n67326), .ZN(
        n66244) );
  OAI22_X1 U46693 ( .A1(n63358), .A2(n67332), .B1(n63088), .B2(n67326), .ZN(
        n66226) );
  OAI22_X1 U46694 ( .A1(n63357), .A2(n67332), .B1(n63087), .B2(n67326), .ZN(
        n66208) );
  OAI22_X1 U46695 ( .A1(n63356), .A2(n67332), .B1(n63086), .B2(n67326), .ZN(
        n66190) );
  OAI22_X1 U46696 ( .A1(n63355), .A2(n67332), .B1(n63085), .B2(n67326), .ZN(
        n66172) );
  OAI22_X1 U46697 ( .A1(n63354), .A2(n67332), .B1(n63084), .B2(n67326), .ZN(
        n66154) );
  OAI22_X1 U46698 ( .A1(n63353), .A2(n67332), .B1(n63083), .B2(n67326), .ZN(
        n66136) );
  OAI22_X1 U46699 ( .A1(n63352), .A2(n67332), .B1(n63082), .B2(n67326), .ZN(
        n66118) );
  OAI22_X1 U46700 ( .A1(n63351), .A2(n67332), .B1(n63081), .B2(n67326), .ZN(
        n66100) );
  OAI22_X1 U46701 ( .A1(n63350), .A2(n67332), .B1(n63080), .B2(n67326), .ZN(
        n66082) );
  OAI22_X1 U46702 ( .A1(n63349), .A2(n67333), .B1(n63079), .B2(n67327), .ZN(
        n66064) );
  OAI22_X1 U46703 ( .A1(n63348), .A2(n67333), .B1(n63078), .B2(n67327), .ZN(
        n66046) );
  OAI22_X1 U46704 ( .A1(n63347), .A2(n67333), .B1(n63077), .B2(n67327), .ZN(
        n66028) );
  OAI22_X1 U46705 ( .A1(n63346), .A2(n67333), .B1(n63076), .B2(n67327), .ZN(
        n66010) );
  OAI22_X1 U46706 ( .A1(n63345), .A2(n67333), .B1(n63075), .B2(n67327), .ZN(
        n65992) );
  OAI22_X1 U46707 ( .A1(n63344), .A2(n67333), .B1(n63074), .B2(n67327), .ZN(
        n65974) );
  OAI22_X1 U46708 ( .A1(n63343), .A2(n67333), .B1(n63073), .B2(n67327), .ZN(
        n65956) );
  OAI22_X1 U46709 ( .A1(n63342), .A2(n67333), .B1(n63072), .B2(n67327), .ZN(
        n65938) );
  OAI22_X1 U46710 ( .A1(n63341), .A2(n67333), .B1(n63071), .B2(n67327), .ZN(
        n65920) );
  OAI22_X1 U46711 ( .A1(n63340), .A2(n67333), .B1(n63070), .B2(n67327), .ZN(
        n65902) );
  OAI22_X1 U46712 ( .A1(n63339), .A2(n67333), .B1(n63069), .B2(n67327), .ZN(
        n65884) );
  OAI22_X1 U46713 ( .A1(n63338), .A2(n67333), .B1(n63068), .B2(n67327), .ZN(
        n65866) );
  OAI22_X1 U46714 ( .A1(n63337), .A2(n67334), .B1(n63067), .B2(n67328), .ZN(
        n65848) );
  OAI22_X1 U46715 ( .A1(n63336), .A2(n67334), .B1(n63066), .B2(n67328), .ZN(
        n65830) );
  OAI22_X1 U46716 ( .A1(n63335), .A2(n67334), .B1(n63065), .B2(n67328), .ZN(
        n65812) );
  OAI22_X1 U46717 ( .A1(n63334), .A2(n67334), .B1(n63064), .B2(n67328), .ZN(
        n65794) );
  OAI22_X1 U46718 ( .A1(n63333), .A2(n67334), .B1(n63063), .B2(n67328), .ZN(
        n65776) );
  OAI22_X1 U46719 ( .A1(n63332), .A2(n67334), .B1(n63062), .B2(n67328), .ZN(
        n65758) );
  OAI22_X1 U46720 ( .A1(n63331), .A2(n67334), .B1(n63061), .B2(n67328), .ZN(
        n65740) );
  OAI22_X1 U46721 ( .A1(n63330), .A2(n67334), .B1(n63060), .B2(n67328), .ZN(
        n65722) );
  OAI22_X1 U46722 ( .A1(n63329), .A2(n67334), .B1(n63059), .B2(n67328), .ZN(
        n65704) );
  OAI22_X1 U46723 ( .A1(n63328), .A2(n67334), .B1(n63058), .B2(n67328), .ZN(
        n65686) );
  OAI22_X1 U46724 ( .A1(n63327), .A2(n67334), .B1(n63057), .B2(n67328), .ZN(
        n65668) );
  OAI22_X1 U46725 ( .A1(n63326), .A2(n67334), .B1(n63056), .B2(n67328), .ZN(
        n65650) );
  OAI22_X1 U46726 ( .A1(n63325), .A2(n67335), .B1(n63055), .B2(n67329), .ZN(
        n65632) );
  OAI22_X1 U46727 ( .A1(n63324), .A2(n67335), .B1(n63054), .B2(n67329), .ZN(
        n65614) );
  OAI22_X1 U46728 ( .A1(n63323), .A2(n67335), .B1(n63053), .B2(n67329), .ZN(
        n65596) );
  OAI22_X1 U46729 ( .A1(n63322), .A2(n67335), .B1(n63052), .B2(n67329), .ZN(
        n65578) );
  OAI22_X1 U46730 ( .A1(n63321), .A2(n67335), .B1(n63051), .B2(n67329), .ZN(
        n65560) );
  OAI22_X1 U46731 ( .A1(n63320), .A2(n67335), .B1(n63050), .B2(n67329), .ZN(
        n65542) );
  OAI22_X1 U46732 ( .A1(n63319), .A2(n67335), .B1(n63049), .B2(n67329), .ZN(
        n65524) );
  OAI22_X1 U46733 ( .A1(n63318), .A2(n67335), .B1(n63048), .B2(n67329), .ZN(
        n65506) );
  OAI22_X1 U46734 ( .A1(n63317), .A2(n67335), .B1(n63047), .B2(n67329), .ZN(
        n65488) );
  OAI22_X1 U46735 ( .A1(n63316), .A2(n67335), .B1(n63046), .B2(n67329), .ZN(
        n65470) );
  OAI22_X1 U46736 ( .A1(n63315), .A2(n67335), .B1(n63045), .B2(n67329), .ZN(
        n65452) );
  OAI22_X1 U46737 ( .A1(n63314), .A2(n67335), .B1(n63044), .B2(n67329), .ZN(
        n65434) );
  OAI22_X1 U46738 ( .A1(n63313), .A2(n67336), .B1(n63043), .B2(n67330), .ZN(
        n65416) );
  OAI22_X1 U46739 ( .A1(n63312), .A2(n67336), .B1(n63042), .B2(n67330), .ZN(
        n65398) );
  OAI22_X1 U46740 ( .A1(n63311), .A2(n67336), .B1(n63041), .B2(n67330), .ZN(
        n65380) );
  OAI22_X1 U46741 ( .A1(n63310), .A2(n67336), .B1(n63040), .B2(n67330), .ZN(
        n65362) );
  OAI22_X1 U46742 ( .A1(n63309), .A2(n67336), .B1(n63039), .B2(n67330), .ZN(
        n65344) );
  OAI22_X1 U46743 ( .A1(n63308), .A2(n67336), .B1(n63038), .B2(n67330), .ZN(
        n65326) );
  OAI22_X1 U46744 ( .A1(n63307), .A2(n67336), .B1(n63037), .B2(n67330), .ZN(
        n65308) );
  OAI22_X1 U46745 ( .A1(n63306), .A2(n67336), .B1(n63036), .B2(n67330), .ZN(
        n65290) );
  OAI22_X1 U46746 ( .A1(n63305), .A2(n67336), .B1(n63035), .B2(n67330), .ZN(
        n65272) );
  OAI22_X1 U46747 ( .A1(n63304), .A2(n67336), .B1(n63034), .B2(n67330), .ZN(
        n65254) );
  OAI22_X1 U46748 ( .A1(n63303), .A2(n67336), .B1(n63033), .B2(n67330), .ZN(
        n65236) );
  OAI22_X1 U46749 ( .A1(n63302), .A2(n67336), .B1(n63032), .B2(n67330), .ZN(
        n65218) );
  OAI22_X1 U46750 ( .A1(n63024), .A2(n67530), .B1(n62624), .B2(n67524), .ZN(
        n65090) );
  OAI22_X1 U46751 ( .A1(n63023), .A2(n67530), .B1(n62623), .B2(n67524), .ZN(
        n65058) );
  OAI22_X1 U46752 ( .A1(n63022), .A2(n67530), .B1(n62622), .B2(n67524), .ZN(
        n65038) );
  OAI22_X1 U46753 ( .A1(n63021), .A2(n67530), .B1(n62621), .B2(n67524), .ZN(
        n65018) );
  OAI22_X1 U46754 ( .A1(n63020), .A2(n67530), .B1(n62620), .B2(n67524), .ZN(
        n64998) );
  OAI22_X1 U46755 ( .A1(n63019), .A2(n67530), .B1(n62619), .B2(n67524), .ZN(
        n64978) );
  OAI22_X1 U46756 ( .A1(n63018), .A2(n67530), .B1(n62618), .B2(n67524), .ZN(
        n64958) );
  OAI22_X1 U46757 ( .A1(n63017), .A2(n67530), .B1(n62617), .B2(n67524), .ZN(
        n64938) );
  OAI22_X1 U46758 ( .A1(n63016), .A2(n67530), .B1(n62616), .B2(n67524), .ZN(
        n64918) );
  OAI22_X1 U46759 ( .A1(n63015), .A2(n67530), .B1(n62615), .B2(n67524), .ZN(
        n64898) );
  OAI22_X1 U46760 ( .A1(n63014), .A2(n67530), .B1(n62614), .B2(n67524), .ZN(
        n64878) );
  OAI22_X1 U46761 ( .A1(n63013), .A2(n67530), .B1(n62613), .B2(n67524), .ZN(
        n64858) );
  OAI22_X1 U46762 ( .A1(n63012), .A2(n67531), .B1(n62612), .B2(n67525), .ZN(
        n64838) );
  OAI22_X1 U46763 ( .A1(n63011), .A2(n67531), .B1(n62611), .B2(n67525), .ZN(
        n64818) );
  OAI22_X1 U46764 ( .A1(n63010), .A2(n67531), .B1(n62610), .B2(n67525), .ZN(
        n64798) );
  OAI22_X1 U46765 ( .A1(n63009), .A2(n67531), .B1(n62609), .B2(n67525), .ZN(
        n64778) );
  OAI22_X1 U46766 ( .A1(n63008), .A2(n67531), .B1(n62608), .B2(n67525), .ZN(
        n64758) );
  OAI22_X1 U46767 ( .A1(n63007), .A2(n67531), .B1(n62607), .B2(n67525), .ZN(
        n64738) );
  OAI22_X1 U46768 ( .A1(n63006), .A2(n67531), .B1(n62606), .B2(n67525), .ZN(
        n64718) );
  OAI22_X1 U46769 ( .A1(n63005), .A2(n67531), .B1(n62605), .B2(n67525), .ZN(
        n64698) );
  OAI22_X1 U46770 ( .A1(n63004), .A2(n67531), .B1(n62604), .B2(n67525), .ZN(
        n64678) );
  OAI22_X1 U46771 ( .A1(n63003), .A2(n67531), .B1(n62603), .B2(n67525), .ZN(
        n64658) );
  OAI22_X1 U46772 ( .A1(n63002), .A2(n67531), .B1(n62602), .B2(n67525), .ZN(
        n64638) );
  OAI22_X1 U46773 ( .A1(n63001), .A2(n67531), .B1(n62601), .B2(n67525), .ZN(
        n64618) );
  OAI22_X1 U46774 ( .A1(n63000), .A2(n67532), .B1(n62600), .B2(n67526), .ZN(
        n64598) );
  OAI22_X1 U46775 ( .A1(n62999), .A2(n67532), .B1(n62599), .B2(n67526), .ZN(
        n64578) );
  OAI22_X1 U46776 ( .A1(n62998), .A2(n67532), .B1(n62598), .B2(n67526), .ZN(
        n64558) );
  OAI22_X1 U46777 ( .A1(n62997), .A2(n67532), .B1(n62597), .B2(n67526), .ZN(
        n64538) );
  OAI22_X1 U46778 ( .A1(n62996), .A2(n67532), .B1(n62596), .B2(n67526), .ZN(
        n64518) );
  OAI22_X1 U46779 ( .A1(n62995), .A2(n67532), .B1(n62595), .B2(n67526), .ZN(
        n64498) );
  OAI22_X1 U46780 ( .A1(n62994), .A2(n67532), .B1(n62594), .B2(n67526), .ZN(
        n64478) );
  OAI22_X1 U46781 ( .A1(n62993), .A2(n67532), .B1(n62593), .B2(n67526), .ZN(
        n64458) );
  OAI22_X1 U46782 ( .A1(n62992), .A2(n67532), .B1(n62592), .B2(n67526), .ZN(
        n64438) );
  OAI22_X1 U46783 ( .A1(n62991), .A2(n67532), .B1(n62591), .B2(n67526), .ZN(
        n64418) );
  OAI22_X1 U46784 ( .A1(n62990), .A2(n67532), .B1(n62590), .B2(n67526), .ZN(
        n64398) );
  OAI22_X1 U46785 ( .A1(n62989), .A2(n67532), .B1(n62589), .B2(n67526), .ZN(
        n64378) );
  OAI22_X1 U46786 ( .A1(n62988), .A2(n67533), .B1(n62588), .B2(n67527), .ZN(
        n64358) );
  OAI22_X1 U46787 ( .A1(n62987), .A2(n67533), .B1(n62587), .B2(n67527), .ZN(
        n64338) );
  OAI22_X1 U46788 ( .A1(n62986), .A2(n67533), .B1(n62586), .B2(n67527), .ZN(
        n64318) );
  OAI22_X1 U46789 ( .A1(n62985), .A2(n67533), .B1(n62585), .B2(n67527), .ZN(
        n64298) );
  OAI22_X1 U46790 ( .A1(n62984), .A2(n67533), .B1(n62584), .B2(n67527), .ZN(
        n64278) );
  OAI22_X1 U46791 ( .A1(n62983), .A2(n67533), .B1(n62583), .B2(n67527), .ZN(
        n64258) );
  OAI22_X1 U46792 ( .A1(n62982), .A2(n67533), .B1(n62582), .B2(n67527), .ZN(
        n64238) );
  OAI22_X1 U46793 ( .A1(n62981), .A2(n67533), .B1(n62581), .B2(n67527), .ZN(
        n64218) );
  OAI22_X1 U46794 ( .A1(n62980), .A2(n67533), .B1(n62580), .B2(n67527), .ZN(
        n64198) );
  OAI22_X1 U46795 ( .A1(n62979), .A2(n67533), .B1(n62579), .B2(n67527), .ZN(
        n64178) );
  OAI22_X1 U46796 ( .A1(n62978), .A2(n67533), .B1(n62578), .B2(n67527), .ZN(
        n64158) );
  OAI22_X1 U46797 ( .A1(n62977), .A2(n67533), .B1(n62577), .B2(n67527), .ZN(
        n64138) );
  OAI22_X1 U46798 ( .A1(n62976), .A2(n67534), .B1(n62576), .B2(n67528), .ZN(
        n64118) );
  OAI22_X1 U46799 ( .A1(n62975), .A2(n67534), .B1(n62575), .B2(n67528), .ZN(
        n64098) );
  OAI22_X1 U46800 ( .A1(n62974), .A2(n67534), .B1(n62574), .B2(n67528), .ZN(
        n64078) );
  OAI22_X1 U46801 ( .A1(n62973), .A2(n67534), .B1(n62573), .B2(n67528), .ZN(
        n64058) );
  OAI22_X1 U46802 ( .A1(n62972), .A2(n67534), .B1(n62572), .B2(n67528), .ZN(
        n64038) );
  OAI22_X1 U46803 ( .A1(n62971), .A2(n67534), .B1(n62571), .B2(n67528), .ZN(
        n64018) );
  OAI22_X1 U46804 ( .A1(n62970), .A2(n67534), .B1(n62570), .B2(n67528), .ZN(
        n63998) );
  OAI22_X1 U46805 ( .A1(n62969), .A2(n67534), .B1(n62569), .B2(n67528), .ZN(
        n63978) );
  OAI22_X1 U46806 ( .A1(n62968), .A2(n67534), .B1(n62568), .B2(n67528), .ZN(
        n63958) );
  OAI22_X1 U46807 ( .A1(n62967), .A2(n67534), .B1(n62567), .B2(n67528), .ZN(
        n63938) );
  OAI22_X1 U46808 ( .A1(n62966), .A2(n67534), .B1(n62566), .B2(n67528), .ZN(
        n63918) );
  OAI22_X1 U46809 ( .A1(n62965), .A2(n67534), .B1(n62565), .B2(n67528), .ZN(
        n63898) );
  NAND2_X1 U46810 ( .A1(n66277), .A2(n66279), .ZN(n65138) );
  NAND2_X1 U46811 ( .A1(n65082), .A2(n65074), .ZN(n63813) );
  BUF_X1 U46812 ( .A(n61966), .Z(n68239) );
  BUF_X1 U46813 ( .A(n61964), .Z(n68242) );
  BUF_X1 U46814 ( .A(n61962), .Z(n68245) );
  BUF_X1 U46815 ( .A(n61960), .Z(n68248) );
  BUF_X1 U46816 ( .A(n62086), .Z(n68059) );
  BUF_X1 U46817 ( .A(n62084), .Z(n68062) );
  BUF_X1 U46818 ( .A(n62082), .Z(n68065) );
  BUF_X1 U46819 ( .A(n62080), .Z(n68068) );
  BUF_X1 U46820 ( .A(n62078), .Z(n68071) );
  BUF_X1 U46821 ( .A(n62076), .Z(n68074) );
  BUF_X1 U46822 ( .A(n62074), .Z(n68077) );
  BUF_X1 U46823 ( .A(n62072), .Z(n68080) );
  BUF_X1 U46824 ( .A(n62070), .Z(n68083) );
  BUF_X1 U46825 ( .A(n62068), .Z(n68086) );
  BUF_X1 U46826 ( .A(n62066), .Z(n68089) );
  BUF_X1 U46827 ( .A(n62064), .Z(n68092) );
  BUF_X1 U46828 ( .A(n62062), .Z(n68095) );
  BUF_X1 U46829 ( .A(n62060), .Z(n68098) );
  BUF_X1 U46830 ( .A(n62058), .Z(n68101) );
  BUF_X1 U46831 ( .A(n62056), .Z(n68104) );
  BUF_X1 U46832 ( .A(n62054), .Z(n68107) );
  BUF_X1 U46833 ( .A(n62052), .Z(n68110) );
  BUF_X1 U46834 ( .A(n62050), .Z(n68113) );
  BUF_X1 U46835 ( .A(n62048), .Z(n68116) );
  BUF_X1 U46836 ( .A(n62046), .Z(n68119) );
  BUF_X1 U46837 ( .A(n62044), .Z(n68122) );
  BUF_X1 U46838 ( .A(n62042), .Z(n68125) );
  BUF_X1 U46839 ( .A(n62040), .Z(n68128) );
  BUF_X1 U46840 ( .A(n62038), .Z(n68131) );
  BUF_X1 U46841 ( .A(n62036), .Z(n68134) );
  BUF_X1 U46842 ( .A(n62034), .Z(n68137) );
  BUF_X1 U46843 ( .A(n62032), .Z(n68140) );
  BUF_X1 U46844 ( .A(n62030), .Z(n68143) );
  BUF_X1 U46845 ( .A(n62028), .Z(n68146) );
  BUF_X1 U46846 ( .A(n62026), .Z(n68149) );
  BUF_X1 U46847 ( .A(n62024), .Z(n68152) );
  BUF_X1 U46848 ( .A(n62022), .Z(n68155) );
  BUF_X1 U46849 ( .A(n62020), .Z(n68158) );
  BUF_X1 U46850 ( .A(n62018), .Z(n68161) );
  BUF_X1 U46851 ( .A(n62016), .Z(n68164) );
  BUF_X1 U46852 ( .A(n62014), .Z(n68167) );
  BUF_X1 U46853 ( .A(n62012), .Z(n68170) );
  BUF_X1 U46854 ( .A(n62010), .Z(n68173) );
  BUF_X1 U46855 ( .A(n62008), .Z(n68176) );
  BUF_X1 U46856 ( .A(n62006), .Z(n68179) );
  BUF_X1 U46857 ( .A(n62004), .Z(n68182) );
  BUF_X1 U46858 ( .A(n62002), .Z(n68185) );
  BUF_X1 U46859 ( .A(n62000), .Z(n68188) );
  BUF_X1 U46860 ( .A(n61998), .Z(n68191) );
  BUF_X1 U46861 ( .A(n61996), .Z(n68194) );
  BUF_X1 U46862 ( .A(n61994), .Z(n68197) );
  BUF_X1 U46863 ( .A(n61992), .Z(n68200) );
  BUF_X1 U46864 ( .A(n61990), .Z(n68203) );
  BUF_X1 U46865 ( .A(n61988), .Z(n68206) );
  BUF_X1 U46866 ( .A(n61986), .Z(n68209) );
  BUF_X1 U46867 ( .A(n61984), .Z(n68212) );
  BUF_X1 U46868 ( .A(n61982), .Z(n68215) );
  BUF_X1 U46869 ( .A(n61980), .Z(n68218) );
  BUF_X1 U46870 ( .A(n61978), .Z(n68221) );
  BUF_X1 U46871 ( .A(n61976), .Z(n68224) );
  BUF_X1 U46872 ( .A(n61974), .Z(n68227) );
  BUF_X1 U46873 ( .A(n61972), .Z(n68230) );
  BUF_X1 U46874 ( .A(n61970), .Z(n68233) );
  BUF_X1 U46875 ( .A(n61968), .Z(n68236) );
  BUF_X1 U46876 ( .A(n65112), .Z(n67438) );
  NAND2_X1 U46877 ( .A1(n65085), .A2(n65075), .ZN(n63786) );
  NAND2_X1 U46878 ( .A1(n65080), .A2(n65075), .ZN(n63818) );
  NAND2_X1 U46879 ( .A1(n65087), .A2(n65075), .ZN(n63819) );
  NAND2_X1 U46880 ( .A1(n66280), .A2(n66283), .ZN(n65113) );
  NAND2_X1 U46881 ( .A1(n65075), .A2(n65077), .ZN(n63802) );
  NAND2_X1 U46882 ( .A1(n65075), .A2(n65076), .ZN(n63776) );
  NAND2_X1 U46883 ( .A1(n65075), .A2(n65081), .ZN(n63781) );
  BUF_X1 U46884 ( .A(n61966), .Z(n68238) );
  BUF_X1 U46885 ( .A(n61964), .Z(n68241) );
  BUF_X1 U46886 ( .A(n61962), .Z(n68244) );
  BUF_X1 U46887 ( .A(n61960), .Z(n68247) );
  BUF_X1 U46888 ( .A(n62086), .Z(n68058) );
  BUF_X1 U46889 ( .A(n62084), .Z(n68061) );
  BUF_X1 U46890 ( .A(n62082), .Z(n68064) );
  BUF_X1 U46891 ( .A(n62080), .Z(n68067) );
  BUF_X1 U46892 ( .A(n62078), .Z(n68070) );
  BUF_X1 U46893 ( .A(n62076), .Z(n68073) );
  BUF_X1 U46894 ( .A(n62074), .Z(n68076) );
  BUF_X1 U46895 ( .A(n62072), .Z(n68079) );
  BUF_X1 U46896 ( .A(n62070), .Z(n68082) );
  BUF_X1 U46897 ( .A(n62068), .Z(n68085) );
  BUF_X1 U46898 ( .A(n62066), .Z(n68088) );
  BUF_X1 U46899 ( .A(n62064), .Z(n68091) );
  BUF_X1 U46900 ( .A(n62062), .Z(n68094) );
  BUF_X1 U46901 ( .A(n62060), .Z(n68097) );
  BUF_X1 U46902 ( .A(n62058), .Z(n68100) );
  BUF_X1 U46903 ( .A(n62056), .Z(n68103) );
  BUF_X1 U46904 ( .A(n62054), .Z(n68106) );
  BUF_X1 U46905 ( .A(n62052), .Z(n68109) );
  BUF_X1 U46906 ( .A(n62050), .Z(n68112) );
  BUF_X1 U46907 ( .A(n62048), .Z(n68115) );
  BUF_X1 U46908 ( .A(n62046), .Z(n68118) );
  BUF_X1 U46909 ( .A(n62044), .Z(n68121) );
  BUF_X1 U46910 ( .A(n62042), .Z(n68124) );
  BUF_X1 U46911 ( .A(n62040), .Z(n68127) );
  BUF_X1 U46912 ( .A(n62038), .Z(n68130) );
  BUF_X1 U46913 ( .A(n62036), .Z(n68133) );
  BUF_X1 U46914 ( .A(n62034), .Z(n68136) );
  BUF_X1 U46915 ( .A(n62032), .Z(n68139) );
  BUF_X1 U46916 ( .A(n62030), .Z(n68142) );
  BUF_X1 U46917 ( .A(n62028), .Z(n68145) );
  BUF_X1 U46918 ( .A(n62026), .Z(n68148) );
  BUF_X1 U46919 ( .A(n62024), .Z(n68151) );
  BUF_X1 U46920 ( .A(n62022), .Z(n68154) );
  BUF_X1 U46921 ( .A(n62020), .Z(n68157) );
  BUF_X1 U46922 ( .A(n62018), .Z(n68160) );
  BUF_X1 U46923 ( .A(n62016), .Z(n68163) );
  BUF_X1 U46924 ( .A(n62014), .Z(n68166) );
  BUF_X1 U46925 ( .A(n62012), .Z(n68169) );
  BUF_X1 U46926 ( .A(n62010), .Z(n68172) );
  BUF_X1 U46927 ( .A(n62008), .Z(n68175) );
  BUF_X1 U46928 ( .A(n62006), .Z(n68178) );
  BUF_X1 U46929 ( .A(n62004), .Z(n68181) );
  BUF_X1 U46930 ( .A(n62002), .Z(n68184) );
  BUF_X1 U46931 ( .A(n62000), .Z(n68187) );
  BUF_X1 U46932 ( .A(n61998), .Z(n68190) );
  BUF_X1 U46933 ( .A(n61996), .Z(n68193) );
  BUF_X1 U46934 ( .A(n61994), .Z(n68196) );
  BUF_X1 U46935 ( .A(n61992), .Z(n68199) );
  BUF_X1 U46936 ( .A(n61990), .Z(n68202) );
  BUF_X1 U46937 ( .A(n61988), .Z(n68205) );
  BUF_X1 U46938 ( .A(n61986), .Z(n68208) );
  BUF_X1 U46939 ( .A(n61984), .Z(n68211) );
  BUF_X1 U46940 ( .A(n61982), .Z(n68214) );
  BUF_X1 U46941 ( .A(n61980), .Z(n68217) );
  BUF_X1 U46942 ( .A(n61978), .Z(n68220) );
  BUF_X1 U46943 ( .A(n61976), .Z(n68223) );
  BUF_X1 U46944 ( .A(n61974), .Z(n68226) );
  BUF_X1 U46945 ( .A(n61972), .Z(n68229) );
  BUF_X1 U46946 ( .A(n61970), .Z(n68232) );
  BUF_X1 U46947 ( .A(n61968), .Z(n68235) );
  OAI22_X1 U46948 ( .A1(n67934), .A2(n62694), .B1(n68247), .B2(n67928), .ZN(
        n6846) );
  NAND2_X1 U46949 ( .A1(n65077), .A2(n65078), .ZN(n63775) );
  OAI22_X1 U46950 ( .A1(n67947), .A2(n62631), .B1(n68238), .B2(n67940), .ZN(
        n6907) );
  OAI22_X1 U46951 ( .A1(n67947), .A2(n62630), .B1(n68241), .B2(n67940), .ZN(
        n6908) );
  OAI22_X1 U46952 ( .A1(n67947), .A2(n62629), .B1(n68244), .B2(n67940), .ZN(
        n6909) );
  OAI22_X1 U46953 ( .A1(n67947), .A2(n62627), .B1(n68247), .B2(n67940), .ZN(
        n6910) );
  OAI22_X1 U46954 ( .A1(n67960), .A2(n62564), .B1(n68238), .B2(n67953), .ZN(
        n6971) );
  OAI22_X1 U46955 ( .A1(n67960), .A2(n62563), .B1(n68241), .B2(n67953), .ZN(
        n6972) );
  OAI22_X1 U46956 ( .A1(n67960), .A2(n62562), .B1(n68244), .B2(n67953), .ZN(
        n6973) );
  OAI22_X1 U46957 ( .A1(n67960), .A2(n62560), .B1(n68247), .B2(n67953), .ZN(
        n6974) );
  OAI22_X1 U46958 ( .A1(n68051), .A2(n62095), .B1(n68238), .B2(n68044), .ZN(
        n7419) );
  OAI22_X1 U46959 ( .A1(n68051), .A2(n62094), .B1(n68241), .B2(n68044), .ZN(
        n7420) );
  OAI22_X1 U46960 ( .A1(n68051), .A2(n62093), .B1(n68244), .B2(n68044), .ZN(
        n7421) );
  OAI22_X1 U46961 ( .A1(n68051), .A2(n62091), .B1(n68247), .B2(n68044), .ZN(
        n7422) );
  OAI22_X1 U46962 ( .A1(n68012), .A2(n62295), .B1(n68238), .B2(n68005), .ZN(
        n7227) );
  OAI22_X1 U46963 ( .A1(n68012), .A2(n62294), .B1(n68241), .B2(n68005), .ZN(
        n7228) );
  OAI22_X1 U46964 ( .A1(n68012), .A2(n62293), .B1(n68244), .B2(n68005), .ZN(
        n7229) );
  OAI22_X1 U46965 ( .A1(n68012), .A2(n62291), .B1(n68247), .B2(n68005), .ZN(
        n7230) );
  OAI22_X1 U46966 ( .A1(n67973), .A2(n62498), .B1(n68238), .B2(n67966), .ZN(
        n7035) );
  OAI22_X1 U46967 ( .A1(n67973), .A2(n62497), .B1(n68241), .B2(n67966), .ZN(
        n7036) );
  OAI22_X1 U46968 ( .A1(n67973), .A2(n62496), .B1(n68244), .B2(n67966), .ZN(
        n7037) );
  OAI22_X1 U46969 ( .A1(n67973), .A2(n62494), .B1(n68247), .B2(n67966), .ZN(
        n7038) );
  OAI22_X1 U46970 ( .A1(n67807), .A2(n63166), .B1(n68239), .B2(n67800), .ZN(
        n6203) );
  OAI22_X1 U46971 ( .A1(n67807), .A2(n63165), .B1(n68242), .B2(n67800), .ZN(
        n6204) );
  OAI22_X1 U46972 ( .A1(n67807), .A2(n63164), .B1(n68245), .B2(n67800), .ZN(
        n6205) );
  OAI22_X1 U46973 ( .A1(n67807), .A2(n63162), .B1(n68248), .B2(n67800), .ZN(
        n6206) );
  OAI22_X1 U46974 ( .A1(n67858), .A2(n62964), .B1(n68239), .B2(n67851), .ZN(
        n6459) );
  OAI22_X1 U46975 ( .A1(n67858), .A2(n62963), .B1(n68242), .B2(n67851), .ZN(
        n6460) );
  OAI22_X1 U46976 ( .A1(n67858), .A2(n62962), .B1(n68245), .B2(n67851), .ZN(
        n6461) );
  OAI22_X1 U46977 ( .A1(n67858), .A2(n62960), .B1(n68248), .B2(n67851), .ZN(
        n6462) );
  OAI22_X1 U46978 ( .A1(n67845), .A2(n63031), .B1(n68239), .B2(n67838), .ZN(
        n6395) );
  OAI22_X1 U46979 ( .A1(n67845), .A2(n63030), .B1(n68242), .B2(n67838), .ZN(
        n6396) );
  OAI22_X1 U46980 ( .A1(n67845), .A2(n63029), .B1(n68245), .B2(n67838), .ZN(
        n6397) );
  OAI22_X1 U46981 ( .A1(n67845), .A2(n63027), .B1(n68248), .B2(n67838), .ZN(
        n6398) );
  OAI22_X1 U46982 ( .A1(n67756), .A2(n63367), .B1(n68239), .B2(n67749), .ZN(
        n5947) );
  OAI22_X1 U46983 ( .A1(n67756), .A2(n63366), .B1(n68242), .B2(n67749), .ZN(
        n5948) );
  OAI22_X1 U46984 ( .A1(n67756), .A2(n63365), .B1(n68245), .B2(n67749), .ZN(
        n5949) );
  OAI22_X1 U46985 ( .A1(n67756), .A2(n63363), .B1(n68248), .B2(n67749), .ZN(
        n5950) );
  OAI22_X1 U46986 ( .A1(n67743), .A2(n63434), .B1(n68240), .B2(n67736), .ZN(
        n5883) );
  OAI22_X1 U46987 ( .A1(n67743), .A2(n63433), .B1(n68243), .B2(n67736), .ZN(
        n5884) );
  OAI22_X1 U46988 ( .A1(n67743), .A2(n63432), .B1(n68246), .B2(n67736), .ZN(
        n5885) );
  OAI22_X1 U46989 ( .A1(n67743), .A2(n63430), .B1(n68249), .B2(n67736), .ZN(
        n5886) );
  OAI22_X1 U46990 ( .A1(n67884), .A2(n62831), .B1(n68239), .B2(n67877), .ZN(
        n6587) );
  OAI22_X1 U46991 ( .A1(n67884), .A2(n62830), .B1(n68242), .B2(n67877), .ZN(
        n6588) );
  OAI22_X1 U46992 ( .A1(n67884), .A2(n62829), .B1(n68245), .B2(n67877), .ZN(
        n6589) );
  OAI22_X1 U46993 ( .A1(n67884), .A2(n62827), .B1(n68248), .B2(n67877), .ZN(
        n6590) );
  OAI22_X1 U46994 ( .A1(n68038), .A2(n62162), .B1(n68238), .B2(n68031), .ZN(
        n7355) );
  OAI22_X1 U46995 ( .A1(n68038), .A2(n62161), .B1(n68241), .B2(n68031), .ZN(
        n7356) );
  OAI22_X1 U46996 ( .A1(n68038), .A2(n62160), .B1(n68244), .B2(n68031), .ZN(
        n7357) );
  OAI22_X1 U46997 ( .A1(n68038), .A2(n62158), .B1(n68247), .B2(n68031), .ZN(
        n7358) );
  OAI22_X1 U46998 ( .A1(n68025), .A2(n62229), .B1(n68238), .B2(n68018), .ZN(
        n7291) );
  OAI22_X1 U46999 ( .A1(n68025), .A2(n62228), .B1(n68241), .B2(n68018), .ZN(
        n7292) );
  OAI22_X1 U47000 ( .A1(n68025), .A2(n62227), .B1(n68244), .B2(n68018), .ZN(
        n7293) );
  OAI22_X1 U47001 ( .A1(n68025), .A2(n62225), .B1(n68247), .B2(n68018), .ZN(
        n7294) );
  OAI22_X1 U47002 ( .A1(n67999), .A2(n62362), .B1(n68238), .B2(n67992), .ZN(
        n7163) );
  OAI22_X1 U47003 ( .A1(n67999), .A2(n62361), .B1(n68241), .B2(n67992), .ZN(
        n7164) );
  OAI22_X1 U47004 ( .A1(n67999), .A2(n62360), .B1(n68244), .B2(n67992), .ZN(
        n7165) );
  OAI22_X1 U47005 ( .A1(n67999), .A2(n62358), .B1(n68247), .B2(n67992), .ZN(
        n7166) );
  OAI22_X1 U47006 ( .A1(n67820), .A2(n63100), .B1(n68239), .B2(n67813), .ZN(
        n6267) );
  OAI22_X1 U47007 ( .A1(n67820), .A2(n63099), .B1(n68242), .B2(n67813), .ZN(
        n6268) );
  OAI22_X1 U47008 ( .A1(n67820), .A2(n63098), .B1(n68245), .B2(n67813), .ZN(
        n6269) );
  OAI22_X1 U47009 ( .A1(n67820), .A2(n63096), .B1(n68248), .B2(n67813), .ZN(
        n6270) );
  OAI22_X1 U47010 ( .A1(n67692), .A2(n63637), .B1(n68240), .B2(n67685), .ZN(
        n5627) );
  OAI22_X1 U47011 ( .A1(n67692), .A2(n63636), .B1(n68243), .B2(n67685), .ZN(
        n5628) );
  OAI22_X1 U47012 ( .A1(n67692), .A2(n63635), .B1(n68246), .B2(n67685), .ZN(
        n5629) );
  OAI22_X1 U47013 ( .A1(n67692), .A2(n63633), .B1(n68249), .B2(n67685), .ZN(
        n5630) );
  OAI22_X1 U47014 ( .A1(n67871), .A2(n62897), .B1(n68239), .B2(n67864), .ZN(
        n6523) );
  OAI22_X1 U47015 ( .A1(n67871), .A2(n62896), .B1(n68242), .B2(n67864), .ZN(
        n6524) );
  OAI22_X1 U47016 ( .A1(n67871), .A2(n62895), .B1(n68245), .B2(n67864), .ZN(
        n6525) );
  OAI22_X1 U47017 ( .A1(n67871), .A2(n62893), .B1(n68248), .B2(n67864), .ZN(
        n6526) );
  OAI22_X1 U47018 ( .A1(n67922), .A2(n62701), .B1(n68238), .B2(n67915), .ZN(
        n6779) );
  OAI22_X1 U47019 ( .A1(n67922), .A2(n62700), .B1(n68241), .B2(n67915), .ZN(
        n6780) );
  OAI22_X1 U47020 ( .A1(n67922), .A2(n62699), .B1(n68244), .B2(n67915), .ZN(
        n6781) );
  OAI22_X1 U47021 ( .A1(n67922), .A2(n62697), .B1(n68247), .B2(n67915), .ZN(
        n6782) );
  OAI22_X1 U47022 ( .A1(n67986), .A2(n62428), .B1(n68238), .B2(n67979), .ZN(
        n7099) );
  OAI22_X1 U47023 ( .A1(n67986), .A2(n62427), .B1(n68241), .B2(n67979), .ZN(
        n7100) );
  OAI22_X1 U47024 ( .A1(n67986), .A2(n62426), .B1(n68244), .B2(n67979), .ZN(
        n7101) );
  OAI22_X1 U47025 ( .A1(n67986), .A2(n62424), .B1(n68247), .B2(n67979), .ZN(
        n7102) );
  OAI22_X1 U47026 ( .A1(n67769), .A2(n63301), .B1(n68239), .B2(n67762), .ZN(
        n6011) );
  OAI22_X1 U47027 ( .A1(n67769), .A2(n63300), .B1(n68242), .B2(n67762), .ZN(
        n6012) );
  OAI22_X1 U47028 ( .A1(n67769), .A2(n63299), .B1(n68245), .B2(n67762), .ZN(
        n6013) );
  OAI22_X1 U47029 ( .A1(n67769), .A2(n63297), .B1(n68248), .B2(n67762), .ZN(
        n6014) );
  OAI22_X1 U47030 ( .A1(n67718), .A2(n63505), .B1(n68240), .B2(n67711), .ZN(
        n5755) );
  OAI22_X1 U47031 ( .A1(n67718), .A2(n63504), .B1(n68243), .B2(n67711), .ZN(
        n5756) );
  OAI22_X1 U47032 ( .A1(n67718), .A2(n63503), .B1(n68246), .B2(n67711), .ZN(
        n5757) );
  OAI22_X1 U47033 ( .A1(n67718), .A2(n63501), .B1(n68249), .B2(n67711), .ZN(
        n5758) );
  OAI22_X1 U47034 ( .A1(n67705), .A2(n63571), .B1(n68240), .B2(n67698), .ZN(
        n5691) );
  OAI22_X1 U47035 ( .A1(n67705), .A2(n63570), .B1(n68243), .B2(n67698), .ZN(
        n5692) );
  OAI22_X1 U47036 ( .A1(n67705), .A2(n63569), .B1(n68246), .B2(n67698), .ZN(
        n5693) );
  OAI22_X1 U47037 ( .A1(n67705), .A2(n63567), .B1(n68249), .B2(n67698), .ZN(
        n5694) );
  NAND2_X1 U47038 ( .A1(n66280), .A2(n66278), .ZN(n65123) );
  OAI22_X1 U47039 ( .A1(n67739), .A2(n63494), .B1(n68060), .B2(n67731), .ZN(
        n5823) );
  OAI22_X1 U47040 ( .A1(n67739), .A2(n63493), .B1(n68063), .B2(n67731), .ZN(
        n5824) );
  OAI22_X1 U47041 ( .A1(n67739), .A2(n63492), .B1(n68066), .B2(n67731), .ZN(
        n5825) );
  OAI22_X1 U47042 ( .A1(n67739), .A2(n63491), .B1(n68069), .B2(n67731), .ZN(
        n5826) );
  OAI22_X1 U47043 ( .A1(n67739), .A2(n63490), .B1(n68072), .B2(n67731), .ZN(
        n5827) );
  OAI22_X1 U47044 ( .A1(n67739), .A2(n63489), .B1(n68075), .B2(n67731), .ZN(
        n5828) );
  OAI22_X1 U47045 ( .A1(n67739), .A2(n63488), .B1(n68078), .B2(n67731), .ZN(
        n5829) );
  OAI22_X1 U47046 ( .A1(n67739), .A2(n63487), .B1(n68081), .B2(n67731), .ZN(
        n5830) );
  OAI22_X1 U47047 ( .A1(n67739), .A2(n63486), .B1(n68084), .B2(n67731), .ZN(
        n5831) );
  OAI22_X1 U47048 ( .A1(n67739), .A2(n63485), .B1(n68087), .B2(n67731), .ZN(
        n5832) );
  OAI22_X1 U47049 ( .A1(n67739), .A2(n63484), .B1(n68090), .B2(n67731), .ZN(
        n5833) );
  OAI22_X1 U47050 ( .A1(n67739), .A2(n63483), .B1(n68093), .B2(n67731), .ZN(
        n5834) );
  OAI22_X1 U47051 ( .A1(n67740), .A2(n63482), .B1(n68096), .B2(n67732), .ZN(
        n5835) );
  OAI22_X1 U47052 ( .A1(n67740), .A2(n63481), .B1(n68099), .B2(n67732), .ZN(
        n5836) );
  OAI22_X1 U47053 ( .A1(n67740), .A2(n63480), .B1(n68102), .B2(n67732), .ZN(
        n5837) );
  OAI22_X1 U47054 ( .A1(n67740), .A2(n63479), .B1(n68105), .B2(n67732), .ZN(
        n5838) );
  OAI22_X1 U47055 ( .A1(n67740), .A2(n63478), .B1(n68108), .B2(n67732), .ZN(
        n5839) );
  OAI22_X1 U47056 ( .A1(n67740), .A2(n63477), .B1(n68111), .B2(n67732), .ZN(
        n5840) );
  OAI22_X1 U47057 ( .A1(n67740), .A2(n63476), .B1(n68114), .B2(n67732), .ZN(
        n5841) );
  OAI22_X1 U47058 ( .A1(n67740), .A2(n63475), .B1(n68117), .B2(n67732), .ZN(
        n5842) );
  OAI22_X1 U47059 ( .A1(n67740), .A2(n63474), .B1(n68120), .B2(n67732), .ZN(
        n5843) );
  OAI22_X1 U47060 ( .A1(n67740), .A2(n63473), .B1(n68123), .B2(n67732), .ZN(
        n5844) );
  OAI22_X1 U47061 ( .A1(n67740), .A2(n63472), .B1(n68126), .B2(n67732), .ZN(
        n5845) );
  OAI22_X1 U47062 ( .A1(n67740), .A2(n63471), .B1(n68129), .B2(n67732), .ZN(
        n5846) );
  OAI22_X1 U47063 ( .A1(n67740), .A2(n63470), .B1(n68132), .B2(n67733), .ZN(
        n5847) );
  OAI22_X1 U47064 ( .A1(n67741), .A2(n63469), .B1(n68135), .B2(n67733), .ZN(
        n5848) );
  OAI22_X1 U47065 ( .A1(n67741), .A2(n63468), .B1(n68138), .B2(n67733), .ZN(
        n5849) );
  OAI22_X1 U47066 ( .A1(n67741), .A2(n63467), .B1(n68141), .B2(n67733), .ZN(
        n5850) );
  OAI22_X1 U47067 ( .A1(n67741), .A2(n63466), .B1(n68144), .B2(n67733), .ZN(
        n5851) );
  OAI22_X1 U47068 ( .A1(n67741), .A2(n63465), .B1(n68147), .B2(n67733), .ZN(
        n5852) );
  OAI22_X1 U47069 ( .A1(n67741), .A2(n63464), .B1(n68150), .B2(n67733), .ZN(
        n5853) );
  OAI22_X1 U47070 ( .A1(n67741), .A2(n63463), .B1(n68153), .B2(n67733), .ZN(
        n5854) );
  OAI22_X1 U47071 ( .A1(n67741), .A2(n63462), .B1(n68156), .B2(n67733), .ZN(
        n5855) );
  OAI22_X1 U47072 ( .A1(n67741), .A2(n63461), .B1(n68159), .B2(n67733), .ZN(
        n5856) );
  OAI22_X1 U47073 ( .A1(n67741), .A2(n63460), .B1(n68162), .B2(n67733), .ZN(
        n5857) );
  OAI22_X1 U47074 ( .A1(n67741), .A2(n63459), .B1(n68165), .B2(n67733), .ZN(
        n5858) );
  OAI22_X1 U47075 ( .A1(n67741), .A2(n63458), .B1(n68168), .B2(n67734), .ZN(
        n5859) );
  OAI22_X1 U47076 ( .A1(n67741), .A2(n63457), .B1(n68171), .B2(n67734), .ZN(
        n5860) );
  OAI22_X1 U47077 ( .A1(n67742), .A2(n63456), .B1(n68174), .B2(n67734), .ZN(
        n5861) );
  OAI22_X1 U47078 ( .A1(n67742), .A2(n63455), .B1(n68177), .B2(n67734), .ZN(
        n5862) );
  OAI22_X1 U47079 ( .A1(n67742), .A2(n63454), .B1(n68180), .B2(n67734), .ZN(
        n5863) );
  OAI22_X1 U47080 ( .A1(n67742), .A2(n63453), .B1(n68183), .B2(n67734), .ZN(
        n5864) );
  OAI22_X1 U47081 ( .A1(n67742), .A2(n63452), .B1(n68186), .B2(n67734), .ZN(
        n5865) );
  OAI22_X1 U47082 ( .A1(n67742), .A2(n63451), .B1(n68189), .B2(n67734), .ZN(
        n5866) );
  OAI22_X1 U47083 ( .A1(n67742), .A2(n63450), .B1(n68192), .B2(n67734), .ZN(
        n5867) );
  OAI22_X1 U47084 ( .A1(n67742), .A2(n63449), .B1(n68195), .B2(n67734), .ZN(
        n5868) );
  OAI22_X1 U47085 ( .A1(n67742), .A2(n63448), .B1(n68198), .B2(n67734), .ZN(
        n5869) );
  OAI22_X1 U47086 ( .A1(n67742), .A2(n63447), .B1(n68201), .B2(n67734), .ZN(
        n5870) );
  OAI22_X1 U47087 ( .A1(n67742), .A2(n63446), .B1(n68204), .B2(n67735), .ZN(
        n5871) );
  OAI22_X1 U47088 ( .A1(n67742), .A2(n63445), .B1(n68207), .B2(n67735), .ZN(
        n5872) );
  OAI22_X1 U47089 ( .A1(n67742), .A2(n63444), .B1(n68210), .B2(n67735), .ZN(
        n5873) );
  OAI22_X1 U47090 ( .A1(n67743), .A2(n63443), .B1(n68213), .B2(n67735), .ZN(
        n5874) );
  OAI22_X1 U47091 ( .A1(n67743), .A2(n63442), .B1(n68216), .B2(n67735), .ZN(
        n5875) );
  OAI22_X1 U47092 ( .A1(n67743), .A2(n63441), .B1(n68219), .B2(n67735), .ZN(
        n5876) );
  OAI22_X1 U47093 ( .A1(n67743), .A2(n63440), .B1(n68222), .B2(n67735), .ZN(
        n5877) );
  OAI22_X1 U47094 ( .A1(n67743), .A2(n63439), .B1(n68225), .B2(n67735), .ZN(
        n5878) );
  OAI22_X1 U47095 ( .A1(n67743), .A2(n63438), .B1(n68228), .B2(n67735), .ZN(
        n5879) );
  OAI22_X1 U47096 ( .A1(n67743), .A2(n63437), .B1(n68231), .B2(n67735), .ZN(
        n5880) );
  OAI22_X1 U47097 ( .A1(n67743), .A2(n63436), .B1(n68234), .B2(n67735), .ZN(
        n5881) );
  OAI22_X1 U47098 ( .A1(n67743), .A2(n63435), .B1(n68237), .B2(n67735), .ZN(
        n5882) );
  OAI22_X1 U47099 ( .A1(n67688), .A2(n63697), .B1(n68060), .B2(n67680), .ZN(
        n5567) );
  OAI22_X1 U47100 ( .A1(n67688), .A2(n63696), .B1(n68063), .B2(n67680), .ZN(
        n5568) );
  OAI22_X1 U47101 ( .A1(n67688), .A2(n63695), .B1(n68066), .B2(n67680), .ZN(
        n5569) );
  OAI22_X1 U47102 ( .A1(n67688), .A2(n63694), .B1(n68069), .B2(n67680), .ZN(
        n5570) );
  OAI22_X1 U47103 ( .A1(n67688), .A2(n63693), .B1(n68072), .B2(n67680), .ZN(
        n5571) );
  OAI22_X1 U47104 ( .A1(n67688), .A2(n63692), .B1(n68075), .B2(n67680), .ZN(
        n5572) );
  OAI22_X1 U47105 ( .A1(n67688), .A2(n63691), .B1(n68078), .B2(n67680), .ZN(
        n5573) );
  OAI22_X1 U47106 ( .A1(n67688), .A2(n63690), .B1(n68081), .B2(n67680), .ZN(
        n5574) );
  OAI22_X1 U47107 ( .A1(n67688), .A2(n63689), .B1(n68084), .B2(n67680), .ZN(
        n5575) );
  OAI22_X1 U47108 ( .A1(n67688), .A2(n63688), .B1(n68087), .B2(n67680), .ZN(
        n5576) );
  OAI22_X1 U47109 ( .A1(n67688), .A2(n63687), .B1(n68090), .B2(n67680), .ZN(
        n5577) );
  OAI22_X1 U47110 ( .A1(n67688), .A2(n63686), .B1(n68093), .B2(n67680), .ZN(
        n5578) );
  OAI22_X1 U47111 ( .A1(n67689), .A2(n63685), .B1(n68096), .B2(n67681), .ZN(
        n5579) );
  OAI22_X1 U47112 ( .A1(n67689), .A2(n63684), .B1(n68099), .B2(n67681), .ZN(
        n5580) );
  OAI22_X1 U47113 ( .A1(n67689), .A2(n63683), .B1(n68102), .B2(n67681), .ZN(
        n5581) );
  OAI22_X1 U47114 ( .A1(n67689), .A2(n63682), .B1(n68105), .B2(n67681), .ZN(
        n5582) );
  OAI22_X1 U47115 ( .A1(n67689), .A2(n63681), .B1(n68108), .B2(n67681), .ZN(
        n5583) );
  OAI22_X1 U47116 ( .A1(n67689), .A2(n63680), .B1(n68111), .B2(n67681), .ZN(
        n5584) );
  OAI22_X1 U47117 ( .A1(n67689), .A2(n63679), .B1(n68114), .B2(n67681), .ZN(
        n5585) );
  OAI22_X1 U47118 ( .A1(n67689), .A2(n63678), .B1(n68117), .B2(n67681), .ZN(
        n5586) );
  OAI22_X1 U47119 ( .A1(n67689), .A2(n63677), .B1(n68120), .B2(n67681), .ZN(
        n5587) );
  OAI22_X1 U47120 ( .A1(n67689), .A2(n63676), .B1(n68123), .B2(n67681), .ZN(
        n5588) );
  OAI22_X1 U47121 ( .A1(n67689), .A2(n63675), .B1(n68126), .B2(n67681), .ZN(
        n5589) );
  OAI22_X1 U47122 ( .A1(n67689), .A2(n63674), .B1(n68129), .B2(n67681), .ZN(
        n5590) );
  OAI22_X1 U47123 ( .A1(n67689), .A2(n63673), .B1(n68132), .B2(n67682), .ZN(
        n5591) );
  OAI22_X1 U47124 ( .A1(n67690), .A2(n63672), .B1(n68135), .B2(n67682), .ZN(
        n5592) );
  OAI22_X1 U47125 ( .A1(n67690), .A2(n63671), .B1(n68138), .B2(n67682), .ZN(
        n5593) );
  OAI22_X1 U47126 ( .A1(n67690), .A2(n63670), .B1(n68141), .B2(n67682), .ZN(
        n5594) );
  OAI22_X1 U47127 ( .A1(n67690), .A2(n63669), .B1(n68144), .B2(n67682), .ZN(
        n5595) );
  OAI22_X1 U47128 ( .A1(n67690), .A2(n63668), .B1(n68147), .B2(n67682), .ZN(
        n5596) );
  OAI22_X1 U47129 ( .A1(n67690), .A2(n63667), .B1(n68150), .B2(n67682), .ZN(
        n5597) );
  OAI22_X1 U47130 ( .A1(n67690), .A2(n63666), .B1(n68153), .B2(n67682), .ZN(
        n5598) );
  OAI22_X1 U47131 ( .A1(n67690), .A2(n63665), .B1(n68156), .B2(n67682), .ZN(
        n5599) );
  OAI22_X1 U47132 ( .A1(n67690), .A2(n63664), .B1(n68159), .B2(n67682), .ZN(
        n5600) );
  OAI22_X1 U47133 ( .A1(n67690), .A2(n63663), .B1(n68162), .B2(n67682), .ZN(
        n5601) );
  OAI22_X1 U47134 ( .A1(n67690), .A2(n63662), .B1(n68165), .B2(n67682), .ZN(
        n5602) );
  OAI22_X1 U47135 ( .A1(n67690), .A2(n63661), .B1(n68168), .B2(n67683), .ZN(
        n5603) );
  OAI22_X1 U47136 ( .A1(n67690), .A2(n63660), .B1(n68171), .B2(n67683), .ZN(
        n5604) );
  OAI22_X1 U47137 ( .A1(n67691), .A2(n63659), .B1(n68174), .B2(n67683), .ZN(
        n5605) );
  OAI22_X1 U47138 ( .A1(n67691), .A2(n63658), .B1(n68177), .B2(n67683), .ZN(
        n5606) );
  OAI22_X1 U47139 ( .A1(n67691), .A2(n63657), .B1(n68180), .B2(n67683), .ZN(
        n5607) );
  OAI22_X1 U47140 ( .A1(n67691), .A2(n63656), .B1(n68183), .B2(n67683), .ZN(
        n5608) );
  OAI22_X1 U47141 ( .A1(n67691), .A2(n63655), .B1(n68186), .B2(n67683), .ZN(
        n5609) );
  OAI22_X1 U47142 ( .A1(n67691), .A2(n63654), .B1(n68189), .B2(n67683), .ZN(
        n5610) );
  OAI22_X1 U47143 ( .A1(n67691), .A2(n63653), .B1(n68192), .B2(n67683), .ZN(
        n5611) );
  OAI22_X1 U47144 ( .A1(n67691), .A2(n63652), .B1(n68195), .B2(n67683), .ZN(
        n5612) );
  OAI22_X1 U47145 ( .A1(n67691), .A2(n63651), .B1(n68198), .B2(n67683), .ZN(
        n5613) );
  OAI22_X1 U47146 ( .A1(n67691), .A2(n63650), .B1(n68201), .B2(n67683), .ZN(
        n5614) );
  OAI22_X1 U47147 ( .A1(n67691), .A2(n63649), .B1(n68204), .B2(n67684), .ZN(
        n5615) );
  OAI22_X1 U47148 ( .A1(n67691), .A2(n63648), .B1(n68207), .B2(n67684), .ZN(
        n5616) );
  OAI22_X1 U47149 ( .A1(n67691), .A2(n63647), .B1(n68210), .B2(n67684), .ZN(
        n5617) );
  OAI22_X1 U47150 ( .A1(n67692), .A2(n63646), .B1(n68213), .B2(n67684), .ZN(
        n5618) );
  OAI22_X1 U47151 ( .A1(n67692), .A2(n63645), .B1(n68216), .B2(n67684), .ZN(
        n5619) );
  OAI22_X1 U47152 ( .A1(n67692), .A2(n63644), .B1(n68219), .B2(n67684), .ZN(
        n5620) );
  OAI22_X1 U47153 ( .A1(n67692), .A2(n63643), .B1(n68222), .B2(n67684), .ZN(
        n5621) );
  OAI22_X1 U47154 ( .A1(n67692), .A2(n63642), .B1(n68225), .B2(n67684), .ZN(
        n5622) );
  OAI22_X1 U47155 ( .A1(n67692), .A2(n63641), .B1(n68228), .B2(n67684), .ZN(
        n5623) );
  OAI22_X1 U47156 ( .A1(n67692), .A2(n63640), .B1(n68231), .B2(n67684), .ZN(
        n5624) );
  OAI22_X1 U47157 ( .A1(n67692), .A2(n63639), .B1(n68234), .B2(n67684), .ZN(
        n5625) );
  OAI22_X1 U47158 ( .A1(n67692), .A2(n63638), .B1(n68237), .B2(n67684), .ZN(
        n5626) );
  OAI22_X1 U47159 ( .A1(n67714), .A2(n63565), .B1(n68060), .B2(n67706), .ZN(
        n5695) );
  OAI22_X1 U47160 ( .A1(n67714), .A2(n63564), .B1(n68063), .B2(n67706), .ZN(
        n5696) );
  OAI22_X1 U47161 ( .A1(n67714), .A2(n63563), .B1(n68066), .B2(n67706), .ZN(
        n5697) );
  OAI22_X1 U47162 ( .A1(n67714), .A2(n63562), .B1(n68069), .B2(n67706), .ZN(
        n5698) );
  OAI22_X1 U47163 ( .A1(n67714), .A2(n63561), .B1(n68072), .B2(n67706), .ZN(
        n5699) );
  OAI22_X1 U47164 ( .A1(n67714), .A2(n63560), .B1(n68075), .B2(n67706), .ZN(
        n5700) );
  OAI22_X1 U47165 ( .A1(n67714), .A2(n63559), .B1(n68078), .B2(n67706), .ZN(
        n5701) );
  OAI22_X1 U47166 ( .A1(n67714), .A2(n63558), .B1(n68081), .B2(n67706), .ZN(
        n5702) );
  OAI22_X1 U47167 ( .A1(n67714), .A2(n63557), .B1(n68084), .B2(n67706), .ZN(
        n5703) );
  OAI22_X1 U47168 ( .A1(n67714), .A2(n63556), .B1(n68087), .B2(n67706), .ZN(
        n5704) );
  OAI22_X1 U47169 ( .A1(n67714), .A2(n63555), .B1(n68090), .B2(n67706), .ZN(
        n5705) );
  OAI22_X1 U47170 ( .A1(n67714), .A2(n63554), .B1(n68093), .B2(n67706), .ZN(
        n5706) );
  OAI22_X1 U47171 ( .A1(n67715), .A2(n63553), .B1(n68096), .B2(n67707), .ZN(
        n5707) );
  OAI22_X1 U47172 ( .A1(n67715), .A2(n63552), .B1(n68099), .B2(n67707), .ZN(
        n5708) );
  OAI22_X1 U47173 ( .A1(n67715), .A2(n63551), .B1(n68102), .B2(n67707), .ZN(
        n5709) );
  OAI22_X1 U47174 ( .A1(n67715), .A2(n63550), .B1(n68105), .B2(n67707), .ZN(
        n5710) );
  OAI22_X1 U47175 ( .A1(n67715), .A2(n63549), .B1(n68108), .B2(n67707), .ZN(
        n5711) );
  OAI22_X1 U47176 ( .A1(n67715), .A2(n63548), .B1(n68111), .B2(n67707), .ZN(
        n5712) );
  OAI22_X1 U47177 ( .A1(n67715), .A2(n63547), .B1(n68114), .B2(n67707), .ZN(
        n5713) );
  OAI22_X1 U47178 ( .A1(n67715), .A2(n63546), .B1(n68117), .B2(n67707), .ZN(
        n5714) );
  OAI22_X1 U47179 ( .A1(n67715), .A2(n63545), .B1(n68120), .B2(n67707), .ZN(
        n5715) );
  OAI22_X1 U47180 ( .A1(n67715), .A2(n63544), .B1(n68123), .B2(n67707), .ZN(
        n5716) );
  OAI22_X1 U47181 ( .A1(n67715), .A2(n63543), .B1(n68126), .B2(n67707), .ZN(
        n5717) );
  OAI22_X1 U47182 ( .A1(n67715), .A2(n63542), .B1(n68129), .B2(n67707), .ZN(
        n5718) );
  OAI22_X1 U47183 ( .A1(n67715), .A2(n63541), .B1(n68132), .B2(n67708), .ZN(
        n5719) );
  OAI22_X1 U47184 ( .A1(n67716), .A2(n63540), .B1(n68135), .B2(n67708), .ZN(
        n5720) );
  OAI22_X1 U47185 ( .A1(n67716), .A2(n63539), .B1(n68138), .B2(n67708), .ZN(
        n5721) );
  OAI22_X1 U47186 ( .A1(n67716), .A2(n63538), .B1(n68141), .B2(n67708), .ZN(
        n5722) );
  OAI22_X1 U47187 ( .A1(n67716), .A2(n63537), .B1(n68144), .B2(n67708), .ZN(
        n5723) );
  OAI22_X1 U47188 ( .A1(n67716), .A2(n63536), .B1(n68147), .B2(n67708), .ZN(
        n5724) );
  OAI22_X1 U47189 ( .A1(n67716), .A2(n63535), .B1(n68150), .B2(n67708), .ZN(
        n5725) );
  OAI22_X1 U47190 ( .A1(n67716), .A2(n63534), .B1(n68153), .B2(n67708), .ZN(
        n5726) );
  OAI22_X1 U47191 ( .A1(n67716), .A2(n63533), .B1(n68156), .B2(n67708), .ZN(
        n5727) );
  OAI22_X1 U47192 ( .A1(n67716), .A2(n63532), .B1(n68159), .B2(n67708), .ZN(
        n5728) );
  OAI22_X1 U47193 ( .A1(n67716), .A2(n63531), .B1(n68162), .B2(n67708), .ZN(
        n5729) );
  OAI22_X1 U47194 ( .A1(n67716), .A2(n63530), .B1(n68165), .B2(n67708), .ZN(
        n5730) );
  OAI22_X1 U47195 ( .A1(n67716), .A2(n63529), .B1(n68168), .B2(n67709), .ZN(
        n5731) );
  OAI22_X1 U47196 ( .A1(n67716), .A2(n63528), .B1(n68171), .B2(n67709), .ZN(
        n5732) );
  OAI22_X1 U47197 ( .A1(n67717), .A2(n63527), .B1(n68174), .B2(n67709), .ZN(
        n5733) );
  OAI22_X1 U47198 ( .A1(n67717), .A2(n63526), .B1(n68177), .B2(n67709), .ZN(
        n5734) );
  OAI22_X1 U47199 ( .A1(n67717), .A2(n63525), .B1(n68180), .B2(n67709), .ZN(
        n5735) );
  OAI22_X1 U47200 ( .A1(n67717), .A2(n63524), .B1(n68183), .B2(n67709), .ZN(
        n5736) );
  OAI22_X1 U47201 ( .A1(n67717), .A2(n63523), .B1(n68186), .B2(n67709), .ZN(
        n5737) );
  OAI22_X1 U47202 ( .A1(n67717), .A2(n63522), .B1(n68189), .B2(n67709), .ZN(
        n5738) );
  OAI22_X1 U47203 ( .A1(n67717), .A2(n63521), .B1(n68192), .B2(n67709), .ZN(
        n5739) );
  OAI22_X1 U47204 ( .A1(n67717), .A2(n63520), .B1(n68195), .B2(n67709), .ZN(
        n5740) );
  OAI22_X1 U47205 ( .A1(n67717), .A2(n63519), .B1(n68198), .B2(n67709), .ZN(
        n5741) );
  OAI22_X1 U47206 ( .A1(n67717), .A2(n63518), .B1(n68201), .B2(n67709), .ZN(
        n5742) );
  OAI22_X1 U47207 ( .A1(n67717), .A2(n63517), .B1(n68204), .B2(n67710), .ZN(
        n5743) );
  OAI22_X1 U47208 ( .A1(n67717), .A2(n63516), .B1(n68207), .B2(n67710), .ZN(
        n5744) );
  OAI22_X1 U47209 ( .A1(n67717), .A2(n63515), .B1(n68210), .B2(n67710), .ZN(
        n5745) );
  OAI22_X1 U47210 ( .A1(n67718), .A2(n63514), .B1(n68213), .B2(n67710), .ZN(
        n5746) );
  OAI22_X1 U47211 ( .A1(n67718), .A2(n63513), .B1(n68216), .B2(n67710), .ZN(
        n5747) );
  OAI22_X1 U47212 ( .A1(n67718), .A2(n63512), .B1(n68219), .B2(n67710), .ZN(
        n5748) );
  OAI22_X1 U47213 ( .A1(n67718), .A2(n63511), .B1(n68222), .B2(n67710), .ZN(
        n5749) );
  OAI22_X1 U47214 ( .A1(n67718), .A2(n63510), .B1(n68225), .B2(n67710), .ZN(
        n5750) );
  OAI22_X1 U47215 ( .A1(n67718), .A2(n63509), .B1(n68228), .B2(n67710), .ZN(
        n5751) );
  OAI22_X1 U47216 ( .A1(n67718), .A2(n63508), .B1(n68231), .B2(n67710), .ZN(
        n5752) );
  OAI22_X1 U47217 ( .A1(n67718), .A2(n63507), .B1(n68234), .B2(n67710), .ZN(
        n5753) );
  OAI22_X1 U47218 ( .A1(n67718), .A2(n63506), .B1(n68237), .B2(n67710), .ZN(
        n5754) );
  OAI22_X1 U47219 ( .A1(n67701), .A2(n63631), .B1(n68060), .B2(n67693), .ZN(
        n5631) );
  OAI22_X1 U47220 ( .A1(n67701), .A2(n63630), .B1(n68063), .B2(n67693), .ZN(
        n5632) );
  OAI22_X1 U47221 ( .A1(n67701), .A2(n63629), .B1(n68066), .B2(n67693), .ZN(
        n5633) );
  OAI22_X1 U47222 ( .A1(n67701), .A2(n63628), .B1(n68069), .B2(n67693), .ZN(
        n5634) );
  OAI22_X1 U47223 ( .A1(n67701), .A2(n63627), .B1(n68072), .B2(n67693), .ZN(
        n5635) );
  OAI22_X1 U47224 ( .A1(n67701), .A2(n63626), .B1(n68075), .B2(n67693), .ZN(
        n5636) );
  OAI22_X1 U47225 ( .A1(n67701), .A2(n63625), .B1(n68078), .B2(n67693), .ZN(
        n5637) );
  OAI22_X1 U47226 ( .A1(n67701), .A2(n63624), .B1(n68081), .B2(n67693), .ZN(
        n5638) );
  OAI22_X1 U47227 ( .A1(n67701), .A2(n63623), .B1(n68084), .B2(n67693), .ZN(
        n5639) );
  OAI22_X1 U47228 ( .A1(n67701), .A2(n63622), .B1(n68087), .B2(n67693), .ZN(
        n5640) );
  OAI22_X1 U47229 ( .A1(n67701), .A2(n63621), .B1(n68090), .B2(n67693), .ZN(
        n5641) );
  OAI22_X1 U47230 ( .A1(n67701), .A2(n63620), .B1(n68093), .B2(n67693), .ZN(
        n5642) );
  OAI22_X1 U47231 ( .A1(n67702), .A2(n63619), .B1(n68096), .B2(n67694), .ZN(
        n5643) );
  OAI22_X1 U47232 ( .A1(n67702), .A2(n63618), .B1(n68099), .B2(n67694), .ZN(
        n5644) );
  OAI22_X1 U47233 ( .A1(n67702), .A2(n63617), .B1(n68102), .B2(n67694), .ZN(
        n5645) );
  OAI22_X1 U47234 ( .A1(n67702), .A2(n63616), .B1(n68105), .B2(n67694), .ZN(
        n5646) );
  OAI22_X1 U47235 ( .A1(n67702), .A2(n63615), .B1(n68108), .B2(n67694), .ZN(
        n5647) );
  OAI22_X1 U47236 ( .A1(n67702), .A2(n63614), .B1(n68111), .B2(n67694), .ZN(
        n5648) );
  OAI22_X1 U47237 ( .A1(n67702), .A2(n63613), .B1(n68114), .B2(n67694), .ZN(
        n5649) );
  OAI22_X1 U47238 ( .A1(n67702), .A2(n63612), .B1(n68117), .B2(n67694), .ZN(
        n5650) );
  OAI22_X1 U47239 ( .A1(n67702), .A2(n63611), .B1(n68120), .B2(n67694), .ZN(
        n5651) );
  OAI22_X1 U47240 ( .A1(n67702), .A2(n63610), .B1(n68123), .B2(n67694), .ZN(
        n5652) );
  OAI22_X1 U47241 ( .A1(n67702), .A2(n63609), .B1(n68126), .B2(n67694), .ZN(
        n5653) );
  OAI22_X1 U47242 ( .A1(n67702), .A2(n63608), .B1(n68129), .B2(n67694), .ZN(
        n5654) );
  OAI22_X1 U47243 ( .A1(n67702), .A2(n63607), .B1(n68132), .B2(n67695), .ZN(
        n5655) );
  OAI22_X1 U47244 ( .A1(n67703), .A2(n63606), .B1(n68135), .B2(n67695), .ZN(
        n5656) );
  OAI22_X1 U47245 ( .A1(n67703), .A2(n63605), .B1(n68138), .B2(n67695), .ZN(
        n5657) );
  OAI22_X1 U47246 ( .A1(n67703), .A2(n63604), .B1(n68141), .B2(n67695), .ZN(
        n5658) );
  OAI22_X1 U47247 ( .A1(n67703), .A2(n63603), .B1(n68144), .B2(n67695), .ZN(
        n5659) );
  OAI22_X1 U47248 ( .A1(n67703), .A2(n63602), .B1(n68147), .B2(n67695), .ZN(
        n5660) );
  OAI22_X1 U47249 ( .A1(n67703), .A2(n63601), .B1(n68150), .B2(n67695), .ZN(
        n5661) );
  OAI22_X1 U47250 ( .A1(n67703), .A2(n63600), .B1(n68153), .B2(n67695), .ZN(
        n5662) );
  OAI22_X1 U47251 ( .A1(n67703), .A2(n63599), .B1(n68156), .B2(n67695), .ZN(
        n5663) );
  OAI22_X1 U47252 ( .A1(n67703), .A2(n63598), .B1(n68159), .B2(n67695), .ZN(
        n5664) );
  OAI22_X1 U47253 ( .A1(n67703), .A2(n63597), .B1(n68162), .B2(n67695), .ZN(
        n5665) );
  OAI22_X1 U47254 ( .A1(n67703), .A2(n63596), .B1(n68165), .B2(n67695), .ZN(
        n5666) );
  OAI22_X1 U47255 ( .A1(n67703), .A2(n63595), .B1(n68168), .B2(n67696), .ZN(
        n5667) );
  OAI22_X1 U47256 ( .A1(n67703), .A2(n63594), .B1(n68171), .B2(n67696), .ZN(
        n5668) );
  OAI22_X1 U47257 ( .A1(n67704), .A2(n63593), .B1(n68174), .B2(n67696), .ZN(
        n5669) );
  OAI22_X1 U47258 ( .A1(n67704), .A2(n63592), .B1(n68177), .B2(n67696), .ZN(
        n5670) );
  OAI22_X1 U47259 ( .A1(n67704), .A2(n63591), .B1(n68180), .B2(n67696), .ZN(
        n5671) );
  OAI22_X1 U47260 ( .A1(n67704), .A2(n63590), .B1(n68183), .B2(n67696), .ZN(
        n5672) );
  OAI22_X1 U47261 ( .A1(n67704), .A2(n63589), .B1(n68186), .B2(n67696), .ZN(
        n5673) );
  OAI22_X1 U47262 ( .A1(n67704), .A2(n63588), .B1(n68189), .B2(n67696), .ZN(
        n5674) );
  OAI22_X1 U47263 ( .A1(n67704), .A2(n63587), .B1(n68192), .B2(n67696), .ZN(
        n5675) );
  OAI22_X1 U47264 ( .A1(n67704), .A2(n63586), .B1(n68195), .B2(n67696), .ZN(
        n5676) );
  OAI22_X1 U47265 ( .A1(n67704), .A2(n63585), .B1(n68198), .B2(n67696), .ZN(
        n5677) );
  OAI22_X1 U47266 ( .A1(n67704), .A2(n63584), .B1(n68201), .B2(n67696), .ZN(
        n5678) );
  OAI22_X1 U47267 ( .A1(n67704), .A2(n63583), .B1(n68204), .B2(n67697), .ZN(
        n5679) );
  OAI22_X1 U47268 ( .A1(n67704), .A2(n63582), .B1(n68207), .B2(n67697), .ZN(
        n5680) );
  OAI22_X1 U47269 ( .A1(n67704), .A2(n63581), .B1(n68210), .B2(n67697), .ZN(
        n5681) );
  OAI22_X1 U47270 ( .A1(n67705), .A2(n63580), .B1(n68213), .B2(n67697), .ZN(
        n5682) );
  OAI22_X1 U47271 ( .A1(n67705), .A2(n63579), .B1(n68216), .B2(n67697), .ZN(
        n5683) );
  OAI22_X1 U47272 ( .A1(n67705), .A2(n63578), .B1(n68219), .B2(n67697), .ZN(
        n5684) );
  OAI22_X1 U47273 ( .A1(n67705), .A2(n63577), .B1(n68222), .B2(n67697), .ZN(
        n5685) );
  OAI22_X1 U47274 ( .A1(n67705), .A2(n63576), .B1(n68225), .B2(n67697), .ZN(
        n5686) );
  OAI22_X1 U47275 ( .A1(n67705), .A2(n63575), .B1(n68228), .B2(n67697), .ZN(
        n5687) );
  OAI22_X1 U47276 ( .A1(n67705), .A2(n63574), .B1(n68231), .B2(n67697), .ZN(
        n5688) );
  OAI22_X1 U47277 ( .A1(n67705), .A2(n63573), .B1(n68234), .B2(n67697), .ZN(
        n5689) );
  OAI22_X1 U47278 ( .A1(n67705), .A2(n63572), .B1(n68237), .B2(n67697), .ZN(
        n5690) );
  NAND2_X1 U47279 ( .A1(n66280), .A2(n66281), .ZN(n65108) );
  NAND2_X1 U47280 ( .A1(n66287), .A2(n66277), .ZN(n65118) );
  AND2_X1 U47281 ( .A1(n65085), .A2(n65074), .ZN(n63790) );
  OAI22_X1 U47282 ( .A1(n67943), .A2(n62691), .B1(n68058), .B2(n67935), .ZN(
        n6847) );
  OAI22_X1 U47283 ( .A1(n67943), .A2(n62690), .B1(n68061), .B2(n67935), .ZN(
        n6848) );
  OAI22_X1 U47284 ( .A1(n67943), .A2(n62689), .B1(n68064), .B2(n67935), .ZN(
        n6849) );
  OAI22_X1 U47285 ( .A1(n67943), .A2(n62688), .B1(n68067), .B2(n67935), .ZN(
        n6850) );
  OAI22_X1 U47286 ( .A1(n67943), .A2(n62687), .B1(n68070), .B2(n67935), .ZN(
        n6851) );
  OAI22_X1 U47287 ( .A1(n67943), .A2(n62686), .B1(n68073), .B2(n67935), .ZN(
        n6852) );
  OAI22_X1 U47288 ( .A1(n67943), .A2(n62685), .B1(n68076), .B2(n67935), .ZN(
        n6853) );
  OAI22_X1 U47289 ( .A1(n67943), .A2(n62684), .B1(n68079), .B2(n67935), .ZN(
        n6854) );
  OAI22_X1 U47290 ( .A1(n67943), .A2(n62683), .B1(n68082), .B2(n67935), .ZN(
        n6855) );
  OAI22_X1 U47291 ( .A1(n67943), .A2(n62682), .B1(n68085), .B2(n67935), .ZN(
        n6856) );
  OAI22_X1 U47292 ( .A1(n67943), .A2(n62681), .B1(n68088), .B2(n67935), .ZN(
        n6857) );
  OAI22_X1 U47293 ( .A1(n67943), .A2(n62680), .B1(n68091), .B2(n67935), .ZN(
        n6858) );
  OAI22_X1 U47294 ( .A1(n67944), .A2(n62679), .B1(n68094), .B2(n67936), .ZN(
        n6859) );
  OAI22_X1 U47295 ( .A1(n67944), .A2(n62678), .B1(n68097), .B2(n67936), .ZN(
        n6860) );
  OAI22_X1 U47296 ( .A1(n67944), .A2(n62677), .B1(n68100), .B2(n67936), .ZN(
        n6861) );
  OAI22_X1 U47297 ( .A1(n67944), .A2(n62676), .B1(n68103), .B2(n67936), .ZN(
        n6862) );
  OAI22_X1 U47298 ( .A1(n67944), .A2(n62675), .B1(n68106), .B2(n67936), .ZN(
        n6863) );
  OAI22_X1 U47299 ( .A1(n67944), .A2(n62674), .B1(n68109), .B2(n67936), .ZN(
        n6864) );
  OAI22_X1 U47300 ( .A1(n67944), .A2(n62673), .B1(n68112), .B2(n67936), .ZN(
        n6865) );
  OAI22_X1 U47301 ( .A1(n67944), .A2(n62672), .B1(n68115), .B2(n67936), .ZN(
        n6866) );
  OAI22_X1 U47302 ( .A1(n67944), .A2(n62671), .B1(n68118), .B2(n67936), .ZN(
        n6867) );
  OAI22_X1 U47303 ( .A1(n67944), .A2(n62670), .B1(n68121), .B2(n67936), .ZN(
        n6868) );
  OAI22_X1 U47304 ( .A1(n67944), .A2(n62669), .B1(n68124), .B2(n67936), .ZN(
        n6869) );
  OAI22_X1 U47305 ( .A1(n67944), .A2(n62668), .B1(n68127), .B2(n67936), .ZN(
        n6870) );
  OAI22_X1 U47306 ( .A1(n67944), .A2(n62667), .B1(n68130), .B2(n67937), .ZN(
        n6871) );
  OAI22_X1 U47307 ( .A1(n67945), .A2(n62666), .B1(n68133), .B2(n67937), .ZN(
        n6872) );
  OAI22_X1 U47308 ( .A1(n67945), .A2(n62665), .B1(n68136), .B2(n67937), .ZN(
        n6873) );
  OAI22_X1 U47309 ( .A1(n67945), .A2(n62664), .B1(n68139), .B2(n67937), .ZN(
        n6874) );
  OAI22_X1 U47310 ( .A1(n67945), .A2(n62663), .B1(n68142), .B2(n67937), .ZN(
        n6875) );
  OAI22_X1 U47311 ( .A1(n67945), .A2(n62662), .B1(n68145), .B2(n67937), .ZN(
        n6876) );
  OAI22_X1 U47312 ( .A1(n67945), .A2(n62661), .B1(n68148), .B2(n67937), .ZN(
        n6877) );
  OAI22_X1 U47313 ( .A1(n67945), .A2(n62660), .B1(n68151), .B2(n67937), .ZN(
        n6878) );
  OAI22_X1 U47314 ( .A1(n67945), .A2(n62659), .B1(n68154), .B2(n67937), .ZN(
        n6879) );
  OAI22_X1 U47315 ( .A1(n67945), .A2(n62658), .B1(n68157), .B2(n67937), .ZN(
        n6880) );
  OAI22_X1 U47316 ( .A1(n67945), .A2(n62657), .B1(n68160), .B2(n67937), .ZN(
        n6881) );
  OAI22_X1 U47317 ( .A1(n67945), .A2(n62656), .B1(n68163), .B2(n67937), .ZN(
        n6882) );
  OAI22_X1 U47318 ( .A1(n67945), .A2(n62655), .B1(n68166), .B2(n67938), .ZN(
        n6883) );
  OAI22_X1 U47319 ( .A1(n67945), .A2(n62654), .B1(n68169), .B2(n67938), .ZN(
        n6884) );
  OAI22_X1 U47320 ( .A1(n67946), .A2(n62653), .B1(n68172), .B2(n67938), .ZN(
        n6885) );
  OAI22_X1 U47321 ( .A1(n67946), .A2(n62652), .B1(n68175), .B2(n67938), .ZN(
        n6886) );
  OAI22_X1 U47322 ( .A1(n67946), .A2(n62651), .B1(n68178), .B2(n67938), .ZN(
        n6887) );
  OAI22_X1 U47323 ( .A1(n67946), .A2(n62650), .B1(n68181), .B2(n67938), .ZN(
        n6888) );
  OAI22_X1 U47324 ( .A1(n67946), .A2(n62649), .B1(n68184), .B2(n67938), .ZN(
        n6889) );
  OAI22_X1 U47325 ( .A1(n67946), .A2(n62648), .B1(n68187), .B2(n67938), .ZN(
        n6890) );
  OAI22_X1 U47326 ( .A1(n67946), .A2(n62647), .B1(n68190), .B2(n67938), .ZN(
        n6891) );
  OAI22_X1 U47327 ( .A1(n67946), .A2(n62646), .B1(n68193), .B2(n67938), .ZN(
        n6892) );
  OAI22_X1 U47328 ( .A1(n67946), .A2(n62645), .B1(n68196), .B2(n67938), .ZN(
        n6893) );
  OAI22_X1 U47329 ( .A1(n67946), .A2(n62644), .B1(n68199), .B2(n67938), .ZN(
        n6894) );
  OAI22_X1 U47330 ( .A1(n67946), .A2(n62643), .B1(n68202), .B2(n67939), .ZN(
        n6895) );
  OAI22_X1 U47331 ( .A1(n67946), .A2(n62642), .B1(n68205), .B2(n67939), .ZN(
        n6896) );
  OAI22_X1 U47332 ( .A1(n67946), .A2(n62641), .B1(n68208), .B2(n67939), .ZN(
        n6897) );
  OAI22_X1 U47333 ( .A1(n67947), .A2(n62640), .B1(n68211), .B2(n67939), .ZN(
        n6898) );
  OAI22_X1 U47334 ( .A1(n67947), .A2(n62639), .B1(n68214), .B2(n67939), .ZN(
        n6899) );
  OAI22_X1 U47335 ( .A1(n67947), .A2(n62638), .B1(n68217), .B2(n67939), .ZN(
        n6900) );
  OAI22_X1 U47336 ( .A1(n67947), .A2(n62637), .B1(n68220), .B2(n67939), .ZN(
        n6901) );
  OAI22_X1 U47337 ( .A1(n67947), .A2(n62636), .B1(n68223), .B2(n67939), .ZN(
        n6902) );
  OAI22_X1 U47338 ( .A1(n67947), .A2(n62635), .B1(n68226), .B2(n67939), .ZN(
        n6903) );
  OAI22_X1 U47339 ( .A1(n67947), .A2(n62634), .B1(n68229), .B2(n67939), .ZN(
        n6904) );
  OAI22_X1 U47340 ( .A1(n67947), .A2(n62633), .B1(n68232), .B2(n67939), .ZN(
        n6905) );
  OAI22_X1 U47341 ( .A1(n67947), .A2(n62632), .B1(n68235), .B2(n67939), .ZN(
        n6906) );
  OAI22_X1 U47342 ( .A1(n67956), .A2(n62624), .B1(n68058), .B2(n67948), .ZN(
        n6911) );
  OAI22_X1 U47343 ( .A1(n67956), .A2(n62623), .B1(n68061), .B2(n67948), .ZN(
        n6912) );
  OAI22_X1 U47344 ( .A1(n67956), .A2(n62622), .B1(n68064), .B2(n67948), .ZN(
        n6913) );
  OAI22_X1 U47345 ( .A1(n67956), .A2(n62621), .B1(n68067), .B2(n67948), .ZN(
        n6914) );
  OAI22_X1 U47346 ( .A1(n67956), .A2(n62620), .B1(n68070), .B2(n67948), .ZN(
        n6915) );
  OAI22_X1 U47347 ( .A1(n67956), .A2(n62619), .B1(n68073), .B2(n67948), .ZN(
        n6916) );
  OAI22_X1 U47348 ( .A1(n67956), .A2(n62618), .B1(n68076), .B2(n67948), .ZN(
        n6917) );
  OAI22_X1 U47349 ( .A1(n67956), .A2(n62617), .B1(n68079), .B2(n67948), .ZN(
        n6918) );
  OAI22_X1 U47350 ( .A1(n67956), .A2(n62616), .B1(n68082), .B2(n67948), .ZN(
        n6919) );
  OAI22_X1 U47351 ( .A1(n67956), .A2(n62615), .B1(n68085), .B2(n67948), .ZN(
        n6920) );
  OAI22_X1 U47352 ( .A1(n67956), .A2(n62614), .B1(n68088), .B2(n67948), .ZN(
        n6921) );
  OAI22_X1 U47353 ( .A1(n67956), .A2(n62613), .B1(n68091), .B2(n67948), .ZN(
        n6922) );
  OAI22_X1 U47354 ( .A1(n67957), .A2(n62612), .B1(n68094), .B2(n67949), .ZN(
        n6923) );
  OAI22_X1 U47355 ( .A1(n67957), .A2(n62611), .B1(n68097), .B2(n67949), .ZN(
        n6924) );
  OAI22_X1 U47356 ( .A1(n67957), .A2(n62610), .B1(n68100), .B2(n67949), .ZN(
        n6925) );
  OAI22_X1 U47357 ( .A1(n67957), .A2(n62609), .B1(n68103), .B2(n67949), .ZN(
        n6926) );
  OAI22_X1 U47358 ( .A1(n67957), .A2(n62608), .B1(n68106), .B2(n67949), .ZN(
        n6927) );
  OAI22_X1 U47359 ( .A1(n67957), .A2(n62607), .B1(n68109), .B2(n67949), .ZN(
        n6928) );
  OAI22_X1 U47360 ( .A1(n67957), .A2(n62606), .B1(n68112), .B2(n67949), .ZN(
        n6929) );
  OAI22_X1 U47361 ( .A1(n67957), .A2(n62605), .B1(n68115), .B2(n67949), .ZN(
        n6930) );
  OAI22_X1 U47362 ( .A1(n67957), .A2(n62604), .B1(n68118), .B2(n67949), .ZN(
        n6931) );
  OAI22_X1 U47363 ( .A1(n67957), .A2(n62603), .B1(n68121), .B2(n67949), .ZN(
        n6932) );
  OAI22_X1 U47364 ( .A1(n67957), .A2(n62602), .B1(n68124), .B2(n67949), .ZN(
        n6933) );
  OAI22_X1 U47365 ( .A1(n67957), .A2(n62601), .B1(n68127), .B2(n67949), .ZN(
        n6934) );
  OAI22_X1 U47366 ( .A1(n67957), .A2(n62600), .B1(n68130), .B2(n67950), .ZN(
        n6935) );
  OAI22_X1 U47367 ( .A1(n67958), .A2(n62599), .B1(n68133), .B2(n67950), .ZN(
        n6936) );
  OAI22_X1 U47368 ( .A1(n67958), .A2(n62598), .B1(n68136), .B2(n67950), .ZN(
        n6937) );
  OAI22_X1 U47369 ( .A1(n67958), .A2(n62597), .B1(n68139), .B2(n67950), .ZN(
        n6938) );
  OAI22_X1 U47370 ( .A1(n67958), .A2(n62596), .B1(n68142), .B2(n67950), .ZN(
        n6939) );
  OAI22_X1 U47371 ( .A1(n67958), .A2(n62595), .B1(n68145), .B2(n67950), .ZN(
        n6940) );
  OAI22_X1 U47372 ( .A1(n67958), .A2(n62594), .B1(n68148), .B2(n67950), .ZN(
        n6941) );
  OAI22_X1 U47373 ( .A1(n67958), .A2(n62593), .B1(n68151), .B2(n67950), .ZN(
        n6942) );
  OAI22_X1 U47374 ( .A1(n67958), .A2(n62592), .B1(n68154), .B2(n67950), .ZN(
        n6943) );
  OAI22_X1 U47375 ( .A1(n67958), .A2(n62591), .B1(n68157), .B2(n67950), .ZN(
        n6944) );
  OAI22_X1 U47376 ( .A1(n67958), .A2(n62590), .B1(n68160), .B2(n67950), .ZN(
        n6945) );
  OAI22_X1 U47377 ( .A1(n67958), .A2(n62589), .B1(n68163), .B2(n67950), .ZN(
        n6946) );
  OAI22_X1 U47378 ( .A1(n67958), .A2(n62588), .B1(n68166), .B2(n67951), .ZN(
        n6947) );
  OAI22_X1 U47379 ( .A1(n67958), .A2(n62587), .B1(n68169), .B2(n67951), .ZN(
        n6948) );
  OAI22_X1 U47380 ( .A1(n67959), .A2(n62586), .B1(n68172), .B2(n67951), .ZN(
        n6949) );
  OAI22_X1 U47381 ( .A1(n67959), .A2(n62585), .B1(n68175), .B2(n67951), .ZN(
        n6950) );
  OAI22_X1 U47382 ( .A1(n67959), .A2(n62584), .B1(n68178), .B2(n67951), .ZN(
        n6951) );
  OAI22_X1 U47383 ( .A1(n67959), .A2(n62583), .B1(n68181), .B2(n67951), .ZN(
        n6952) );
  OAI22_X1 U47384 ( .A1(n67959), .A2(n62582), .B1(n68184), .B2(n67951), .ZN(
        n6953) );
  OAI22_X1 U47385 ( .A1(n67959), .A2(n62581), .B1(n68187), .B2(n67951), .ZN(
        n6954) );
  OAI22_X1 U47386 ( .A1(n67959), .A2(n62580), .B1(n68190), .B2(n67951), .ZN(
        n6955) );
  OAI22_X1 U47387 ( .A1(n67959), .A2(n62579), .B1(n68193), .B2(n67951), .ZN(
        n6956) );
  OAI22_X1 U47388 ( .A1(n67959), .A2(n62578), .B1(n68196), .B2(n67951), .ZN(
        n6957) );
  OAI22_X1 U47389 ( .A1(n67959), .A2(n62577), .B1(n68199), .B2(n67951), .ZN(
        n6958) );
  OAI22_X1 U47390 ( .A1(n67959), .A2(n62576), .B1(n68202), .B2(n67952), .ZN(
        n6959) );
  OAI22_X1 U47391 ( .A1(n67959), .A2(n62575), .B1(n68205), .B2(n67952), .ZN(
        n6960) );
  OAI22_X1 U47392 ( .A1(n67959), .A2(n62574), .B1(n68208), .B2(n67952), .ZN(
        n6961) );
  OAI22_X1 U47393 ( .A1(n67960), .A2(n62573), .B1(n68211), .B2(n67952), .ZN(
        n6962) );
  OAI22_X1 U47394 ( .A1(n67960), .A2(n62572), .B1(n68214), .B2(n67952), .ZN(
        n6963) );
  OAI22_X1 U47395 ( .A1(n67960), .A2(n62571), .B1(n68217), .B2(n67952), .ZN(
        n6964) );
  OAI22_X1 U47396 ( .A1(n67960), .A2(n62570), .B1(n68220), .B2(n67952), .ZN(
        n6965) );
  OAI22_X1 U47397 ( .A1(n67960), .A2(n62569), .B1(n68223), .B2(n67952), .ZN(
        n6966) );
  OAI22_X1 U47398 ( .A1(n67960), .A2(n62568), .B1(n68226), .B2(n67952), .ZN(
        n6967) );
  OAI22_X1 U47399 ( .A1(n67960), .A2(n62567), .B1(n68229), .B2(n67952), .ZN(
        n6968) );
  OAI22_X1 U47400 ( .A1(n67960), .A2(n62566), .B1(n68232), .B2(n67952), .ZN(
        n6969) );
  OAI22_X1 U47401 ( .A1(n67960), .A2(n62565), .B1(n68235), .B2(n67952), .ZN(
        n6970) );
  OAI22_X1 U47402 ( .A1(n68047), .A2(n62155), .B1(n68058), .B2(n68039), .ZN(
        n7359) );
  OAI22_X1 U47403 ( .A1(n68047), .A2(n62154), .B1(n68061), .B2(n68039), .ZN(
        n7360) );
  OAI22_X1 U47404 ( .A1(n68047), .A2(n62153), .B1(n68064), .B2(n68039), .ZN(
        n7361) );
  OAI22_X1 U47405 ( .A1(n68047), .A2(n62152), .B1(n68067), .B2(n68039), .ZN(
        n7362) );
  OAI22_X1 U47406 ( .A1(n68047), .A2(n62151), .B1(n68070), .B2(n68039), .ZN(
        n7363) );
  OAI22_X1 U47407 ( .A1(n68047), .A2(n62150), .B1(n68073), .B2(n68039), .ZN(
        n7364) );
  OAI22_X1 U47408 ( .A1(n68047), .A2(n62149), .B1(n68076), .B2(n68039), .ZN(
        n7365) );
  OAI22_X1 U47409 ( .A1(n68047), .A2(n62148), .B1(n68079), .B2(n68039), .ZN(
        n7366) );
  OAI22_X1 U47410 ( .A1(n68047), .A2(n62147), .B1(n68082), .B2(n68039), .ZN(
        n7367) );
  OAI22_X1 U47411 ( .A1(n68047), .A2(n62146), .B1(n68085), .B2(n68039), .ZN(
        n7368) );
  OAI22_X1 U47412 ( .A1(n68047), .A2(n62145), .B1(n68088), .B2(n68039), .ZN(
        n7369) );
  OAI22_X1 U47413 ( .A1(n68047), .A2(n62144), .B1(n68091), .B2(n68039), .ZN(
        n7370) );
  OAI22_X1 U47414 ( .A1(n68048), .A2(n62143), .B1(n68094), .B2(n68040), .ZN(
        n7371) );
  OAI22_X1 U47415 ( .A1(n68048), .A2(n62142), .B1(n68097), .B2(n68040), .ZN(
        n7372) );
  OAI22_X1 U47416 ( .A1(n68048), .A2(n62141), .B1(n68100), .B2(n68040), .ZN(
        n7373) );
  OAI22_X1 U47417 ( .A1(n68048), .A2(n62140), .B1(n68103), .B2(n68040), .ZN(
        n7374) );
  OAI22_X1 U47418 ( .A1(n68048), .A2(n62139), .B1(n68106), .B2(n68040), .ZN(
        n7375) );
  OAI22_X1 U47419 ( .A1(n68048), .A2(n62138), .B1(n68109), .B2(n68040), .ZN(
        n7376) );
  OAI22_X1 U47420 ( .A1(n68048), .A2(n62137), .B1(n68112), .B2(n68040), .ZN(
        n7377) );
  OAI22_X1 U47421 ( .A1(n68048), .A2(n62136), .B1(n68115), .B2(n68040), .ZN(
        n7378) );
  OAI22_X1 U47422 ( .A1(n68048), .A2(n62135), .B1(n68118), .B2(n68040), .ZN(
        n7379) );
  OAI22_X1 U47423 ( .A1(n68048), .A2(n62134), .B1(n68121), .B2(n68040), .ZN(
        n7380) );
  OAI22_X1 U47424 ( .A1(n68048), .A2(n62133), .B1(n68124), .B2(n68040), .ZN(
        n7381) );
  OAI22_X1 U47425 ( .A1(n68048), .A2(n62132), .B1(n68127), .B2(n68040), .ZN(
        n7382) );
  OAI22_X1 U47426 ( .A1(n68048), .A2(n62131), .B1(n68130), .B2(n68041), .ZN(
        n7383) );
  OAI22_X1 U47427 ( .A1(n68049), .A2(n62130), .B1(n68133), .B2(n68041), .ZN(
        n7384) );
  OAI22_X1 U47428 ( .A1(n68049), .A2(n62129), .B1(n68136), .B2(n68041), .ZN(
        n7385) );
  OAI22_X1 U47429 ( .A1(n68049), .A2(n62128), .B1(n68139), .B2(n68041), .ZN(
        n7386) );
  OAI22_X1 U47430 ( .A1(n68049), .A2(n62127), .B1(n68142), .B2(n68041), .ZN(
        n7387) );
  OAI22_X1 U47431 ( .A1(n68049), .A2(n62126), .B1(n68145), .B2(n68041), .ZN(
        n7388) );
  OAI22_X1 U47432 ( .A1(n68049), .A2(n62125), .B1(n68148), .B2(n68041), .ZN(
        n7389) );
  OAI22_X1 U47433 ( .A1(n68049), .A2(n62124), .B1(n68151), .B2(n68041), .ZN(
        n7390) );
  OAI22_X1 U47434 ( .A1(n68049), .A2(n62123), .B1(n68154), .B2(n68041), .ZN(
        n7391) );
  OAI22_X1 U47435 ( .A1(n68049), .A2(n62122), .B1(n68157), .B2(n68041), .ZN(
        n7392) );
  OAI22_X1 U47436 ( .A1(n68049), .A2(n62121), .B1(n68160), .B2(n68041), .ZN(
        n7393) );
  OAI22_X1 U47437 ( .A1(n68049), .A2(n62120), .B1(n68163), .B2(n68041), .ZN(
        n7394) );
  OAI22_X1 U47438 ( .A1(n68049), .A2(n62119), .B1(n68166), .B2(n68042), .ZN(
        n7395) );
  OAI22_X1 U47439 ( .A1(n68049), .A2(n62118), .B1(n68169), .B2(n68042), .ZN(
        n7396) );
  OAI22_X1 U47440 ( .A1(n68050), .A2(n62117), .B1(n68172), .B2(n68042), .ZN(
        n7397) );
  OAI22_X1 U47441 ( .A1(n68050), .A2(n62116), .B1(n68175), .B2(n68042), .ZN(
        n7398) );
  OAI22_X1 U47442 ( .A1(n68050), .A2(n62115), .B1(n68178), .B2(n68042), .ZN(
        n7399) );
  OAI22_X1 U47443 ( .A1(n68050), .A2(n62114), .B1(n68181), .B2(n68042), .ZN(
        n7400) );
  OAI22_X1 U47444 ( .A1(n68050), .A2(n62113), .B1(n68184), .B2(n68042), .ZN(
        n7401) );
  OAI22_X1 U47445 ( .A1(n68050), .A2(n62112), .B1(n68187), .B2(n68042), .ZN(
        n7402) );
  OAI22_X1 U47446 ( .A1(n68050), .A2(n62111), .B1(n68190), .B2(n68042), .ZN(
        n7403) );
  OAI22_X1 U47447 ( .A1(n68050), .A2(n62110), .B1(n68193), .B2(n68042), .ZN(
        n7404) );
  OAI22_X1 U47448 ( .A1(n68050), .A2(n62109), .B1(n68196), .B2(n68042), .ZN(
        n7405) );
  OAI22_X1 U47449 ( .A1(n68050), .A2(n62108), .B1(n68199), .B2(n68042), .ZN(
        n7406) );
  OAI22_X1 U47450 ( .A1(n68050), .A2(n62107), .B1(n68202), .B2(n68043), .ZN(
        n7407) );
  OAI22_X1 U47451 ( .A1(n68050), .A2(n62106), .B1(n68205), .B2(n68043), .ZN(
        n7408) );
  OAI22_X1 U47452 ( .A1(n68050), .A2(n62105), .B1(n68208), .B2(n68043), .ZN(
        n7409) );
  OAI22_X1 U47453 ( .A1(n68051), .A2(n62104), .B1(n68211), .B2(n68043), .ZN(
        n7410) );
  OAI22_X1 U47454 ( .A1(n68051), .A2(n62103), .B1(n68214), .B2(n68043), .ZN(
        n7411) );
  OAI22_X1 U47455 ( .A1(n68051), .A2(n62102), .B1(n68217), .B2(n68043), .ZN(
        n7412) );
  OAI22_X1 U47456 ( .A1(n68051), .A2(n62101), .B1(n68220), .B2(n68043), .ZN(
        n7413) );
  OAI22_X1 U47457 ( .A1(n68051), .A2(n62100), .B1(n68223), .B2(n68043), .ZN(
        n7414) );
  OAI22_X1 U47458 ( .A1(n68051), .A2(n62099), .B1(n68226), .B2(n68043), .ZN(
        n7415) );
  OAI22_X1 U47459 ( .A1(n68051), .A2(n62098), .B1(n68229), .B2(n68043), .ZN(
        n7416) );
  OAI22_X1 U47460 ( .A1(n68051), .A2(n62097), .B1(n68232), .B2(n68043), .ZN(
        n7417) );
  OAI22_X1 U47461 ( .A1(n68051), .A2(n62096), .B1(n68235), .B2(n68043), .ZN(
        n7418) );
  OAI22_X1 U47462 ( .A1(n68008), .A2(n62355), .B1(n68058), .B2(n68000), .ZN(
        n7167) );
  OAI22_X1 U47463 ( .A1(n68008), .A2(n62354), .B1(n68061), .B2(n68000), .ZN(
        n7168) );
  OAI22_X1 U47464 ( .A1(n68008), .A2(n62353), .B1(n68064), .B2(n68000), .ZN(
        n7169) );
  OAI22_X1 U47465 ( .A1(n68008), .A2(n62352), .B1(n68067), .B2(n68000), .ZN(
        n7170) );
  OAI22_X1 U47466 ( .A1(n68008), .A2(n62351), .B1(n68070), .B2(n68000), .ZN(
        n7171) );
  OAI22_X1 U47467 ( .A1(n68008), .A2(n62350), .B1(n68073), .B2(n68000), .ZN(
        n7172) );
  OAI22_X1 U47468 ( .A1(n68008), .A2(n62349), .B1(n68076), .B2(n68000), .ZN(
        n7173) );
  OAI22_X1 U47469 ( .A1(n68008), .A2(n62348), .B1(n68079), .B2(n68000), .ZN(
        n7174) );
  OAI22_X1 U47470 ( .A1(n68008), .A2(n62347), .B1(n68082), .B2(n68000), .ZN(
        n7175) );
  OAI22_X1 U47471 ( .A1(n68008), .A2(n62346), .B1(n68085), .B2(n68000), .ZN(
        n7176) );
  OAI22_X1 U47472 ( .A1(n68008), .A2(n62345), .B1(n68088), .B2(n68000), .ZN(
        n7177) );
  OAI22_X1 U47473 ( .A1(n68008), .A2(n62344), .B1(n68091), .B2(n68000), .ZN(
        n7178) );
  OAI22_X1 U47474 ( .A1(n68009), .A2(n62343), .B1(n68094), .B2(n68001), .ZN(
        n7179) );
  OAI22_X1 U47475 ( .A1(n68009), .A2(n62342), .B1(n68097), .B2(n68001), .ZN(
        n7180) );
  OAI22_X1 U47476 ( .A1(n68009), .A2(n62341), .B1(n68100), .B2(n68001), .ZN(
        n7181) );
  OAI22_X1 U47477 ( .A1(n68009), .A2(n62340), .B1(n68103), .B2(n68001), .ZN(
        n7182) );
  OAI22_X1 U47478 ( .A1(n68009), .A2(n62339), .B1(n68106), .B2(n68001), .ZN(
        n7183) );
  OAI22_X1 U47479 ( .A1(n68009), .A2(n62338), .B1(n68109), .B2(n68001), .ZN(
        n7184) );
  OAI22_X1 U47480 ( .A1(n68009), .A2(n62337), .B1(n68112), .B2(n68001), .ZN(
        n7185) );
  OAI22_X1 U47481 ( .A1(n68009), .A2(n62336), .B1(n68115), .B2(n68001), .ZN(
        n7186) );
  OAI22_X1 U47482 ( .A1(n68009), .A2(n62335), .B1(n68118), .B2(n68001), .ZN(
        n7187) );
  OAI22_X1 U47483 ( .A1(n68009), .A2(n62334), .B1(n68121), .B2(n68001), .ZN(
        n7188) );
  OAI22_X1 U47484 ( .A1(n68009), .A2(n62333), .B1(n68124), .B2(n68001), .ZN(
        n7189) );
  OAI22_X1 U47485 ( .A1(n68009), .A2(n62332), .B1(n68127), .B2(n68001), .ZN(
        n7190) );
  OAI22_X1 U47486 ( .A1(n68009), .A2(n62331), .B1(n68130), .B2(n68002), .ZN(
        n7191) );
  OAI22_X1 U47487 ( .A1(n68010), .A2(n62330), .B1(n68133), .B2(n68002), .ZN(
        n7192) );
  OAI22_X1 U47488 ( .A1(n68010), .A2(n62329), .B1(n68136), .B2(n68002), .ZN(
        n7193) );
  OAI22_X1 U47489 ( .A1(n68010), .A2(n62328), .B1(n68139), .B2(n68002), .ZN(
        n7194) );
  OAI22_X1 U47490 ( .A1(n68010), .A2(n62327), .B1(n68142), .B2(n68002), .ZN(
        n7195) );
  OAI22_X1 U47491 ( .A1(n68010), .A2(n62326), .B1(n68145), .B2(n68002), .ZN(
        n7196) );
  OAI22_X1 U47492 ( .A1(n68010), .A2(n62325), .B1(n68148), .B2(n68002), .ZN(
        n7197) );
  OAI22_X1 U47493 ( .A1(n68010), .A2(n62324), .B1(n68151), .B2(n68002), .ZN(
        n7198) );
  OAI22_X1 U47494 ( .A1(n68010), .A2(n62323), .B1(n68154), .B2(n68002), .ZN(
        n7199) );
  OAI22_X1 U47495 ( .A1(n68010), .A2(n62322), .B1(n68157), .B2(n68002), .ZN(
        n7200) );
  OAI22_X1 U47496 ( .A1(n68010), .A2(n62321), .B1(n68160), .B2(n68002), .ZN(
        n7201) );
  OAI22_X1 U47497 ( .A1(n68010), .A2(n62320), .B1(n68163), .B2(n68002), .ZN(
        n7202) );
  OAI22_X1 U47498 ( .A1(n68010), .A2(n62319), .B1(n68166), .B2(n68003), .ZN(
        n7203) );
  OAI22_X1 U47499 ( .A1(n68010), .A2(n62318), .B1(n68169), .B2(n68003), .ZN(
        n7204) );
  OAI22_X1 U47500 ( .A1(n68011), .A2(n62317), .B1(n68172), .B2(n68003), .ZN(
        n7205) );
  OAI22_X1 U47501 ( .A1(n68011), .A2(n62316), .B1(n68175), .B2(n68003), .ZN(
        n7206) );
  OAI22_X1 U47502 ( .A1(n68011), .A2(n62315), .B1(n68178), .B2(n68003), .ZN(
        n7207) );
  OAI22_X1 U47503 ( .A1(n68011), .A2(n62314), .B1(n68181), .B2(n68003), .ZN(
        n7208) );
  OAI22_X1 U47504 ( .A1(n68011), .A2(n62313), .B1(n68184), .B2(n68003), .ZN(
        n7209) );
  OAI22_X1 U47505 ( .A1(n68011), .A2(n62312), .B1(n68187), .B2(n68003), .ZN(
        n7210) );
  OAI22_X1 U47506 ( .A1(n68011), .A2(n62311), .B1(n68190), .B2(n68003), .ZN(
        n7211) );
  OAI22_X1 U47507 ( .A1(n68011), .A2(n62310), .B1(n68193), .B2(n68003), .ZN(
        n7212) );
  OAI22_X1 U47508 ( .A1(n68011), .A2(n62309), .B1(n68196), .B2(n68003), .ZN(
        n7213) );
  OAI22_X1 U47509 ( .A1(n68011), .A2(n62308), .B1(n68199), .B2(n68003), .ZN(
        n7214) );
  OAI22_X1 U47510 ( .A1(n68011), .A2(n62307), .B1(n68202), .B2(n68004), .ZN(
        n7215) );
  OAI22_X1 U47511 ( .A1(n68011), .A2(n62306), .B1(n68205), .B2(n68004), .ZN(
        n7216) );
  OAI22_X1 U47512 ( .A1(n68011), .A2(n62305), .B1(n68208), .B2(n68004), .ZN(
        n7217) );
  OAI22_X1 U47513 ( .A1(n68012), .A2(n62304), .B1(n68211), .B2(n68004), .ZN(
        n7218) );
  OAI22_X1 U47514 ( .A1(n68012), .A2(n62303), .B1(n68214), .B2(n68004), .ZN(
        n7219) );
  OAI22_X1 U47515 ( .A1(n68012), .A2(n62302), .B1(n68217), .B2(n68004), .ZN(
        n7220) );
  OAI22_X1 U47516 ( .A1(n68012), .A2(n62301), .B1(n68220), .B2(n68004), .ZN(
        n7221) );
  OAI22_X1 U47517 ( .A1(n68012), .A2(n62300), .B1(n68223), .B2(n68004), .ZN(
        n7222) );
  OAI22_X1 U47518 ( .A1(n68012), .A2(n62299), .B1(n68226), .B2(n68004), .ZN(
        n7223) );
  OAI22_X1 U47519 ( .A1(n68012), .A2(n62298), .B1(n68229), .B2(n68004), .ZN(
        n7224) );
  OAI22_X1 U47520 ( .A1(n68012), .A2(n62297), .B1(n68232), .B2(n68004), .ZN(
        n7225) );
  OAI22_X1 U47521 ( .A1(n68012), .A2(n62296), .B1(n68235), .B2(n68004), .ZN(
        n7226) );
  OAI22_X1 U47522 ( .A1(n67969), .A2(n62558), .B1(n68058), .B2(n67961), .ZN(
        n6975) );
  OAI22_X1 U47523 ( .A1(n67969), .A2(n62557), .B1(n68061), .B2(n67961), .ZN(
        n6976) );
  OAI22_X1 U47524 ( .A1(n67969), .A2(n62556), .B1(n68064), .B2(n67961), .ZN(
        n6977) );
  OAI22_X1 U47525 ( .A1(n67969), .A2(n62555), .B1(n68067), .B2(n67961), .ZN(
        n6978) );
  OAI22_X1 U47526 ( .A1(n67969), .A2(n62554), .B1(n68070), .B2(n67961), .ZN(
        n6979) );
  OAI22_X1 U47527 ( .A1(n67969), .A2(n62553), .B1(n68073), .B2(n67961), .ZN(
        n6980) );
  OAI22_X1 U47528 ( .A1(n67969), .A2(n62552), .B1(n68076), .B2(n67961), .ZN(
        n6981) );
  OAI22_X1 U47529 ( .A1(n67969), .A2(n62551), .B1(n68079), .B2(n67961), .ZN(
        n6982) );
  OAI22_X1 U47530 ( .A1(n67969), .A2(n62550), .B1(n68082), .B2(n67961), .ZN(
        n6983) );
  OAI22_X1 U47531 ( .A1(n67969), .A2(n62549), .B1(n68085), .B2(n67961), .ZN(
        n6984) );
  OAI22_X1 U47532 ( .A1(n67969), .A2(n62548), .B1(n68088), .B2(n67961), .ZN(
        n6985) );
  OAI22_X1 U47533 ( .A1(n67969), .A2(n62547), .B1(n68091), .B2(n67961), .ZN(
        n6986) );
  OAI22_X1 U47534 ( .A1(n67970), .A2(n62546), .B1(n68094), .B2(n67962), .ZN(
        n6987) );
  OAI22_X1 U47535 ( .A1(n67970), .A2(n62545), .B1(n68097), .B2(n67962), .ZN(
        n6988) );
  OAI22_X1 U47536 ( .A1(n67970), .A2(n62544), .B1(n68100), .B2(n67962), .ZN(
        n6989) );
  OAI22_X1 U47537 ( .A1(n67970), .A2(n62543), .B1(n68103), .B2(n67962), .ZN(
        n6990) );
  OAI22_X1 U47538 ( .A1(n67970), .A2(n62542), .B1(n68106), .B2(n67962), .ZN(
        n6991) );
  OAI22_X1 U47539 ( .A1(n67970), .A2(n62541), .B1(n68109), .B2(n67962), .ZN(
        n6992) );
  OAI22_X1 U47540 ( .A1(n67970), .A2(n62540), .B1(n68112), .B2(n67962), .ZN(
        n6993) );
  OAI22_X1 U47541 ( .A1(n67970), .A2(n62539), .B1(n68115), .B2(n67962), .ZN(
        n6994) );
  OAI22_X1 U47542 ( .A1(n67970), .A2(n62538), .B1(n68118), .B2(n67962), .ZN(
        n6995) );
  OAI22_X1 U47543 ( .A1(n67970), .A2(n62537), .B1(n68121), .B2(n67962), .ZN(
        n6996) );
  OAI22_X1 U47544 ( .A1(n67970), .A2(n62536), .B1(n68124), .B2(n67962), .ZN(
        n6997) );
  OAI22_X1 U47545 ( .A1(n67970), .A2(n62535), .B1(n68127), .B2(n67962), .ZN(
        n6998) );
  OAI22_X1 U47546 ( .A1(n67970), .A2(n62534), .B1(n68130), .B2(n67963), .ZN(
        n6999) );
  OAI22_X1 U47547 ( .A1(n67971), .A2(n62533), .B1(n68133), .B2(n67963), .ZN(
        n7000) );
  OAI22_X1 U47548 ( .A1(n67971), .A2(n62532), .B1(n68136), .B2(n67963), .ZN(
        n7001) );
  OAI22_X1 U47549 ( .A1(n67971), .A2(n62531), .B1(n68139), .B2(n67963), .ZN(
        n7002) );
  OAI22_X1 U47550 ( .A1(n67971), .A2(n62530), .B1(n68142), .B2(n67963), .ZN(
        n7003) );
  OAI22_X1 U47551 ( .A1(n67971), .A2(n62529), .B1(n68145), .B2(n67963), .ZN(
        n7004) );
  OAI22_X1 U47552 ( .A1(n67971), .A2(n62528), .B1(n68148), .B2(n67963), .ZN(
        n7005) );
  OAI22_X1 U47553 ( .A1(n67971), .A2(n62527), .B1(n68151), .B2(n67963), .ZN(
        n7006) );
  OAI22_X1 U47554 ( .A1(n67971), .A2(n62526), .B1(n68154), .B2(n67963), .ZN(
        n7007) );
  OAI22_X1 U47555 ( .A1(n67971), .A2(n62525), .B1(n68157), .B2(n67963), .ZN(
        n7008) );
  OAI22_X1 U47556 ( .A1(n67971), .A2(n62524), .B1(n68160), .B2(n67963), .ZN(
        n7009) );
  OAI22_X1 U47557 ( .A1(n67971), .A2(n62523), .B1(n68163), .B2(n67963), .ZN(
        n7010) );
  OAI22_X1 U47558 ( .A1(n67971), .A2(n62522), .B1(n68166), .B2(n67964), .ZN(
        n7011) );
  OAI22_X1 U47559 ( .A1(n67971), .A2(n62521), .B1(n68169), .B2(n67964), .ZN(
        n7012) );
  OAI22_X1 U47560 ( .A1(n67972), .A2(n62520), .B1(n68172), .B2(n67964), .ZN(
        n7013) );
  OAI22_X1 U47561 ( .A1(n67972), .A2(n62519), .B1(n68175), .B2(n67964), .ZN(
        n7014) );
  OAI22_X1 U47562 ( .A1(n67972), .A2(n62518), .B1(n68178), .B2(n67964), .ZN(
        n7015) );
  OAI22_X1 U47563 ( .A1(n67972), .A2(n62517), .B1(n68181), .B2(n67964), .ZN(
        n7016) );
  OAI22_X1 U47564 ( .A1(n67972), .A2(n62516), .B1(n68184), .B2(n67964), .ZN(
        n7017) );
  OAI22_X1 U47565 ( .A1(n67972), .A2(n62515), .B1(n68187), .B2(n67964), .ZN(
        n7018) );
  OAI22_X1 U47566 ( .A1(n67972), .A2(n62514), .B1(n68190), .B2(n67964), .ZN(
        n7019) );
  OAI22_X1 U47567 ( .A1(n67972), .A2(n62513), .B1(n68193), .B2(n67964), .ZN(
        n7020) );
  OAI22_X1 U47568 ( .A1(n67972), .A2(n62512), .B1(n68196), .B2(n67964), .ZN(
        n7021) );
  OAI22_X1 U47569 ( .A1(n67972), .A2(n62511), .B1(n68199), .B2(n67964), .ZN(
        n7022) );
  OAI22_X1 U47570 ( .A1(n67972), .A2(n62510), .B1(n68202), .B2(n67965), .ZN(
        n7023) );
  OAI22_X1 U47571 ( .A1(n67972), .A2(n62509), .B1(n68205), .B2(n67965), .ZN(
        n7024) );
  OAI22_X1 U47572 ( .A1(n67972), .A2(n62508), .B1(n68208), .B2(n67965), .ZN(
        n7025) );
  OAI22_X1 U47573 ( .A1(n67973), .A2(n62507), .B1(n68211), .B2(n67965), .ZN(
        n7026) );
  OAI22_X1 U47574 ( .A1(n67973), .A2(n62506), .B1(n68214), .B2(n67965), .ZN(
        n7027) );
  OAI22_X1 U47575 ( .A1(n67973), .A2(n62505), .B1(n68217), .B2(n67965), .ZN(
        n7028) );
  OAI22_X1 U47576 ( .A1(n67973), .A2(n62504), .B1(n68220), .B2(n67965), .ZN(
        n7029) );
  OAI22_X1 U47577 ( .A1(n67973), .A2(n62503), .B1(n68223), .B2(n67965), .ZN(
        n7030) );
  OAI22_X1 U47578 ( .A1(n67973), .A2(n62502), .B1(n68226), .B2(n67965), .ZN(
        n7031) );
  OAI22_X1 U47579 ( .A1(n67973), .A2(n62501), .B1(n68229), .B2(n67965), .ZN(
        n7032) );
  OAI22_X1 U47580 ( .A1(n67973), .A2(n62500), .B1(n68232), .B2(n67965), .ZN(
        n7033) );
  OAI22_X1 U47581 ( .A1(n67973), .A2(n62499), .B1(n68235), .B2(n67965), .ZN(
        n7034) );
  OAI22_X1 U47582 ( .A1(n67803), .A2(n63226), .B1(n68059), .B2(n67795), .ZN(
        n6143) );
  OAI22_X1 U47583 ( .A1(n67803), .A2(n63225), .B1(n68062), .B2(n67795), .ZN(
        n6144) );
  OAI22_X1 U47584 ( .A1(n67803), .A2(n63224), .B1(n68065), .B2(n67795), .ZN(
        n6145) );
  OAI22_X1 U47585 ( .A1(n67803), .A2(n63223), .B1(n68068), .B2(n67795), .ZN(
        n6146) );
  OAI22_X1 U47586 ( .A1(n67803), .A2(n63222), .B1(n68071), .B2(n67795), .ZN(
        n6147) );
  OAI22_X1 U47587 ( .A1(n67803), .A2(n63221), .B1(n68074), .B2(n67795), .ZN(
        n6148) );
  OAI22_X1 U47588 ( .A1(n67803), .A2(n63220), .B1(n68077), .B2(n67795), .ZN(
        n6149) );
  OAI22_X1 U47589 ( .A1(n67803), .A2(n63219), .B1(n68080), .B2(n67795), .ZN(
        n6150) );
  OAI22_X1 U47590 ( .A1(n67803), .A2(n63218), .B1(n68083), .B2(n67795), .ZN(
        n6151) );
  OAI22_X1 U47591 ( .A1(n67803), .A2(n63217), .B1(n68086), .B2(n67795), .ZN(
        n6152) );
  OAI22_X1 U47592 ( .A1(n67803), .A2(n63216), .B1(n68089), .B2(n67795), .ZN(
        n6153) );
  OAI22_X1 U47593 ( .A1(n67803), .A2(n63215), .B1(n68092), .B2(n67795), .ZN(
        n6154) );
  OAI22_X1 U47594 ( .A1(n67804), .A2(n63214), .B1(n68095), .B2(n67796), .ZN(
        n6155) );
  OAI22_X1 U47595 ( .A1(n67804), .A2(n63213), .B1(n68098), .B2(n67796), .ZN(
        n6156) );
  OAI22_X1 U47596 ( .A1(n67804), .A2(n63212), .B1(n68101), .B2(n67796), .ZN(
        n6157) );
  OAI22_X1 U47597 ( .A1(n67804), .A2(n63211), .B1(n68104), .B2(n67796), .ZN(
        n6158) );
  OAI22_X1 U47598 ( .A1(n67804), .A2(n63210), .B1(n68107), .B2(n67796), .ZN(
        n6159) );
  OAI22_X1 U47599 ( .A1(n67804), .A2(n63209), .B1(n68110), .B2(n67796), .ZN(
        n6160) );
  OAI22_X1 U47600 ( .A1(n67804), .A2(n63208), .B1(n68113), .B2(n67796), .ZN(
        n6161) );
  OAI22_X1 U47601 ( .A1(n67804), .A2(n63207), .B1(n68116), .B2(n67796), .ZN(
        n6162) );
  OAI22_X1 U47602 ( .A1(n67804), .A2(n63206), .B1(n68119), .B2(n67796), .ZN(
        n6163) );
  OAI22_X1 U47603 ( .A1(n67804), .A2(n63205), .B1(n68122), .B2(n67796), .ZN(
        n6164) );
  OAI22_X1 U47604 ( .A1(n67804), .A2(n63204), .B1(n68125), .B2(n67796), .ZN(
        n6165) );
  OAI22_X1 U47605 ( .A1(n67804), .A2(n63203), .B1(n68128), .B2(n67796), .ZN(
        n6166) );
  OAI22_X1 U47606 ( .A1(n67804), .A2(n63202), .B1(n68131), .B2(n67797), .ZN(
        n6167) );
  OAI22_X1 U47607 ( .A1(n67805), .A2(n63201), .B1(n68134), .B2(n67797), .ZN(
        n6168) );
  OAI22_X1 U47608 ( .A1(n67805), .A2(n63200), .B1(n68137), .B2(n67797), .ZN(
        n6169) );
  OAI22_X1 U47609 ( .A1(n67805), .A2(n63199), .B1(n68140), .B2(n67797), .ZN(
        n6170) );
  OAI22_X1 U47610 ( .A1(n67805), .A2(n63198), .B1(n68143), .B2(n67797), .ZN(
        n6171) );
  OAI22_X1 U47611 ( .A1(n67805), .A2(n63197), .B1(n68146), .B2(n67797), .ZN(
        n6172) );
  OAI22_X1 U47612 ( .A1(n67805), .A2(n63196), .B1(n68149), .B2(n67797), .ZN(
        n6173) );
  OAI22_X1 U47613 ( .A1(n67805), .A2(n63195), .B1(n68152), .B2(n67797), .ZN(
        n6174) );
  OAI22_X1 U47614 ( .A1(n67805), .A2(n63194), .B1(n68155), .B2(n67797), .ZN(
        n6175) );
  OAI22_X1 U47615 ( .A1(n67805), .A2(n63193), .B1(n68158), .B2(n67797), .ZN(
        n6176) );
  OAI22_X1 U47616 ( .A1(n67805), .A2(n63192), .B1(n68161), .B2(n67797), .ZN(
        n6177) );
  OAI22_X1 U47617 ( .A1(n67805), .A2(n63191), .B1(n68164), .B2(n67797), .ZN(
        n6178) );
  OAI22_X1 U47618 ( .A1(n67805), .A2(n63190), .B1(n68167), .B2(n67798), .ZN(
        n6179) );
  OAI22_X1 U47619 ( .A1(n67805), .A2(n63189), .B1(n68170), .B2(n67798), .ZN(
        n6180) );
  OAI22_X1 U47620 ( .A1(n67806), .A2(n63188), .B1(n68173), .B2(n67798), .ZN(
        n6181) );
  OAI22_X1 U47621 ( .A1(n67806), .A2(n63187), .B1(n68176), .B2(n67798), .ZN(
        n6182) );
  OAI22_X1 U47622 ( .A1(n67806), .A2(n63186), .B1(n68179), .B2(n67798), .ZN(
        n6183) );
  OAI22_X1 U47623 ( .A1(n67806), .A2(n63185), .B1(n68182), .B2(n67798), .ZN(
        n6184) );
  OAI22_X1 U47624 ( .A1(n67806), .A2(n63184), .B1(n68185), .B2(n67798), .ZN(
        n6185) );
  OAI22_X1 U47625 ( .A1(n67806), .A2(n63183), .B1(n68188), .B2(n67798), .ZN(
        n6186) );
  OAI22_X1 U47626 ( .A1(n67806), .A2(n63182), .B1(n68191), .B2(n67798), .ZN(
        n6187) );
  OAI22_X1 U47627 ( .A1(n67806), .A2(n63181), .B1(n68194), .B2(n67798), .ZN(
        n6188) );
  OAI22_X1 U47628 ( .A1(n67806), .A2(n63180), .B1(n68197), .B2(n67798), .ZN(
        n6189) );
  OAI22_X1 U47629 ( .A1(n67806), .A2(n63179), .B1(n68200), .B2(n67798), .ZN(
        n6190) );
  OAI22_X1 U47630 ( .A1(n67806), .A2(n63178), .B1(n68203), .B2(n67799), .ZN(
        n6191) );
  OAI22_X1 U47631 ( .A1(n67806), .A2(n63177), .B1(n68206), .B2(n67799), .ZN(
        n6192) );
  OAI22_X1 U47632 ( .A1(n67806), .A2(n63176), .B1(n68209), .B2(n67799), .ZN(
        n6193) );
  OAI22_X1 U47633 ( .A1(n67807), .A2(n63175), .B1(n68212), .B2(n67799), .ZN(
        n6194) );
  OAI22_X1 U47634 ( .A1(n67807), .A2(n63174), .B1(n68215), .B2(n67799), .ZN(
        n6195) );
  OAI22_X1 U47635 ( .A1(n67807), .A2(n63173), .B1(n68218), .B2(n67799), .ZN(
        n6196) );
  OAI22_X1 U47636 ( .A1(n67807), .A2(n63172), .B1(n68221), .B2(n67799), .ZN(
        n6197) );
  OAI22_X1 U47637 ( .A1(n67807), .A2(n63171), .B1(n68224), .B2(n67799), .ZN(
        n6198) );
  OAI22_X1 U47638 ( .A1(n67807), .A2(n63170), .B1(n68227), .B2(n67799), .ZN(
        n6199) );
  OAI22_X1 U47639 ( .A1(n67807), .A2(n63169), .B1(n68230), .B2(n67799), .ZN(
        n6200) );
  OAI22_X1 U47640 ( .A1(n67807), .A2(n63168), .B1(n68233), .B2(n67799), .ZN(
        n6201) );
  OAI22_X1 U47641 ( .A1(n67807), .A2(n63167), .B1(n68236), .B2(n67799), .ZN(
        n6202) );
  OAI22_X1 U47642 ( .A1(n67854), .A2(n63024), .B1(n68059), .B2(n67846), .ZN(
        n6399) );
  OAI22_X1 U47643 ( .A1(n67854), .A2(n63023), .B1(n68062), .B2(n67846), .ZN(
        n6400) );
  OAI22_X1 U47644 ( .A1(n67854), .A2(n63022), .B1(n68065), .B2(n67846), .ZN(
        n6401) );
  OAI22_X1 U47645 ( .A1(n67854), .A2(n63021), .B1(n68068), .B2(n67846), .ZN(
        n6402) );
  OAI22_X1 U47646 ( .A1(n67854), .A2(n63020), .B1(n68071), .B2(n67846), .ZN(
        n6403) );
  OAI22_X1 U47647 ( .A1(n67854), .A2(n63019), .B1(n68074), .B2(n67846), .ZN(
        n6404) );
  OAI22_X1 U47648 ( .A1(n67854), .A2(n63018), .B1(n68077), .B2(n67846), .ZN(
        n6405) );
  OAI22_X1 U47649 ( .A1(n67854), .A2(n63017), .B1(n68080), .B2(n67846), .ZN(
        n6406) );
  OAI22_X1 U47650 ( .A1(n67854), .A2(n63016), .B1(n68083), .B2(n67846), .ZN(
        n6407) );
  OAI22_X1 U47651 ( .A1(n67854), .A2(n63015), .B1(n68086), .B2(n67846), .ZN(
        n6408) );
  OAI22_X1 U47652 ( .A1(n67854), .A2(n63014), .B1(n68089), .B2(n67846), .ZN(
        n6409) );
  OAI22_X1 U47653 ( .A1(n67854), .A2(n63013), .B1(n68092), .B2(n67846), .ZN(
        n6410) );
  OAI22_X1 U47654 ( .A1(n67855), .A2(n63012), .B1(n68095), .B2(n67847), .ZN(
        n6411) );
  OAI22_X1 U47655 ( .A1(n67855), .A2(n63011), .B1(n68098), .B2(n67847), .ZN(
        n6412) );
  OAI22_X1 U47656 ( .A1(n67855), .A2(n63010), .B1(n68101), .B2(n67847), .ZN(
        n6413) );
  OAI22_X1 U47657 ( .A1(n67855), .A2(n63009), .B1(n68104), .B2(n67847), .ZN(
        n6414) );
  OAI22_X1 U47658 ( .A1(n67855), .A2(n63008), .B1(n68107), .B2(n67847), .ZN(
        n6415) );
  OAI22_X1 U47659 ( .A1(n67855), .A2(n63007), .B1(n68110), .B2(n67847), .ZN(
        n6416) );
  OAI22_X1 U47660 ( .A1(n67855), .A2(n63006), .B1(n68113), .B2(n67847), .ZN(
        n6417) );
  OAI22_X1 U47661 ( .A1(n67855), .A2(n63005), .B1(n68116), .B2(n67847), .ZN(
        n6418) );
  OAI22_X1 U47662 ( .A1(n67855), .A2(n63004), .B1(n68119), .B2(n67847), .ZN(
        n6419) );
  OAI22_X1 U47663 ( .A1(n67855), .A2(n63003), .B1(n68122), .B2(n67847), .ZN(
        n6420) );
  OAI22_X1 U47664 ( .A1(n67855), .A2(n63002), .B1(n68125), .B2(n67847), .ZN(
        n6421) );
  OAI22_X1 U47665 ( .A1(n67855), .A2(n63001), .B1(n68128), .B2(n67847), .ZN(
        n6422) );
  OAI22_X1 U47666 ( .A1(n67855), .A2(n63000), .B1(n68131), .B2(n67848), .ZN(
        n6423) );
  OAI22_X1 U47667 ( .A1(n67856), .A2(n62999), .B1(n68134), .B2(n67848), .ZN(
        n6424) );
  OAI22_X1 U47668 ( .A1(n67856), .A2(n62998), .B1(n68137), .B2(n67848), .ZN(
        n6425) );
  OAI22_X1 U47669 ( .A1(n67856), .A2(n62997), .B1(n68140), .B2(n67848), .ZN(
        n6426) );
  OAI22_X1 U47670 ( .A1(n67856), .A2(n62996), .B1(n68143), .B2(n67848), .ZN(
        n6427) );
  OAI22_X1 U47671 ( .A1(n67856), .A2(n62995), .B1(n68146), .B2(n67848), .ZN(
        n6428) );
  OAI22_X1 U47672 ( .A1(n67856), .A2(n62994), .B1(n68149), .B2(n67848), .ZN(
        n6429) );
  OAI22_X1 U47673 ( .A1(n67856), .A2(n62993), .B1(n68152), .B2(n67848), .ZN(
        n6430) );
  OAI22_X1 U47674 ( .A1(n67856), .A2(n62992), .B1(n68155), .B2(n67848), .ZN(
        n6431) );
  OAI22_X1 U47675 ( .A1(n67856), .A2(n62991), .B1(n68158), .B2(n67848), .ZN(
        n6432) );
  OAI22_X1 U47676 ( .A1(n67856), .A2(n62990), .B1(n68161), .B2(n67848), .ZN(
        n6433) );
  OAI22_X1 U47677 ( .A1(n67856), .A2(n62989), .B1(n68164), .B2(n67848), .ZN(
        n6434) );
  OAI22_X1 U47678 ( .A1(n67856), .A2(n62988), .B1(n68167), .B2(n67849), .ZN(
        n6435) );
  OAI22_X1 U47679 ( .A1(n67856), .A2(n62987), .B1(n68170), .B2(n67849), .ZN(
        n6436) );
  OAI22_X1 U47680 ( .A1(n67857), .A2(n62986), .B1(n68173), .B2(n67849), .ZN(
        n6437) );
  OAI22_X1 U47681 ( .A1(n67857), .A2(n62985), .B1(n68176), .B2(n67849), .ZN(
        n6438) );
  OAI22_X1 U47682 ( .A1(n67857), .A2(n62984), .B1(n68179), .B2(n67849), .ZN(
        n6439) );
  OAI22_X1 U47683 ( .A1(n67857), .A2(n62983), .B1(n68182), .B2(n67849), .ZN(
        n6440) );
  OAI22_X1 U47684 ( .A1(n67857), .A2(n62982), .B1(n68185), .B2(n67849), .ZN(
        n6441) );
  OAI22_X1 U47685 ( .A1(n67857), .A2(n62981), .B1(n68188), .B2(n67849), .ZN(
        n6442) );
  OAI22_X1 U47686 ( .A1(n67857), .A2(n62980), .B1(n68191), .B2(n67849), .ZN(
        n6443) );
  OAI22_X1 U47687 ( .A1(n67857), .A2(n62979), .B1(n68194), .B2(n67849), .ZN(
        n6444) );
  OAI22_X1 U47688 ( .A1(n67857), .A2(n62978), .B1(n68197), .B2(n67849), .ZN(
        n6445) );
  OAI22_X1 U47689 ( .A1(n67857), .A2(n62977), .B1(n68200), .B2(n67849), .ZN(
        n6446) );
  OAI22_X1 U47690 ( .A1(n67857), .A2(n62976), .B1(n68203), .B2(n67850), .ZN(
        n6447) );
  OAI22_X1 U47691 ( .A1(n67857), .A2(n62975), .B1(n68206), .B2(n67850), .ZN(
        n6448) );
  OAI22_X1 U47692 ( .A1(n67857), .A2(n62974), .B1(n68209), .B2(n67850), .ZN(
        n6449) );
  OAI22_X1 U47693 ( .A1(n67858), .A2(n62973), .B1(n68212), .B2(n67850), .ZN(
        n6450) );
  OAI22_X1 U47694 ( .A1(n67858), .A2(n62972), .B1(n68215), .B2(n67850), .ZN(
        n6451) );
  OAI22_X1 U47695 ( .A1(n67858), .A2(n62971), .B1(n68218), .B2(n67850), .ZN(
        n6452) );
  OAI22_X1 U47696 ( .A1(n67858), .A2(n62970), .B1(n68221), .B2(n67850), .ZN(
        n6453) );
  OAI22_X1 U47697 ( .A1(n67858), .A2(n62969), .B1(n68224), .B2(n67850), .ZN(
        n6454) );
  OAI22_X1 U47698 ( .A1(n67858), .A2(n62968), .B1(n68227), .B2(n67850), .ZN(
        n6455) );
  OAI22_X1 U47699 ( .A1(n67858), .A2(n62967), .B1(n68230), .B2(n67850), .ZN(
        n6456) );
  OAI22_X1 U47700 ( .A1(n67858), .A2(n62966), .B1(n68233), .B2(n67850), .ZN(
        n6457) );
  OAI22_X1 U47701 ( .A1(n67858), .A2(n62965), .B1(n68236), .B2(n67850), .ZN(
        n6458) );
  OAI22_X1 U47702 ( .A1(n67841), .A2(n63091), .B1(n68059), .B2(n67833), .ZN(
        n6335) );
  OAI22_X1 U47703 ( .A1(n67841), .A2(n63090), .B1(n68062), .B2(n67833), .ZN(
        n6336) );
  OAI22_X1 U47704 ( .A1(n67841), .A2(n63089), .B1(n68065), .B2(n67833), .ZN(
        n6337) );
  OAI22_X1 U47705 ( .A1(n67841), .A2(n63088), .B1(n68068), .B2(n67833), .ZN(
        n6338) );
  OAI22_X1 U47706 ( .A1(n67841), .A2(n63087), .B1(n68071), .B2(n67833), .ZN(
        n6339) );
  OAI22_X1 U47707 ( .A1(n67841), .A2(n63086), .B1(n68074), .B2(n67833), .ZN(
        n6340) );
  OAI22_X1 U47708 ( .A1(n67841), .A2(n63085), .B1(n68077), .B2(n67833), .ZN(
        n6341) );
  OAI22_X1 U47709 ( .A1(n67841), .A2(n63084), .B1(n68080), .B2(n67833), .ZN(
        n6342) );
  OAI22_X1 U47710 ( .A1(n67841), .A2(n63083), .B1(n68083), .B2(n67833), .ZN(
        n6343) );
  OAI22_X1 U47711 ( .A1(n67841), .A2(n63082), .B1(n68086), .B2(n67833), .ZN(
        n6344) );
  OAI22_X1 U47712 ( .A1(n67841), .A2(n63081), .B1(n68089), .B2(n67833), .ZN(
        n6345) );
  OAI22_X1 U47713 ( .A1(n67841), .A2(n63080), .B1(n68092), .B2(n67833), .ZN(
        n6346) );
  OAI22_X1 U47714 ( .A1(n67842), .A2(n63079), .B1(n68095), .B2(n67834), .ZN(
        n6347) );
  OAI22_X1 U47715 ( .A1(n67842), .A2(n63078), .B1(n68098), .B2(n67834), .ZN(
        n6348) );
  OAI22_X1 U47716 ( .A1(n67842), .A2(n63077), .B1(n68101), .B2(n67834), .ZN(
        n6349) );
  OAI22_X1 U47717 ( .A1(n67842), .A2(n63076), .B1(n68104), .B2(n67834), .ZN(
        n6350) );
  OAI22_X1 U47718 ( .A1(n67842), .A2(n63075), .B1(n68107), .B2(n67834), .ZN(
        n6351) );
  OAI22_X1 U47719 ( .A1(n67842), .A2(n63074), .B1(n68110), .B2(n67834), .ZN(
        n6352) );
  OAI22_X1 U47720 ( .A1(n67842), .A2(n63073), .B1(n68113), .B2(n67834), .ZN(
        n6353) );
  OAI22_X1 U47721 ( .A1(n67842), .A2(n63072), .B1(n68116), .B2(n67834), .ZN(
        n6354) );
  OAI22_X1 U47722 ( .A1(n67842), .A2(n63071), .B1(n68119), .B2(n67834), .ZN(
        n6355) );
  OAI22_X1 U47723 ( .A1(n67842), .A2(n63070), .B1(n68122), .B2(n67834), .ZN(
        n6356) );
  OAI22_X1 U47724 ( .A1(n67842), .A2(n63069), .B1(n68125), .B2(n67834), .ZN(
        n6357) );
  OAI22_X1 U47725 ( .A1(n67842), .A2(n63068), .B1(n68128), .B2(n67834), .ZN(
        n6358) );
  OAI22_X1 U47726 ( .A1(n67842), .A2(n63067), .B1(n68131), .B2(n67835), .ZN(
        n6359) );
  OAI22_X1 U47727 ( .A1(n67843), .A2(n63066), .B1(n68134), .B2(n67835), .ZN(
        n6360) );
  OAI22_X1 U47728 ( .A1(n67843), .A2(n63065), .B1(n68137), .B2(n67835), .ZN(
        n6361) );
  OAI22_X1 U47729 ( .A1(n67843), .A2(n63064), .B1(n68140), .B2(n67835), .ZN(
        n6362) );
  OAI22_X1 U47730 ( .A1(n67843), .A2(n63063), .B1(n68143), .B2(n67835), .ZN(
        n6363) );
  OAI22_X1 U47731 ( .A1(n67843), .A2(n63062), .B1(n68146), .B2(n67835), .ZN(
        n6364) );
  OAI22_X1 U47732 ( .A1(n67843), .A2(n63061), .B1(n68149), .B2(n67835), .ZN(
        n6365) );
  OAI22_X1 U47733 ( .A1(n67843), .A2(n63060), .B1(n68152), .B2(n67835), .ZN(
        n6366) );
  OAI22_X1 U47734 ( .A1(n67843), .A2(n63059), .B1(n68155), .B2(n67835), .ZN(
        n6367) );
  OAI22_X1 U47735 ( .A1(n67843), .A2(n63058), .B1(n68158), .B2(n67835), .ZN(
        n6368) );
  OAI22_X1 U47736 ( .A1(n67843), .A2(n63057), .B1(n68161), .B2(n67835), .ZN(
        n6369) );
  OAI22_X1 U47737 ( .A1(n67843), .A2(n63056), .B1(n68164), .B2(n67835), .ZN(
        n6370) );
  OAI22_X1 U47738 ( .A1(n67843), .A2(n63055), .B1(n68167), .B2(n67836), .ZN(
        n6371) );
  OAI22_X1 U47739 ( .A1(n67843), .A2(n63054), .B1(n68170), .B2(n67836), .ZN(
        n6372) );
  OAI22_X1 U47740 ( .A1(n67844), .A2(n63053), .B1(n68173), .B2(n67836), .ZN(
        n6373) );
  OAI22_X1 U47741 ( .A1(n67844), .A2(n63052), .B1(n68176), .B2(n67836), .ZN(
        n6374) );
  OAI22_X1 U47742 ( .A1(n67844), .A2(n63051), .B1(n68179), .B2(n67836), .ZN(
        n6375) );
  OAI22_X1 U47743 ( .A1(n67844), .A2(n63050), .B1(n68182), .B2(n67836), .ZN(
        n6376) );
  OAI22_X1 U47744 ( .A1(n67844), .A2(n63049), .B1(n68185), .B2(n67836), .ZN(
        n6377) );
  OAI22_X1 U47745 ( .A1(n67844), .A2(n63048), .B1(n68188), .B2(n67836), .ZN(
        n6378) );
  OAI22_X1 U47746 ( .A1(n67844), .A2(n63047), .B1(n68191), .B2(n67836), .ZN(
        n6379) );
  OAI22_X1 U47747 ( .A1(n67844), .A2(n63046), .B1(n68194), .B2(n67836), .ZN(
        n6380) );
  OAI22_X1 U47748 ( .A1(n67844), .A2(n63045), .B1(n68197), .B2(n67836), .ZN(
        n6381) );
  OAI22_X1 U47749 ( .A1(n67844), .A2(n63044), .B1(n68200), .B2(n67836), .ZN(
        n6382) );
  OAI22_X1 U47750 ( .A1(n67844), .A2(n63043), .B1(n68203), .B2(n67837), .ZN(
        n6383) );
  OAI22_X1 U47751 ( .A1(n67844), .A2(n63042), .B1(n68206), .B2(n67837), .ZN(
        n6384) );
  OAI22_X1 U47752 ( .A1(n67844), .A2(n63041), .B1(n68209), .B2(n67837), .ZN(
        n6385) );
  OAI22_X1 U47753 ( .A1(n67845), .A2(n63040), .B1(n68212), .B2(n67837), .ZN(
        n6386) );
  OAI22_X1 U47754 ( .A1(n67845), .A2(n63039), .B1(n68215), .B2(n67837), .ZN(
        n6387) );
  OAI22_X1 U47755 ( .A1(n67845), .A2(n63038), .B1(n68218), .B2(n67837), .ZN(
        n6388) );
  OAI22_X1 U47756 ( .A1(n67845), .A2(n63037), .B1(n68221), .B2(n67837), .ZN(
        n6389) );
  OAI22_X1 U47757 ( .A1(n67845), .A2(n63036), .B1(n68224), .B2(n67837), .ZN(
        n6390) );
  OAI22_X1 U47758 ( .A1(n67845), .A2(n63035), .B1(n68227), .B2(n67837), .ZN(
        n6391) );
  OAI22_X1 U47759 ( .A1(n67845), .A2(n63034), .B1(n68230), .B2(n67837), .ZN(
        n6392) );
  OAI22_X1 U47760 ( .A1(n67845), .A2(n63033), .B1(n68233), .B2(n67837), .ZN(
        n6393) );
  OAI22_X1 U47761 ( .A1(n67845), .A2(n63032), .B1(n68236), .B2(n67837), .ZN(
        n6394) );
  OAI22_X1 U47762 ( .A1(n67752), .A2(n63427), .B1(n68059), .B2(n67744), .ZN(
        n5887) );
  OAI22_X1 U47763 ( .A1(n67752), .A2(n63426), .B1(n68062), .B2(n67744), .ZN(
        n5888) );
  OAI22_X1 U47764 ( .A1(n67752), .A2(n63425), .B1(n68065), .B2(n67744), .ZN(
        n5889) );
  OAI22_X1 U47765 ( .A1(n67752), .A2(n63424), .B1(n68068), .B2(n67744), .ZN(
        n5890) );
  OAI22_X1 U47766 ( .A1(n67752), .A2(n63423), .B1(n68071), .B2(n67744), .ZN(
        n5891) );
  OAI22_X1 U47767 ( .A1(n67752), .A2(n63422), .B1(n68074), .B2(n67744), .ZN(
        n5892) );
  OAI22_X1 U47768 ( .A1(n67752), .A2(n63421), .B1(n68077), .B2(n67744), .ZN(
        n5893) );
  OAI22_X1 U47769 ( .A1(n67752), .A2(n63420), .B1(n68080), .B2(n67744), .ZN(
        n5894) );
  OAI22_X1 U47770 ( .A1(n67752), .A2(n63419), .B1(n68083), .B2(n67744), .ZN(
        n5895) );
  OAI22_X1 U47771 ( .A1(n67752), .A2(n63418), .B1(n68086), .B2(n67744), .ZN(
        n5896) );
  OAI22_X1 U47772 ( .A1(n67752), .A2(n63417), .B1(n68089), .B2(n67744), .ZN(
        n5897) );
  OAI22_X1 U47773 ( .A1(n67752), .A2(n63416), .B1(n68092), .B2(n67744), .ZN(
        n5898) );
  OAI22_X1 U47774 ( .A1(n67753), .A2(n63415), .B1(n68095), .B2(n67745), .ZN(
        n5899) );
  OAI22_X1 U47775 ( .A1(n67753), .A2(n63414), .B1(n68098), .B2(n67745), .ZN(
        n5900) );
  OAI22_X1 U47776 ( .A1(n67753), .A2(n63413), .B1(n68101), .B2(n67745), .ZN(
        n5901) );
  OAI22_X1 U47777 ( .A1(n67753), .A2(n63412), .B1(n68104), .B2(n67745), .ZN(
        n5902) );
  OAI22_X1 U47778 ( .A1(n67753), .A2(n63411), .B1(n68107), .B2(n67745), .ZN(
        n5903) );
  OAI22_X1 U47779 ( .A1(n67753), .A2(n63410), .B1(n68110), .B2(n67745), .ZN(
        n5904) );
  OAI22_X1 U47780 ( .A1(n67753), .A2(n63409), .B1(n68113), .B2(n67745), .ZN(
        n5905) );
  OAI22_X1 U47781 ( .A1(n67753), .A2(n63408), .B1(n68116), .B2(n67745), .ZN(
        n5906) );
  OAI22_X1 U47782 ( .A1(n67753), .A2(n63407), .B1(n68119), .B2(n67745), .ZN(
        n5907) );
  OAI22_X1 U47783 ( .A1(n67753), .A2(n63406), .B1(n68122), .B2(n67745), .ZN(
        n5908) );
  OAI22_X1 U47784 ( .A1(n67753), .A2(n63405), .B1(n68125), .B2(n67745), .ZN(
        n5909) );
  OAI22_X1 U47785 ( .A1(n67753), .A2(n63404), .B1(n68128), .B2(n67745), .ZN(
        n5910) );
  OAI22_X1 U47786 ( .A1(n67753), .A2(n63403), .B1(n68131), .B2(n67746), .ZN(
        n5911) );
  OAI22_X1 U47787 ( .A1(n67754), .A2(n63402), .B1(n68134), .B2(n67746), .ZN(
        n5912) );
  OAI22_X1 U47788 ( .A1(n67754), .A2(n63401), .B1(n68137), .B2(n67746), .ZN(
        n5913) );
  OAI22_X1 U47789 ( .A1(n67754), .A2(n63400), .B1(n68140), .B2(n67746), .ZN(
        n5914) );
  OAI22_X1 U47790 ( .A1(n67754), .A2(n63399), .B1(n68143), .B2(n67746), .ZN(
        n5915) );
  OAI22_X1 U47791 ( .A1(n67754), .A2(n63398), .B1(n68146), .B2(n67746), .ZN(
        n5916) );
  OAI22_X1 U47792 ( .A1(n67754), .A2(n63397), .B1(n68149), .B2(n67746), .ZN(
        n5917) );
  OAI22_X1 U47793 ( .A1(n67754), .A2(n63396), .B1(n68152), .B2(n67746), .ZN(
        n5918) );
  OAI22_X1 U47794 ( .A1(n67754), .A2(n63395), .B1(n68155), .B2(n67746), .ZN(
        n5919) );
  OAI22_X1 U47795 ( .A1(n67754), .A2(n63394), .B1(n68158), .B2(n67746), .ZN(
        n5920) );
  OAI22_X1 U47796 ( .A1(n67754), .A2(n63393), .B1(n68161), .B2(n67746), .ZN(
        n5921) );
  OAI22_X1 U47797 ( .A1(n67754), .A2(n63392), .B1(n68164), .B2(n67746), .ZN(
        n5922) );
  OAI22_X1 U47798 ( .A1(n67754), .A2(n63391), .B1(n68167), .B2(n67747), .ZN(
        n5923) );
  OAI22_X1 U47799 ( .A1(n67754), .A2(n63390), .B1(n68170), .B2(n67747), .ZN(
        n5924) );
  OAI22_X1 U47800 ( .A1(n67755), .A2(n63389), .B1(n68173), .B2(n67747), .ZN(
        n5925) );
  OAI22_X1 U47801 ( .A1(n67755), .A2(n63388), .B1(n68176), .B2(n67747), .ZN(
        n5926) );
  OAI22_X1 U47802 ( .A1(n67755), .A2(n63387), .B1(n68179), .B2(n67747), .ZN(
        n5927) );
  OAI22_X1 U47803 ( .A1(n67755), .A2(n63386), .B1(n68182), .B2(n67747), .ZN(
        n5928) );
  OAI22_X1 U47804 ( .A1(n67755), .A2(n63385), .B1(n68185), .B2(n67747), .ZN(
        n5929) );
  OAI22_X1 U47805 ( .A1(n67755), .A2(n63384), .B1(n68188), .B2(n67747), .ZN(
        n5930) );
  OAI22_X1 U47806 ( .A1(n67755), .A2(n63383), .B1(n68191), .B2(n67747), .ZN(
        n5931) );
  OAI22_X1 U47807 ( .A1(n67755), .A2(n63382), .B1(n68194), .B2(n67747), .ZN(
        n5932) );
  OAI22_X1 U47808 ( .A1(n67755), .A2(n63381), .B1(n68197), .B2(n67747), .ZN(
        n5933) );
  OAI22_X1 U47809 ( .A1(n67755), .A2(n63380), .B1(n68200), .B2(n67747), .ZN(
        n5934) );
  OAI22_X1 U47810 ( .A1(n67755), .A2(n63379), .B1(n68203), .B2(n67748), .ZN(
        n5935) );
  OAI22_X1 U47811 ( .A1(n67755), .A2(n63378), .B1(n68206), .B2(n67748), .ZN(
        n5936) );
  OAI22_X1 U47812 ( .A1(n67755), .A2(n63377), .B1(n68209), .B2(n67748), .ZN(
        n5937) );
  OAI22_X1 U47813 ( .A1(n67756), .A2(n63376), .B1(n68212), .B2(n67748), .ZN(
        n5938) );
  OAI22_X1 U47814 ( .A1(n67756), .A2(n63375), .B1(n68215), .B2(n67748), .ZN(
        n5939) );
  OAI22_X1 U47815 ( .A1(n67756), .A2(n63374), .B1(n68218), .B2(n67748), .ZN(
        n5940) );
  OAI22_X1 U47816 ( .A1(n67756), .A2(n63373), .B1(n68221), .B2(n67748), .ZN(
        n5941) );
  OAI22_X1 U47817 ( .A1(n67756), .A2(n63372), .B1(n68224), .B2(n67748), .ZN(
        n5942) );
  OAI22_X1 U47818 ( .A1(n67756), .A2(n63371), .B1(n68227), .B2(n67748), .ZN(
        n5943) );
  OAI22_X1 U47819 ( .A1(n67756), .A2(n63370), .B1(n68230), .B2(n67748), .ZN(
        n5944) );
  OAI22_X1 U47820 ( .A1(n67756), .A2(n63369), .B1(n68233), .B2(n67748), .ZN(
        n5945) );
  OAI22_X1 U47821 ( .A1(n67756), .A2(n63368), .B1(n68236), .B2(n67748), .ZN(
        n5946) );
  OAI22_X1 U47822 ( .A1(n67880), .A2(n62891), .B1(n68059), .B2(n67872), .ZN(
        n6527) );
  OAI22_X1 U47823 ( .A1(n67880), .A2(n62890), .B1(n68062), .B2(n67872), .ZN(
        n6528) );
  OAI22_X1 U47824 ( .A1(n67880), .A2(n62889), .B1(n68065), .B2(n67872), .ZN(
        n6529) );
  OAI22_X1 U47825 ( .A1(n67880), .A2(n62888), .B1(n68068), .B2(n67872), .ZN(
        n6530) );
  OAI22_X1 U47826 ( .A1(n67880), .A2(n62887), .B1(n68071), .B2(n67872), .ZN(
        n6531) );
  OAI22_X1 U47827 ( .A1(n67880), .A2(n62886), .B1(n68074), .B2(n67872), .ZN(
        n6532) );
  OAI22_X1 U47828 ( .A1(n67880), .A2(n62885), .B1(n68077), .B2(n67872), .ZN(
        n6533) );
  OAI22_X1 U47829 ( .A1(n67880), .A2(n62884), .B1(n68080), .B2(n67872), .ZN(
        n6534) );
  OAI22_X1 U47830 ( .A1(n67880), .A2(n62883), .B1(n68083), .B2(n67872), .ZN(
        n6535) );
  OAI22_X1 U47831 ( .A1(n67880), .A2(n62882), .B1(n68086), .B2(n67872), .ZN(
        n6536) );
  OAI22_X1 U47832 ( .A1(n67880), .A2(n62881), .B1(n68089), .B2(n67872), .ZN(
        n6537) );
  OAI22_X1 U47833 ( .A1(n67880), .A2(n62880), .B1(n68092), .B2(n67872), .ZN(
        n6538) );
  OAI22_X1 U47834 ( .A1(n67881), .A2(n62879), .B1(n68095), .B2(n67873), .ZN(
        n6539) );
  OAI22_X1 U47835 ( .A1(n67881), .A2(n62878), .B1(n68098), .B2(n67873), .ZN(
        n6540) );
  OAI22_X1 U47836 ( .A1(n67881), .A2(n62877), .B1(n68101), .B2(n67873), .ZN(
        n6541) );
  OAI22_X1 U47837 ( .A1(n67881), .A2(n62876), .B1(n68104), .B2(n67873), .ZN(
        n6542) );
  OAI22_X1 U47838 ( .A1(n67881), .A2(n62875), .B1(n68107), .B2(n67873), .ZN(
        n6543) );
  OAI22_X1 U47839 ( .A1(n67881), .A2(n62874), .B1(n68110), .B2(n67873), .ZN(
        n6544) );
  OAI22_X1 U47840 ( .A1(n67881), .A2(n62873), .B1(n68113), .B2(n67873), .ZN(
        n6545) );
  OAI22_X1 U47841 ( .A1(n67881), .A2(n62872), .B1(n68116), .B2(n67873), .ZN(
        n6546) );
  OAI22_X1 U47842 ( .A1(n67881), .A2(n62871), .B1(n68119), .B2(n67873), .ZN(
        n6547) );
  OAI22_X1 U47843 ( .A1(n67881), .A2(n62870), .B1(n68122), .B2(n67873), .ZN(
        n6548) );
  OAI22_X1 U47844 ( .A1(n67881), .A2(n62869), .B1(n68125), .B2(n67873), .ZN(
        n6549) );
  OAI22_X1 U47845 ( .A1(n67881), .A2(n62868), .B1(n68128), .B2(n67873), .ZN(
        n6550) );
  OAI22_X1 U47846 ( .A1(n67881), .A2(n62867), .B1(n68131), .B2(n67874), .ZN(
        n6551) );
  OAI22_X1 U47847 ( .A1(n67882), .A2(n62866), .B1(n68134), .B2(n67874), .ZN(
        n6552) );
  OAI22_X1 U47848 ( .A1(n67882), .A2(n62865), .B1(n68137), .B2(n67874), .ZN(
        n6553) );
  OAI22_X1 U47849 ( .A1(n67882), .A2(n62864), .B1(n68140), .B2(n67874), .ZN(
        n6554) );
  OAI22_X1 U47850 ( .A1(n67882), .A2(n62863), .B1(n68143), .B2(n67874), .ZN(
        n6555) );
  OAI22_X1 U47851 ( .A1(n67882), .A2(n62862), .B1(n68146), .B2(n67874), .ZN(
        n6556) );
  OAI22_X1 U47852 ( .A1(n67882), .A2(n62861), .B1(n68149), .B2(n67874), .ZN(
        n6557) );
  OAI22_X1 U47853 ( .A1(n67882), .A2(n62860), .B1(n68152), .B2(n67874), .ZN(
        n6558) );
  OAI22_X1 U47854 ( .A1(n67882), .A2(n62859), .B1(n68155), .B2(n67874), .ZN(
        n6559) );
  OAI22_X1 U47855 ( .A1(n67882), .A2(n62858), .B1(n68158), .B2(n67874), .ZN(
        n6560) );
  OAI22_X1 U47856 ( .A1(n67882), .A2(n62857), .B1(n68161), .B2(n67874), .ZN(
        n6561) );
  OAI22_X1 U47857 ( .A1(n67882), .A2(n62856), .B1(n68164), .B2(n67874), .ZN(
        n6562) );
  OAI22_X1 U47858 ( .A1(n67882), .A2(n62855), .B1(n68167), .B2(n67875), .ZN(
        n6563) );
  OAI22_X1 U47859 ( .A1(n67882), .A2(n62854), .B1(n68170), .B2(n67875), .ZN(
        n6564) );
  OAI22_X1 U47860 ( .A1(n67883), .A2(n62853), .B1(n68173), .B2(n67875), .ZN(
        n6565) );
  OAI22_X1 U47861 ( .A1(n67883), .A2(n62852), .B1(n68176), .B2(n67875), .ZN(
        n6566) );
  OAI22_X1 U47862 ( .A1(n67883), .A2(n62851), .B1(n68179), .B2(n67875), .ZN(
        n6567) );
  OAI22_X1 U47863 ( .A1(n67883), .A2(n62850), .B1(n68182), .B2(n67875), .ZN(
        n6568) );
  OAI22_X1 U47864 ( .A1(n67883), .A2(n62849), .B1(n68185), .B2(n67875), .ZN(
        n6569) );
  OAI22_X1 U47865 ( .A1(n67883), .A2(n62848), .B1(n68188), .B2(n67875), .ZN(
        n6570) );
  OAI22_X1 U47866 ( .A1(n67883), .A2(n62847), .B1(n68191), .B2(n67875), .ZN(
        n6571) );
  OAI22_X1 U47867 ( .A1(n67883), .A2(n62846), .B1(n68194), .B2(n67875), .ZN(
        n6572) );
  OAI22_X1 U47868 ( .A1(n67883), .A2(n62845), .B1(n68197), .B2(n67875), .ZN(
        n6573) );
  OAI22_X1 U47869 ( .A1(n67883), .A2(n62844), .B1(n68200), .B2(n67875), .ZN(
        n6574) );
  OAI22_X1 U47870 ( .A1(n67883), .A2(n62843), .B1(n68203), .B2(n67876), .ZN(
        n6575) );
  OAI22_X1 U47871 ( .A1(n67883), .A2(n62842), .B1(n68206), .B2(n67876), .ZN(
        n6576) );
  OAI22_X1 U47872 ( .A1(n67883), .A2(n62841), .B1(n68209), .B2(n67876), .ZN(
        n6577) );
  OAI22_X1 U47873 ( .A1(n67884), .A2(n62840), .B1(n68212), .B2(n67876), .ZN(
        n6578) );
  OAI22_X1 U47874 ( .A1(n67884), .A2(n62839), .B1(n68215), .B2(n67876), .ZN(
        n6579) );
  OAI22_X1 U47875 ( .A1(n67884), .A2(n62838), .B1(n68218), .B2(n67876), .ZN(
        n6580) );
  OAI22_X1 U47876 ( .A1(n67884), .A2(n62837), .B1(n68221), .B2(n67876), .ZN(
        n6581) );
  OAI22_X1 U47877 ( .A1(n67884), .A2(n62836), .B1(n68224), .B2(n67876), .ZN(
        n6582) );
  OAI22_X1 U47878 ( .A1(n67884), .A2(n62835), .B1(n68227), .B2(n67876), .ZN(
        n6583) );
  OAI22_X1 U47879 ( .A1(n67884), .A2(n62834), .B1(n68230), .B2(n67876), .ZN(
        n6584) );
  OAI22_X1 U47880 ( .A1(n67884), .A2(n62833), .B1(n68233), .B2(n67876), .ZN(
        n6585) );
  OAI22_X1 U47881 ( .A1(n67884), .A2(n62832), .B1(n68236), .B2(n67876), .ZN(
        n6586) );
  OAI22_X1 U47882 ( .A1(n68034), .A2(n62222), .B1(n68058), .B2(n68026), .ZN(
        n7295) );
  OAI22_X1 U47883 ( .A1(n68034), .A2(n62221), .B1(n68061), .B2(n68026), .ZN(
        n7296) );
  OAI22_X1 U47884 ( .A1(n68034), .A2(n62220), .B1(n68064), .B2(n68026), .ZN(
        n7297) );
  OAI22_X1 U47885 ( .A1(n68034), .A2(n62219), .B1(n68067), .B2(n68026), .ZN(
        n7298) );
  OAI22_X1 U47886 ( .A1(n68034), .A2(n62218), .B1(n68070), .B2(n68026), .ZN(
        n7299) );
  OAI22_X1 U47887 ( .A1(n68034), .A2(n62217), .B1(n68073), .B2(n68026), .ZN(
        n7300) );
  OAI22_X1 U47888 ( .A1(n68034), .A2(n62216), .B1(n68076), .B2(n68026), .ZN(
        n7301) );
  OAI22_X1 U47889 ( .A1(n68034), .A2(n62215), .B1(n68079), .B2(n68026), .ZN(
        n7302) );
  OAI22_X1 U47890 ( .A1(n68034), .A2(n62214), .B1(n68082), .B2(n68026), .ZN(
        n7303) );
  OAI22_X1 U47891 ( .A1(n68034), .A2(n62213), .B1(n68085), .B2(n68026), .ZN(
        n7304) );
  OAI22_X1 U47892 ( .A1(n68034), .A2(n62212), .B1(n68088), .B2(n68026), .ZN(
        n7305) );
  OAI22_X1 U47893 ( .A1(n68034), .A2(n62211), .B1(n68091), .B2(n68026), .ZN(
        n7306) );
  OAI22_X1 U47894 ( .A1(n68035), .A2(n62210), .B1(n68094), .B2(n68027), .ZN(
        n7307) );
  OAI22_X1 U47895 ( .A1(n68035), .A2(n62209), .B1(n68097), .B2(n68027), .ZN(
        n7308) );
  OAI22_X1 U47896 ( .A1(n68035), .A2(n62208), .B1(n68100), .B2(n68027), .ZN(
        n7309) );
  OAI22_X1 U47897 ( .A1(n68035), .A2(n62207), .B1(n68103), .B2(n68027), .ZN(
        n7310) );
  OAI22_X1 U47898 ( .A1(n68035), .A2(n62206), .B1(n68106), .B2(n68027), .ZN(
        n7311) );
  OAI22_X1 U47899 ( .A1(n68035), .A2(n62205), .B1(n68109), .B2(n68027), .ZN(
        n7312) );
  OAI22_X1 U47900 ( .A1(n68035), .A2(n62204), .B1(n68112), .B2(n68027), .ZN(
        n7313) );
  OAI22_X1 U47901 ( .A1(n68035), .A2(n62203), .B1(n68115), .B2(n68027), .ZN(
        n7314) );
  OAI22_X1 U47902 ( .A1(n68035), .A2(n62202), .B1(n68118), .B2(n68027), .ZN(
        n7315) );
  OAI22_X1 U47903 ( .A1(n68035), .A2(n62201), .B1(n68121), .B2(n68027), .ZN(
        n7316) );
  OAI22_X1 U47904 ( .A1(n68035), .A2(n62200), .B1(n68124), .B2(n68027), .ZN(
        n7317) );
  OAI22_X1 U47905 ( .A1(n68035), .A2(n62199), .B1(n68127), .B2(n68027), .ZN(
        n7318) );
  OAI22_X1 U47906 ( .A1(n68035), .A2(n62198), .B1(n68130), .B2(n68028), .ZN(
        n7319) );
  OAI22_X1 U47907 ( .A1(n68036), .A2(n62197), .B1(n68133), .B2(n68028), .ZN(
        n7320) );
  OAI22_X1 U47908 ( .A1(n68036), .A2(n62196), .B1(n68136), .B2(n68028), .ZN(
        n7321) );
  OAI22_X1 U47909 ( .A1(n68036), .A2(n62195), .B1(n68139), .B2(n68028), .ZN(
        n7322) );
  OAI22_X1 U47910 ( .A1(n68036), .A2(n62194), .B1(n68142), .B2(n68028), .ZN(
        n7323) );
  OAI22_X1 U47911 ( .A1(n68036), .A2(n62193), .B1(n68145), .B2(n68028), .ZN(
        n7324) );
  OAI22_X1 U47912 ( .A1(n68036), .A2(n62192), .B1(n68148), .B2(n68028), .ZN(
        n7325) );
  OAI22_X1 U47913 ( .A1(n68036), .A2(n62191), .B1(n68151), .B2(n68028), .ZN(
        n7326) );
  OAI22_X1 U47914 ( .A1(n68036), .A2(n62190), .B1(n68154), .B2(n68028), .ZN(
        n7327) );
  OAI22_X1 U47915 ( .A1(n68036), .A2(n62189), .B1(n68157), .B2(n68028), .ZN(
        n7328) );
  OAI22_X1 U47916 ( .A1(n68036), .A2(n62188), .B1(n68160), .B2(n68028), .ZN(
        n7329) );
  OAI22_X1 U47917 ( .A1(n68036), .A2(n62187), .B1(n68163), .B2(n68028), .ZN(
        n7330) );
  OAI22_X1 U47918 ( .A1(n68036), .A2(n62186), .B1(n68166), .B2(n68029), .ZN(
        n7331) );
  OAI22_X1 U47919 ( .A1(n68036), .A2(n62185), .B1(n68169), .B2(n68029), .ZN(
        n7332) );
  OAI22_X1 U47920 ( .A1(n68037), .A2(n62184), .B1(n68172), .B2(n68029), .ZN(
        n7333) );
  OAI22_X1 U47921 ( .A1(n68037), .A2(n62183), .B1(n68175), .B2(n68029), .ZN(
        n7334) );
  OAI22_X1 U47922 ( .A1(n68037), .A2(n62182), .B1(n68178), .B2(n68029), .ZN(
        n7335) );
  OAI22_X1 U47923 ( .A1(n68037), .A2(n62181), .B1(n68181), .B2(n68029), .ZN(
        n7336) );
  OAI22_X1 U47924 ( .A1(n68037), .A2(n62180), .B1(n68184), .B2(n68029), .ZN(
        n7337) );
  OAI22_X1 U47925 ( .A1(n68037), .A2(n62179), .B1(n68187), .B2(n68029), .ZN(
        n7338) );
  OAI22_X1 U47926 ( .A1(n68037), .A2(n62178), .B1(n68190), .B2(n68029), .ZN(
        n7339) );
  OAI22_X1 U47927 ( .A1(n68037), .A2(n62177), .B1(n68193), .B2(n68029), .ZN(
        n7340) );
  OAI22_X1 U47928 ( .A1(n68037), .A2(n62176), .B1(n68196), .B2(n68029), .ZN(
        n7341) );
  OAI22_X1 U47929 ( .A1(n68037), .A2(n62175), .B1(n68199), .B2(n68029), .ZN(
        n7342) );
  OAI22_X1 U47930 ( .A1(n68037), .A2(n62174), .B1(n68202), .B2(n68030), .ZN(
        n7343) );
  OAI22_X1 U47931 ( .A1(n68037), .A2(n62173), .B1(n68205), .B2(n68030), .ZN(
        n7344) );
  OAI22_X1 U47932 ( .A1(n68037), .A2(n62172), .B1(n68208), .B2(n68030), .ZN(
        n7345) );
  OAI22_X1 U47933 ( .A1(n68038), .A2(n62171), .B1(n68211), .B2(n68030), .ZN(
        n7346) );
  OAI22_X1 U47934 ( .A1(n68038), .A2(n62170), .B1(n68214), .B2(n68030), .ZN(
        n7347) );
  OAI22_X1 U47935 ( .A1(n68038), .A2(n62169), .B1(n68217), .B2(n68030), .ZN(
        n7348) );
  OAI22_X1 U47936 ( .A1(n68038), .A2(n62168), .B1(n68220), .B2(n68030), .ZN(
        n7349) );
  OAI22_X1 U47937 ( .A1(n68038), .A2(n62167), .B1(n68223), .B2(n68030), .ZN(
        n7350) );
  OAI22_X1 U47938 ( .A1(n68038), .A2(n62166), .B1(n68226), .B2(n68030), .ZN(
        n7351) );
  OAI22_X1 U47939 ( .A1(n68038), .A2(n62165), .B1(n68229), .B2(n68030), .ZN(
        n7352) );
  OAI22_X1 U47940 ( .A1(n68038), .A2(n62164), .B1(n68232), .B2(n68030), .ZN(
        n7353) );
  OAI22_X1 U47941 ( .A1(n68038), .A2(n62163), .B1(n68235), .B2(n68030), .ZN(
        n7354) );
  OAI22_X1 U47942 ( .A1(n68021), .A2(n62289), .B1(n68058), .B2(n68013), .ZN(
        n7231) );
  OAI22_X1 U47943 ( .A1(n68021), .A2(n62288), .B1(n68061), .B2(n68013), .ZN(
        n7232) );
  OAI22_X1 U47944 ( .A1(n68021), .A2(n62287), .B1(n68064), .B2(n68013), .ZN(
        n7233) );
  OAI22_X1 U47945 ( .A1(n68021), .A2(n62286), .B1(n68067), .B2(n68013), .ZN(
        n7234) );
  OAI22_X1 U47946 ( .A1(n68021), .A2(n62285), .B1(n68070), .B2(n68013), .ZN(
        n7235) );
  OAI22_X1 U47947 ( .A1(n68021), .A2(n62284), .B1(n68073), .B2(n68013), .ZN(
        n7236) );
  OAI22_X1 U47948 ( .A1(n68021), .A2(n62283), .B1(n68076), .B2(n68013), .ZN(
        n7237) );
  OAI22_X1 U47949 ( .A1(n68021), .A2(n62282), .B1(n68079), .B2(n68013), .ZN(
        n7238) );
  OAI22_X1 U47950 ( .A1(n68021), .A2(n62281), .B1(n68082), .B2(n68013), .ZN(
        n7239) );
  OAI22_X1 U47951 ( .A1(n68021), .A2(n62280), .B1(n68085), .B2(n68013), .ZN(
        n7240) );
  OAI22_X1 U47952 ( .A1(n68021), .A2(n62279), .B1(n68088), .B2(n68013), .ZN(
        n7241) );
  OAI22_X1 U47953 ( .A1(n68021), .A2(n62278), .B1(n68091), .B2(n68013), .ZN(
        n7242) );
  OAI22_X1 U47954 ( .A1(n68022), .A2(n62277), .B1(n68094), .B2(n68014), .ZN(
        n7243) );
  OAI22_X1 U47955 ( .A1(n68022), .A2(n62276), .B1(n68097), .B2(n68014), .ZN(
        n7244) );
  OAI22_X1 U47956 ( .A1(n68022), .A2(n62275), .B1(n68100), .B2(n68014), .ZN(
        n7245) );
  OAI22_X1 U47957 ( .A1(n68022), .A2(n62274), .B1(n68103), .B2(n68014), .ZN(
        n7246) );
  OAI22_X1 U47958 ( .A1(n68022), .A2(n62273), .B1(n68106), .B2(n68014), .ZN(
        n7247) );
  OAI22_X1 U47959 ( .A1(n68022), .A2(n62272), .B1(n68109), .B2(n68014), .ZN(
        n7248) );
  OAI22_X1 U47960 ( .A1(n68022), .A2(n62271), .B1(n68112), .B2(n68014), .ZN(
        n7249) );
  OAI22_X1 U47961 ( .A1(n68022), .A2(n62270), .B1(n68115), .B2(n68014), .ZN(
        n7250) );
  OAI22_X1 U47962 ( .A1(n68022), .A2(n62269), .B1(n68118), .B2(n68014), .ZN(
        n7251) );
  OAI22_X1 U47963 ( .A1(n68022), .A2(n62268), .B1(n68121), .B2(n68014), .ZN(
        n7252) );
  OAI22_X1 U47964 ( .A1(n68022), .A2(n62267), .B1(n68124), .B2(n68014), .ZN(
        n7253) );
  OAI22_X1 U47965 ( .A1(n68022), .A2(n62266), .B1(n68127), .B2(n68014), .ZN(
        n7254) );
  OAI22_X1 U47966 ( .A1(n68022), .A2(n62265), .B1(n68130), .B2(n68015), .ZN(
        n7255) );
  OAI22_X1 U47967 ( .A1(n68023), .A2(n62264), .B1(n68133), .B2(n68015), .ZN(
        n7256) );
  OAI22_X1 U47968 ( .A1(n68023), .A2(n62263), .B1(n68136), .B2(n68015), .ZN(
        n7257) );
  OAI22_X1 U47969 ( .A1(n68023), .A2(n62262), .B1(n68139), .B2(n68015), .ZN(
        n7258) );
  OAI22_X1 U47970 ( .A1(n68023), .A2(n62261), .B1(n68142), .B2(n68015), .ZN(
        n7259) );
  OAI22_X1 U47971 ( .A1(n68023), .A2(n62260), .B1(n68145), .B2(n68015), .ZN(
        n7260) );
  OAI22_X1 U47972 ( .A1(n68023), .A2(n62259), .B1(n68148), .B2(n68015), .ZN(
        n7261) );
  OAI22_X1 U47973 ( .A1(n68023), .A2(n62258), .B1(n68151), .B2(n68015), .ZN(
        n7262) );
  OAI22_X1 U47974 ( .A1(n68023), .A2(n62257), .B1(n68154), .B2(n68015), .ZN(
        n7263) );
  OAI22_X1 U47975 ( .A1(n68023), .A2(n62256), .B1(n68157), .B2(n68015), .ZN(
        n7264) );
  OAI22_X1 U47976 ( .A1(n68023), .A2(n62255), .B1(n68160), .B2(n68015), .ZN(
        n7265) );
  OAI22_X1 U47977 ( .A1(n68023), .A2(n62254), .B1(n68163), .B2(n68015), .ZN(
        n7266) );
  OAI22_X1 U47978 ( .A1(n68023), .A2(n62253), .B1(n68166), .B2(n68016), .ZN(
        n7267) );
  OAI22_X1 U47979 ( .A1(n68023), .A2(n62252), .B1(n68169), .B2(n68016), .ZN(
        n7268) );
  OAI22_X1 U47980 ( .A1(n68024), .A2(n62251), .B1(n68172), .B2(n68016), .ZN(
        n7269) );
  OAI22_X1 U47981 ( .A1(n68024), .A2(n62250), .B1(n68175), .B2(n68016), .ZN(
        n7270) );
  OAI22_X1 U47982 ( .A1(n68024), .A2(n62249), .B1(n68178), .B2(n68016), .ZN(
        n7271) );
  OAI22_X1 U47983 ( .A1(n68024), .A2(n62248), .B1(n68181), .B2(n68016), .ZN(
        n7272) );
  OAI22_X1 U47984 ( .A1(n68024), .A2(n62247), .B1(n68184), .B2(n68016), .ZN(
        n7273) );
  OAI22_X1 U47985 ( .A1(n68024), .A2(n62246), .B1(n68187), .B2(n68016), .ZN(
        n7274) );
  OAI22_X1 U47986 ( .A1(n68024), .A2(n62245), .B1(n68190), .B2(n68016), .ZN(
        n7275) );
  OAI22_X1 U47987 ( .A1(n68024), .A2(n62244), .B1(n68193), .B2(n68016), .ZN(
        n7276) );
  OAI22_X1 U47988 ( .A1(n68024), .A2(n62243), .B1(n68196), .B2(n68016), .ZN(
        n7277) );
  OAI22_X1 U47989 ( .A1(n68024), .A2(n62242), .B1(n68199), .B2(n68016), .ZN(
        n7278) );
  OAI22_X1 U47990 ( .A1(n68024), .A2(n62241), .B1(n68202), .B2(n68017), .ZN(
        n7279) );
  OAI22_X1 U47991 ( .A1(n68024), .A2(n62240), .B1(n68205), .B2(n68017), .ZN(
        n7280) );
  OAI22_X1 U47992 ( .A1(n68024), .A2(n62239), .B1(n68208), .B2(n68017), .ZN(
        n7281) );
  OAI22_X1 U47993 ( .A1(n68025), .A2(n62238), .B1(n68211), .B2(n68017), .ZN(
        n7282) );
  OAI22_X1 U47994 ( .A1(n68025), .A2(n62237), .B1(n68214), .B2(n68017), .ZN(
        n7283) );
  OAI22_X1 U47995 ( .A1(n68025), .A2(n62236), .B1(n68217), .B2(n68017), .ZN(
        n7284) );
  OAI22_X1 U47996 ( .A1(n68025), .A2(n62235), .B1(n68220), .B2(n68017), .ZN(
        n7285) );
  OAI22_X1 U47997 ( .A1(n68025), .A2(n62234), .B1(n68223), .B2(n68017), .ZN(
        n7286) );
  OAI22_X1 U47998 ( .A1(n68025), .A2(n62233), .B1(n68226), .B2(n68017), .ZN(
        n7287) );
  OAI22_X1 U47999 ( .A1(n68025), .A2(n62232), .B1(n68229), .B2(n68017), .ZN(
        n7288) );
  OAI22_X1 U48000 ( .A1(n68025), .A2(n62231), .B1(n68232), .B2(n68017), .ZN(
        n7289) );
  OAI22_X1 U48001 ( .A1(n68025), .A2(n62230), .B1(n68235), .B2(n68017), .ZN(
        n7290) );
  OAI22_X1 U48002 ( .A1(n67995), .A2(n62422), .B1(n68058), .B2(n67987), .ZN(
        n7103) );
  OAI22_X1 U48003 ( .A1(n67995), .A2(n62421), .B1(n68061), .B2(n67987), .ZN(
        n7104) );
  OAI22_X1 U48004 ( .A1(n67995), .A2(n62420), .B1(n68064), .B2(n67987), .ZN(
        n7105) );
  OAI22_X1 U48005 ( .A1(n67995), .A2(n62419), .B1(n68067), .B2(n67987), .ZN(
        n7106) );
  OAI22_X1 U48006 ( .A1(n67995), .A2(n62418), .B1(n68070), .B2(n67987), .ZN(
        n7107) );
  OAI22_X1 U48007 ( .A1(n67995), .A2(n62417), .B1(n68073), .B2(n67987), .ZN(
        n7108) );
  OAI22_X1 U48008 ( .A1(n67995), .A2(n62416), .B1(n68076), .B2(n67987), .ZN(
        n7109) );
  OAI22_X1 U48009 ( .A1(n67995), .A2(n62415), .B1(n68079), .B2(n67987), .ZN(
        n7110) );
  OAI22_X1 U48010 ( .A1(n67995), .A2(n62414), .B1(n68082), .B2(n67987), .ZN(
        n7111) );
  OAI22_X1 U48011 ( .A1(n67995), .A2(n62413), .B1(n68085), .B2(n67987), .ZN(
        n7112) );
  OAI22_X1 U48012 ( .A1(n67995), .A2(n62412), .B1(n68088), .B2(n67987), .ZN(
        n7113) );
  OAI22_X1 U48013 ( .A1(n67995), .A2(n62411), .B1(n68091), .B2(n67987), .ZN(
        n7114) );
  OAI22_X1 U48014 ( .A1(n67996), .A2(n62410), .B1(n68094), .B2(n67988), .ZN(
        n7115) );
  OAI22_X1 U48015 ( .A1(n67996), .A2(n62409), .B1(n68097), .B2(n67988), .ZN(
        n7116) );
  OAI22_X1 U48016 ( .A1(n67996), .A2(n62408), .B1(n68100), .B2(n67988), .ZN(
        n7117) );
  OAI22_X1 U48017 ( .A1(n67996), .A2(n62407), .B1(n68103), .B2(n67988), .ZN(
        n7118) );
  OAI22_X1 U48018 ( .A1(n67996), .A2(n62406), .B1(n68106), .B2(n67988), .ZN(
        n7119) );
  OAI22_X1 U48019 ( .A1(n67996), .A2(n62405), .B1(n68109), .B2(n67988), .ZN(
        n7120) );
  OAI22_X1 U48020 ( .A1(n67996), .A2(n62404), .B1(n68112), .B2(n67988), .ZN(
        n7121) );
  OAI22_X1 U48021 ( .A1(n67996), .A2(n62403), .B1(n68115), .B2(n67988), .ZN(
        n7122) );
  OAI22_X1 U48022 ( .A1(n67996), .A2(n62402), .B1(n68118), .B2(n67988), .ZN(
        n7123) );
  OAI22_X1 U48023 ( .A1(n67996), .A2(n62401), .B1(n68121), .B2(n67988), .ZN(
        n7124) );
  OAI22_X1 U48024 ( .A1(n67996), .A2(n62400), .B1(n68124), .B2(n67988), .ZN(
        n7125) );
  OAI22_X1 U48025 ( .A1(n67996), .A2(n62399), .B1(n68127), .B2(n67988), .ZN(
        n7126) );
  OAI22_X1 U48026 ( .A1(n67996), .A2(n62398), .B1(n68130), .B2(n67989), .ZN(
        n7127) );
  OAI22_X1 U48027 ( .A1(n67997), .A2(n62397), .B1(n68133), .B2(n67989), .ZN(
        n7128) );
  OAI22_X1 U48028 ( .A1(n67997), .A2(n62396), .B1(n68136), .B2(n67989), .ZN(
        n7129) );
  OAI22_X1 U48029 ( .A1(n67997), .A2(n62395), .B1(n68139), .B2(n67989), .ZN(
        n7130) );
  OAI22_X1 U48030 ( .A1(n67997), .A2(n62394), .B1(n68142), .B2(n67989), .ZN(
        n7131) );
  OAI22_X1 U48031 ( .A1(n67997), .A2(n62393), .B1(n68145), .B2(n67989), .ZN(
        n7132) );
  OAI22_X1 U48032 ( .A1(n67997), .A2(n62392), .B1(n68148), .B2(n67989), .ZN(
        n7133) );
  OAI22_X1 U48033 ( .A1(n67997), .A2(n62391), .B1(n68151), .B2(n67989), .ZN(
        n7134) );
  OAI22_X1 U48034 ( .A1(n67997), .A2(n62390), .B1(n68154), .B2(n67989), .ZN(
        n7135) );
  OAI22_X1 U48035 ( .A1(n67997), .A2(n62389), .B1(n68157), .B2(n67989), .ZN(
        n7136) );
  OAI22_X1 U48036 ( .A1(n67997), .A2(n62388), .B1(n68160), .B2(n67989), .ZN(
        n7137) );
  OAI22_X1 U48037 ( .A1(n67997), .A2(n62387), .B1(n68163), .B2(n67989), .ZN(
        n7138) );
  OAI22_X1 U48038 ( .A1(n67997), .A2(n62386), .B1(n68166), .B2(n67990), .ZN(
        n7139) );
  OAI22_X1 U48039 ( .A1(n67997), .A2(n62385), .B1(n68169), .B2(n67990), .ZN(
        n7140) );
  OAI22_X1 U48040 ( .A1(n67998), .A2(n62384), .B1(n68172), .B2(n67990), .ZN(
        n7141) );
  OAI22_X1 U48041 ( .A1(n67998), .A2(n62383), .B1(n68175), .B2(n67990), .ZN(
        n7142) );
  OAI22_X1 U48042 ( .A1(n67998), .A2(n62382), .B1(n68178), .B2(n67990), .ZN(
        n7143) );
  OAI22_X1 U48043 ( .A1(n67998), .A2(n62381), .B1(n68181), .B2(n67990), .ZN(
        n7144) );
  OAI22_X1 U48044 ( .A1(n67998), .A2(n62380), .B1(n68184), .B2(n67990), .ZN(
        n7145) );
  OAI22_X1 U48045 ( .A1(n67998), .A2(n62379), .B1(n68187), .B2(n67990), .ZN(
        n7146) );
  OAI22_X1 U48046 ( .A1(n67998), .A2(n62378), .B1(n68190), .B2(n67990), .ZN(
        n7147) );
  OAI22_X1 U48047 ( .A1(n67998), .A2(n62377), .B1(n68193), .B2(n67990), .ZN(
        n7148) );
  OAI22_X1 U48048 ( .A1(n67998), .A2(n62376), .B1(n68196), .B2(n67990), .ZN(
        n7149) );
  OAI22_X1 U48049 ( .A1(n67998), .A2(n62375), .B1(n68199), .B2(n67990), .ZN(
        n7150) );
  OAI22_X1 U48050 ( .A1(n67998), .A2(n62374), .B1(n68202), .B2(n67991), .ZN(
        n7151) );
  OAI22_X1 U48051 ( .A1(n67998), .A2(n62373), .B1(n68205), .B2(n67991), .ZN(
        n7152) );
  OAI22_X1 U48052 ( .A1(n67998), .A2(n62372), .B1(n68208), .B2(n67991), .ZN(
        n7153) );
  OAI22_X1 U48053 ( .A1(n67999), .A2(n62371), .B1(n68211), .B2(n67991), .ZN(
        n7154) );
  OAI22_X1 U48054 ( .A1(n67999), .A2(n62370), .B1(n68214), .B2(n67991), .ZN(
        n7155) );
  OAI22_X1 U48055 ( .A1(n67999), .A2(n62369), .B1(n68217), .B2(n67991), .ZN(
        n7156) );
  OAI22_X1 U48056 ( .A1(n67999), .A2(n62368), .B1(n68220), .B2(n67991), .ZN(
        n7157) );
  OAI22_X1 U48057 ( .A1(n67999), .A2(n62367), .B1(n68223), .B2(n67991), .ZN(
        n7158) );
  OAI22_X1 U48058 ( .A1(n67999), .A2(n62366), .B1(n68226), .B2(n67991), .ZN(
        n7159) );
  OAI22_X1 U48059 ( .A1(n67999), .A2(n62365), .B1(n68229), .B2(n67991), .ZN(
        n7160) );
  OAI22_X1 U48060 ( .A1(n67999), .A2(n62364), .B1(n68232), .B2(n67991), .ZN(
        n7161) );
  OAI22_X1 U48061 ( .A1(n67999), .A2(n62363), .B1(n68235), .B2(n67991), .ZN(
        n7162) );
  OAI22_X1 U48062 ( .A1(n67816), .A2(n63160), .B1(n68059), .B2(n67808), .ZN(
        n6207) );
  OAI22_X1 U48063 ( .A1(n67816), .A2(n63159), .B1(n68062), .B2(n67808), .ZN(
        n6208) );
  OAI22_X1 U48064 ( .A1(n67816), .A2(n63158), .B1(n68065), .B2(n67808), .ZN(
        n6209) );
  OAI22_X1 U48065 ( .A1(n67816), .A2(n63157), .B1(n68068), .B2(n67808), .ZN(
        n6210) );
  OAI22_X1 U48066 ( .A1(n67816), .A2(n63156), .B1(n68071), .B2(n67808), .ZN(
        n6211) );
  OAI22_X1 U48067 ( .A1(n67816), .A2(n63155), .B1(n68074), .B2(n67808), .ZN(
        n6212) );
  OAI22_X1 U48068 ( .A1(n67816), .A2(n63154), .B1(n68077), .B2(n67808), .ZN(
        n6213) );
  OAI22_X1 U48069 ( .A1(n67816), .A2(n63153), .B1(n68080), .B2(n67808), .ZN(
        n6214) );
  OAI22_X1 U48070 ( .A1(n67816), .A2(n63152), .B1(n68083), .B2(n67808), .ZN(
        n6215) );
  OAI22_X1 U48071 ( .A1(n67816), .A2(n63151), .B1(n68086), .B2(n67808), .ZN(
        n6216) );
  OAI22_X1 U48072 ( .A1(n67816), .A2(n63150), .B1(n68089), .B2(n67808), .ZN(
        n6217) );
  OAI22_X1 U48073 ( .A1(n67816), .A2(n63149), .B1(n68092), .B2(n67808), .ZN(
        n6218) );
  OAI22_X1 U48074 ( .A1(n67817), .A2(n63148), .B1(n68095), .B2(n67809), .ZN(
        n6219) );
  OAI22_X1 U48075 ( .A1(n67817), .A2(n63147), .B1(n68098), .B2(n67809), .ZN(
        n6220) );
  OAI22_X1 U48076 ( .A1(n67817), .A2(n63146), .B1(n68101), .B2(n67809), .ZN(
        n6221) );
  OAI22_X1 U48077 ( .A1(n67817), .A2(n63145), .B1(n68104), .B2(n67809), .ZN(
        n6222) );
  OAI22_X1 U48078 ( .A1(n67817), .A2(n63144), .B1(n68107), .B2(n67809), .ZN(
        n6223) );
  OAI22_X1 U48079 ( .A1(n67817), .A2(n63143), .B1(n68110), .B2(n67809), .ZN(
        n6224) );
  OAI22_X1 U48080 ( .A1(n67817), .A2(n63142), .B1(n68113), .B2(n67809), .ZN(
        n6225) );
  OAI22_X1 U48081 ( .A1(n67817), .A2(n63141), .B1(n68116), .B2(n67809), .ZN(
        n6226) );
  OAI22_X1 U48082 ( .A1(n67817), .A2(n63140), .B1(n68119), .B2(n67809), .ZN(
        n6227) );
  OAI22_X1 U48083 ( .A1(n67817), .A2(n63139), .B1(n68122), .B2(n67809), .ZN(
        n6228) );
  OAI22_X1 U48084 ( .A1(n67817), .A2(n63138), .B1(n68125), .B2(n67809), .ZN(
        n6229) );
  OAI22_X1 U48085 ( .A1(n67817), .A2(n63137), .B1(n68128), .B2(n67809), .ZN(
        n6230) );
  OAI22_X1 U48086 ( .A1(n67817), .A2(n63136), .B1(n68131), .B2(n67810), .ZN(
        n6231) );
  OAI22_X1 U48087 ( .A1(n67818), .A2(n63135), .B1(n68134), .B2(n67810), .ZN(
        n6232) );
  OAI22_X1 U48088 ( .A1(n67818), .A2(n63134), .B1(n68137), .B2(n67810), .ZN(
        n6233) );
  OAI22_X1 U48089 ( .A1(n67818), .A2(n63133), .B1(n68140), .B2(n67810), .ZN(
        n6234) );
  OAI22_X1 U48090 ( .A1(n67818), .A2(n63132), .B1(n68143), .B2(n67810), .ZN(
        n6235) );
  OAI22_X1 U48091 ( .A1(n67818), .A2(n63131), .B1(n68146), .B2(n67810), .ZN(
        n6236) );
  OAI22_X1 U48092 ( .A1(n67818), .A2(n63130), .B1(n68149), .B2(n67810), .ZN(
        n6237) );
  OAI22_X1 U48093 ( .A1(n67818), .A2(n63129), .B1(n68152), .B2(n67810), .ZN(
        n6238) );
  OAI22_X1 U48094 ( .A1(n67818), .A2(n63128), .B1(n68155), .B2(n67810), .ZN(
        n6239) );
  OAI22_X1 U48095 ( .A1(n67818), .A2(n63127), .B1(n68158), .B2(n67810), .ZN(
        n6240) );
  OAI22_X1 U48096 ( .A1(n67818), .A2(n63126), .B1(n68161), .B2(n67810), .ZN(
        n6241) );
  OAI22_X1 U48097 ( .A1(n67818), .A2(n63125), .B1(n68164), .B2(n67810), .ZN(
        n6242) );
  OAI22_X1 U48098 ( .A1(n67818), .A2(n63124), .B1(n68167), .B2(n67811), .ZN(
        n6243) );
  OAI22_X1 U48099 ( .A1(n67818), .A2(n63123), .B1(n68170), .B2(n67811), .ZN(
        n6244) );
  OAI22_X1 U48100 ( .A1(n67819), .A2(n63122), .B1(n68173), .B2(n67811), .ZN(
        n6245) );
  OAI22_X1 U48101 ( .A1(n67819), .A2(n63121), .B1(n68176), .B2(n67811), .ZN(
        n6246) );
  OAI22_X1 U48102 ( .A1(n67819), .A2(n63120), .B1(n68179), .B2(n67811), .ZN(
        n6247) );
  OAI22_X1 U48103 ( .A1(n67819), .A2(n63119), .B1(n68182), .B2(n67811), .ZN(
        n6248) );
  OAI22_X1 U48104 ( .A1(n67819), .A2(n63118), .B1(n68185), .B2(n67811), .ZN(
        n6249) );
  OAI22_X1 U48105 ( .A1(n67819), .A2(n63117), .B1(n68188), .B2(n67811), .ZN(
        n6250) );
  OAI22_X1 U48106 ( .A1(n67819), .A2(n63116), .B1(n68191), .B2(n67811), .ZN(
        n6251) );
  OAI22_X1 U48107 ( .A1(n67819), .A2(n63115), .B1(n68194), .B2(n67811), .ZN(
        n6252) );
  OAI22_X1 U48108 ( .A1(n67819), .A2(n63114), .B1(n68197), .B2(n67811), .ZN(
        n6253) );
  OAI22_X1 U48109 ( .A1(n67819), .A2(n63113), .B1(n68200), .B2(n67811), .ZN(
        n6254) );
  OAI22_X1 U48110 ( .A1(n67819), .A2(n63112), .B1(n68203), .B2(n67812), .ZN(
        n6255) );
  OAI22_X1 U48111 ( .A1(n67819), .A2(n63111), .B1(n68206), .B2(n67812), .ZN(
        n6256) );
  OAI22_X1 U48112 ( .A1(n67819), .A2(n63110), .B1(n68209), .B2(n67812), .ZN(
        n6257) );
  OAI22_X1 U48113 ( .A1(n67820), .A2(n63109), .B1(n68212), .B2(n67812), .ZN(
        n6258) );
  OAI22_X1 U48114 ( .A1(n67820), .A2(n63108), .B1(n68215), .B2(n67812), .ZN(
        n6259) );
  OAI22_X1 U48115 ( .A1(n67820), .A2(n63107), .B1(n68218), .B2(n67812), .ZN(
        n6260) );
  OAI22_X1 U48116 ( .A1(n67820), .A2(n63106), .B1(n68221), .B2(n67812), .ZN(
        n6261) );
  OAI22_X1 U48117 ( .A1(n67820), .A2(n63105), .B1(n68224), .B2(n67812), .ZN(
        n6262) );
  OAI22_X1 U48118 ( .A1(n67820), .A2(n63104), .B1(n68227), .B2(n67812), .ZN(
        n6263) );
  OAI22_X1 U48119 ( .A1(n67820), .A2(n63103), .B1(n68230), .B2(n67812), .ZN(
        n6264) );
  OAI22_X1 U48120 ( .A1(n67820), .A2(n63102), .B1(n68233), .B2(n67812), .ZN(
        n6265) );
  OAI22_X1 U48121 ( .A1(n67820), .A2(n63101), .B1(n68236), .B2(n67812), .ZN(
        n6266) );
  OAI22_X1 U48122 ( .A1(n67982), .A2(n62488), .B1(n68058), .B2(n67974), .ZN(
        n7039) );
  OAI22_X1 U48123 ( .A1(n67982), .A2(n62487), .B1(n68061), .B2(n67974), .ZN(
        n7040) );
  OAI22_X1 U48124 ( .A1(n67982), .A2(n62486), .B1(n68064), .B2(n67974), .ZN(
        n7041) );
  OAI22_X1 U48125 ( .A1(n67982), .A2(n62485), .B1(n68067), .B2(n67974), .ZN(
        n7042) );
  OAI22_X1 U48126 ( .A1(n67982), .A2(n62484), .B1(n68070), .B2(n67974), .ZN(
        n7043) );
  OAI22_X1 U48127 ( .A1(n67982), .A2(n62483), .B1(n68073), .B2(n67974), .ZN(
        n7044) );
  OAI22_X1 U48128 ( .A1(n67982), .A2(n62482), .B1(n68076), .B2(n67974), .ZN(
        n7045) );
  OAI22_X1 U48129 ( .A1(n67982), .A2(n62481), .B1(n68079), .B2(n67974), .ZN(
        n7046) );
  OAI22_X1 U48130 ( .A1(n67982), .A2(n62480), .B1(n68082), .B2(n67974), .ZN(
        n7047) );
  OAI22_X1 U48131 ( .A1(n67982), .A2(n62479), .B1(n68085), .B2(n67974), .ZN(
        n7048) );
  OAI22_X1 U48132 ( .A1(n67982), .A2(n62478), .B1(n68088), .B2(n67974), .ZN(
        n7049) );
  OAI22_X1 U48133 ( .A1(n67982), .A2(n62477), .B1(n68091), .B2(n67974), .ZN(
        n7050) );
  OAI22_X1 U48134 ( .A1(n67983), .A2(n62476), .B1(n68094), .B2(n67975), .ZN(
        n7051) );
  OAI22_X1 U48135 ( .A1(n67983), .A2(n62475), .B1(n68097), .B2(n67975), .ZN(
        n7052) );
  OAI22_X1 U48136 ( .A1(n67983), .A2(n62474), .B1(n68100), .B2(n67975), .ZN(
        n7053) );
  OAI22_X1 U48137 ( .A1(n67983), .A2(n62473), .B1(n68103), .B2(n67975), .ZN(
        n7054) );
  OAI22_X1 U48138 ( .A1(n67983), .A2(n62472), .B1(n68106), .B2(n67975), .ZN(
        n7055) );
  OAI22_X1 U48139 ( .A1(n67983), .A2(n62471), .B1(n68109), .B2(n67975), .ZN(
        n7056) );
  OAI22_X1 U48140 ( .A1(n67983), .A2(n62470), .B1(n68112), .B2(n67975), .ZN(
        n7057) );
  OAI22_X1 U48141 ( .A1(n67983), .A2(n62469), .B1(n68115), .B2(n67975), .ZN(
        n7058) );
  OAI22_X1 U48142 ( .A1(n67983), .A2(n62468), .B1(n68118), .B2(n67975), .ZN(
        n7059) );
  OAI22_X1 U48143 ( .A1(n67983), .A2(n62467), .B1(n68121), .B2(n67975), .ZN(
        n7060) );
  OAI22_X1 U48144 ( .A1(n67983), .A2(n62466), .B1(n68124), .B2(n67975), .ZN(
        n7061) );
  OAI22_X1 U48145 ( .A1(n67983), .A2(n62465), .B1(n68127), .B2(n67975), .ZN(
        n7062) );
  OAI22_X1 U48146 ( .A1(n67983), .A2(n62464), .B1(n68130), .B2(n67976), .ZN(
        n7063) );
  OAI22_X1 U48147 ( .A1(n67984), .A2(n62463), .B1(n68133), .B2(n67976), .ZN(
        n7064) );
  OAI22_X1 U48148 ( .A1(n67984), .A2(n62462), .B1(n68136), .B2(n67976), .ZN(
        n7065) );
  OAI22_X1 U48149 ( .A1(n67984), .A2(n62461), .B1(n68139), .B2(n67976), .ZN(
        n7066) );
  OAI22_X1 U48150 ( .A1(n67984), .A2(n62460), .B1(n68142), .B2(n67976), .ZN(
        n7067) );
  OAI22_X1 U48151 ( .A1(n67984), .A2(n62459), .B1(n68145), .B2(n67976), .ZN(
        n7068) );
  OAI22_X1 U48152 ( .A1(n67984), .A2(n62458), .B1(n68148), .B2(n67976), .ZN(
        n7069) );
  OAI22_X1 U48153 ( .A1(n67984), .A2(n62457), .B1(n68151), .B2(n67976), .ZN(
        n7070) );
  OAI22_X1 U48154 ( .A1(n67984), .A2(n62456), .B1(n68154), .B2(n67976), .ZN(
        n7071) );
  OAI22_X1 U48155 ( .A1(n67984), .A2(n62455), .B1(n68157), .B2(n67976), .ZN(
        n7072) );
  OAI22_X1 U48156 ( .A1(n67984), .A2(n62454), .B1(n68160), .B2(n67976), .ZN(
        n7073) );
  OAI22_X1 U48157 ( .A1(n67984), .A2(n62453), .B1(n68163), .B2(n67976), .ZN(
        n7074) );
  OAI22_X1 U48158 ( .A1(n67984), .A2(n62452), .B1(n68166), .B2(n67977), .ZN(
        n7075) );
  OAI22_X1 U48159 ( .A1(n67984), .A2(n62451), .B1(n68169), .B2(n67977), .ZN(
        n7076) );
  OAI22_X1 U48160 ( .A1(n67985), .A2(n62450), .B1(n68172), .B2(n67977), .ZN(
        n7077) );
  OAI22_X1 U48161 ( .A1(n67985), .A2(n62449), .B1(n68175), .B2(n67977), .ZN(
        n7078) );
  OAI22_X1 U48162 ( .A1(n67985), .A2(n62448), .B1(n68178), .B2(n67977), .ZN(
        n7079) );
  OAI22_X1 U48163 ( .A1(n67985), .A2(n62447), .B1(n68181), .B2(n67977), .ZN(
        n7080) );
  OAI22_X1 U48164 ( .A1(n67985), .A2(n62446), .B1(n68184), .B2(n67977), .ZN(
        n7081) );
  OAI22_X1 U48165 ( .A1(n67985), .A2(n62445), .B1(n68187), .B2(n67977), .ZN(
        n7082) );
  OAI22_X1 U48166 ( .A1(n67985), .A2(n62444), .B1(n68190), .B2(n67977), .ZN(
        n7083) );
  OAI22_X1 U48167 ( .A1(n67985), .A2(n62443), .B1(n68193), .B2(n67977), .ZN(
        n7084) );
  OAI22_X1 U48168 ( .A1(n67985), .A2(n62442), .B1(n68196), .B2(n67977), .ZN(
        n7085) );
  OAI22_X1 U48169 ( .A1(n67985), .A2(n62441), .B1(n68199), .B2(n67977), .ZN(
        n7086) );
  OAI22_X1 U48170 ( .A1(n67985), .A2(n62440), .B1(n68202), .B2(n67978), .ZN(
        n7087) );
  OAI22_X1 U48171 ( .A1(n67985), .A2(n62439), .B1(n68205), .B2(n67978), .ZN(
        n7088) );
  OAI22_X1 U48172 ( .A1(n67985), .A2(n62438), .B1(n68208), .B2(n67978), .ZN(
        n7089) );
  OAI22_X1 U48173 ( .A1(n67986), .A2(n62437), .B1(n68211), .B2(n67978), .ZN(
        n7090) );
  OAI22_X1 U48174 ( .A1(n67986), .A2(n62436), .B1(n68214), .B2(n67978), .ZN(
        n7091) );
  OAI22_X1 U48175 ( .A1(n67986), .A2(n62435), .B1(n68217), .B2(n67978), .ZN(
        n7092) );
  OAI22_X1 U48176 ( .A1(n67986), .A2(n62434), .B1(n68220), .B2(n67978), .ZN(
        n7093) );
  OAI22_X1 U48177 ( .A1(n67986), .A2(n62433), .B1(n68223), .B2(n67978), .ZN(
        n7094) );
  OAI22_X1 U48178 ( .A1(n67986), .A2(n62432), .B1(n68226), .B2(n67978), .ZN(
        n7095) );
  OAI22_X1 U48179 ( .A1(n67986), .A2(n62431), .B1(n68229), .B2(n67978), .ZN(
        n7096) );
  OAI22_X1 U48180 ( .A1(n67986), .A2(n62430), .B1(n68232), .B2(n67978), .ZN(
        n7097) );
  OAI22_X1 U48181 ( .A1(n67986), .A2(n62429), .B1(n68235), .B2(n67978), .ZN(
        n7098) );
  OAI22_X1 U48182 ( .A1(n67765), .A2(n63361), .B1(n68059), .B2(n67757), .ZN(
        n5951) );
  OAI22_X1 U48183 ( .A1(n67765), .A2(n63360), .B1(n68062), .B2(n67757), .ZN(
        n5952) );
  OAI22_X1 U48184 ( .A1(n67765), .A2(n63359), .B1(n68065), .B2(n67757), .ZN(
        n5953) );
  OAI22_X1 U48185 ( .A1(n67765), .A2(n63358), .B1(n68068), .B2(n67757), .ZN(
        n5954) );
  OAI22_X1 U48186 ( .A1(n67765), .A2(n63357), .B1(n68071), .B2(n67757), .ZN(
        n5955) );
  OAI22_X1 U48187 ( .A1(n67765), .A2(n63356), .B1(n68074), .B2(n67757), .ZN(
        n5956) );
  OAI22_X1 U48188 ( .A1(n67765), .A2(n63355), .B1(n68077), .B2(n67757), .ZN(
        n5957) );
  OAI22_X1 U48189 ( .A1(n67765), .A2(n63354), .B1(n68080), .B2(n67757), .ZN(
        n5958) );
  OAI22_X1 U48190 ( .A1(n67765), .A2(n63353), .B1(n68083), .B2(n67757), .ZN(
        n5959) );
  OAI22_X1 U48191 ( .A1(n67765), .A2(n63352), .B1(n68086), .B2(n67757), .ZN(
        n5960) );
  OAI22_X1 U48192 ( .A1(n67765), .A2(n63351), .B1(n68089), .B2(n67757), .ZN(
        n5961) );
  OAI22_X1 U48193 ( .A1(n67765), .A2(n63350), .B1(n68092), .B2(n67757), .ZN(
        n5962) );
  OAI22_X1 U48194 ( .A1(n67766), .A2(n63349), .B1(n68095), .B2(n67758), .ZN(
        n5963) );
  OAI22_X1 U48195 ( .A1(n67766), .A2(n63348), .B1(n68098), .B2(n67758), .ZN(
        n5964) );
  OAI22_X1 U48196 ( .A1(n67766), .A2(n63347), .B1(n68101), .B2(n67758), .ZN(
        n5965) );
  OAI22_X1 U48197 ( .A1(n67766), .A2(n63346), .B1(n68104), .B2(n67758), .ZN(
        n5966) );
  OAI22_X1 U48198 ( .A1(n67766), .A2(n63345), .B1(n68107), .B2(n67758), .ZN(
        n5967) );
  OAI22_X1 U48199 ( .A1(n67766), .A2(n63344), .B1(n68110), .B2(n67758), .ZN(
        n5968) );
  OAI22_X1 U48200 ( .A1(n67766), .A2(n63343), .B1(n68113), .B2(n67758), .ZN(
        n5969) );
  OAI22_X1 U48201 ( .A1(n67766), .A2(n63342), .B1(n68116), .B2(n67758), .ZN(
        n5970) );
  OAI22_X1 U48202 ( .A1(n67766), .A2(n63341), .B1(n68119), .B2(n67758), .ZN(
        n5971) );
  OAI22_X1 U48203 ( .A1(n67766), .A2(n63340), .B1(n68122), .B2(n67758), .ZN(
        n5972) );
  OAI22_X1 U48204 ( .A1(n67766), .A2(n63339), .B1(n68125), .B2(n67758), .ZN(
        n5973) );
  OAI22_X1 U48205 ( .A1(n67766), .A2(n63338), .B1(n68128), .B2(n67758), .ZN(
        n5974) );
  OAI22_X1 U48206 ( .A1(n67766), .A2(n63337), .B1(n68131), .B2(n67759), .ZN(
        n5975) );
  OAI22_X1 U48207 ( .A1(n67767), .A2(n63336), .B1(n68134), .B2(n67759), .ZN(
        n5976) );
  OAI22_X1 U48208 ( .A1(n67767), .A2(n63335), .B1(n68137), .B2(n67759), .ZN(
        n5977) );
  OAI22_X1 U48209 ( .A1(n67767), .A2(n63334), .B1(n68140), .B2(n67759), .ZN(
        n5978) );
  OAI22_X1 U48210 ( .A1(n67767), .A2(n63333), .B1(n68143), .B2(n67759), .ZN(
        n5979) );
  OAI22_X1 U48211 ( .A1(n67767), .A2(n63332), .B1(n68146), .B2(n67759), .ZN(
        n5980) );
  OAI22_X1 U48212 ( .A1(n67767), .A2(n63331), .B1(n68149), .B2(n67759), .ZN(
        n5981) );
  OAI22_X1 U48213 ( .A1(n67767), .A2(n63330), .B1(n68152), .B2(n67759), .ZN(
        n5982) );
  OAI22_X1 U48214 ( .A1(n67767), .A2(n63329), .B1(n68155), .B2(n67759), .ZN(
        n5983) );
  OAI22_X1 U48215 ( .A1(n67767), .A2(n63328), .B1(n68158), .B2(n67759), .ZN(
        n5984) );
  OAI22_X1 U48216 ( .A1(n67767), .A2(n63327), .B1(n68161), .B2(n67759), .ZN(
        n5985) );
  OAI22_X1 U48217 ( .A1(n67767), .A2(n63326), .B1(n68164), .B2(n67759), .ZN(
        n5986) );
  OAI22_X1 U48218 ( .A1(n67767), .A2(n63325), .B1(n68167), .B2(n67760), .ZN(
        n5987) );
  OAI22_X1 U48219 ( .A1(n67767), .A2(n63324), .B1(n68170), .B2(n67760), .ZN(
        n5988) );
  OAI22_X1 U48220 ( .A1(n67768), .A2(n63323), .B1(n68173), .B2(n67760), .ZN(
        n5989) );
  OAI22_X1 U48221 ( .A1(n67768), .A2(n63322), .B1(n68176), .B2(n67760), .ZN(
        n5990) );
  OAI22_X1 U48222 ( .A1(n67768), .A2(n63321), .B1(n68179), .B2(n67760), .ZN(
        n5991) );
  OAI22_X1 U48223 ( .A1(n67768), .A2(n63320), .B1(n68182), .B2(n67760), .ZN(
        n5992) );
  OAI22_X1 U48224 ( .A1(n67768), .A2(n63319), .B1(n68185), .B2(n67760), .ZN(
        n5993) );
  OAI22_X1 U48225 ( .A1(n67768), .A2(n63318), .B1(n68188), .B2(n67760), .ZN(
        n5994) );
  OAI22_X1 U48226 ( .A1(n67768), .A2(n63317), .B1(n68191), .B2(n67760), .ZN(
        n5995) );
  OAI22_X1 U48227 ( .A1(n67768), .A2(n63316), .B1(n68194), .B2(n67760), .ZN(
        n5996) );
  OAI22_X1 U48228 ( .A1(n67768), .A2(n63315), .B1(n68197), .B2(n67760), .ZN(
        n5997) );
  OAI22_X1 U48229 ( .A1(n67768), .A2(n63314), .B1(n68200), .B2(n67760), .ZN(
        n5998) );
  OAI22_X1 U48230 ( .A1(n67768), .A2(n63313), .B1(n68203), .B2(n67761), .ZN(
        n5999) );
  OAI22_X1 U48231 ( .A1(n67768), .A2(n63312), .B1(n68206), .B2(n67761), .ZN(
        n6000) );
  OAI22_X1 U48232 ( .A1(n67768), .A2(n63311), .B1(n68209), .B2(n67761), .ZN(
        n6001) );
  OAI22_X1 U48233 ( .A1(n67769), .A2(n63310), .B1(n68212), .B2(n67761), .ZN(
        n6002) );
  OAI22_X1 U48234 ( .A1(n67769), .A2(n63309), .B1(n68215), .B2(n67761), .ZN(
        n6003) );
  OAI22_X1 U48235 ( .A1(n67769), .A2(n63308), .B1(n68218), .B2(n67761), .ZN(
        n6004) );
  OAI22_X1 U48236 ( .A1(n67769), .A2(n63307), .B1(n68221), .B2(n67761), .ZN(
        n6005) );
  OAI22_X1 U48237 ( .A1(n67769), .A2(n63306), .B1(n68224), .B2(n67761), .ZN(
        n6006) );
  OAI22_X1 U48238 ( .A1(n67769), .A2(n63305), .B1(n68227), .B2(n67761), .ZN(
        n6007) );
  OAI22_X1 U48239 ( .A1(n67769), .A2(n63304), .B1(n68230), .B2(n67761), .ZN(
        n6008) );
  OAI22_X1 U48240 ( .A1(n67769), .A2(n63303), .B1(n68233), .B2(n67761), .ZN(
        n6009) );
  OAI22_X1 U48241 ( .A1(n67769), .A2(n63302), .B1(n68236), .B2(n67761), .ZN(
        n6010) );
  OAI22_X1 U48242 ( .A1(n67867), .A2(n62957), .B1(n68059), .B2(n67859), .ZN(
        n6463) );
  OAI22_X1 U48243 ( .A1(n67867), .A2(n62956), .B1(n68062), .B2(n67859), .ZN(
        n6464) );
  OAI22_X1 U48244 ( .A1(n67867), .A2(n62955), .B1(n68065), .B2(n67859), .ZN(
        n6465) );
  OAI22_X1 U48245 ( .A1(n67867), .A2(n62954), .B1(n68068), .B2(n67859), .ZN(
        n6466) );
  OAI22_X1 U48246 ( .A1(n67867), .A2(n62953), .B1(n68071), .B2(n67859), .ZN(
        n6467) );
  OAI22_X1 U48247 ( .A1(n67867), .A2(n62952), .B1(n68074), .B2(n67859), .ZN(
        n6468) );
  OAI22_X1 U48248 ( .A1(n67867), .A2(n62951), .B1(n68077), .B2(n67859), .ZN(
        n6469) );
  OAI22_X1 U48249 ( .A1(n67867), .A2(n62950), .B1(n68080), .B2(n67859), .ZN(
        n6470) );
  OAI22_X1 U48250 ( .A1(n67867), .A2(n62949), .B1(n68083), .B2(n67859), .ZN(
        n6471) );
  OAI22_X1 U48251 ( .A1(n67867), .A2(n62948), .B1(n68086), .B2(n67859), .ZN(
        n6472) );
  OAI22_X1 U48252 ( .A1(n67867), .A2(n62947), .B1(n68089), .B2(n67859), .ZN(
        n6473) );
  OAI22_X1 U48253 ( .A1(n67867), .A2(n62946), .B1(n68092), .B2(n67859), .ZN(
        n6474) );
  OAI22_X1 U48254 ( .A1(n67868), .A2(n62945), .B1(n68095), .B2(n67860), .ZN(
        n6475) );
  OAI22_X1 U48255 ( .A1(n67868), .A2(n62944), .B1(n68098), .B2(n67860), .ZN(
        n6476) );
  OAI22_X1 U48256 ( .A1(n67868), .A2(n62943), .B1(n68101), .B2(n67860), .ZN(
        n6477) );
  OAI22_X1 U48257 ( .A1(n67868), .A2(n62942), .B1(n68104), .B2(n67860), .ZN(
        n6478) );
  OAI22_X1 U48258 ( .A1(n67868), .A2(n62941), .B1(n68107), .B2(n67860), .ZN(
        n6479) );
  OAI22_X1 U48259 ( .A1(n67868), .A2(n62940), .B1(n68110), .B2(n67860), .ZN(
        n6480) );
  OAI22_X1 U48260 ( .A1(n67868), .A2(n62939), .B1(n68113), .B2(n67860), .ZN(
        n6481) );
  OAI22_X1 U48261 ( .A1(n67868), .A2(n62938), .B1(n68116), .B2(n67860), .ZN(
        n6482) );
  OAI22_X1 U48262 ( .A1(n67868), .A2(n62937), .B1(n68119), .B2(n67860), .ZN(
        n6483) );
  OAI22_X1 U48263 ( .A1(n67868), .A2(n62936), .B1(n68122), .B2(n67860), .ZN(
        n6484) );
  OAI22_X1 U48264 ( .A1(n67868), .A2(n62935), .B1(n68125), .B2(n67860), .ZN(
        n6485) );
  OAI22_X1 U48265 ( .A1(n67868), .A2(n62934), .B1(n68128), .B2(n67860), .ZN(
        n6486) );
  OAI22_X1 U48266 ( .A1(n67868), .A2(n62933), .B1(n68131), .B2(n67861), .ZN(
        n6487) );
  OAI22_X1 U48267 ( .A1(n67869), .A2(n62932), .B1(n68134), .B2(n67861), .ZN(
        n6488) );
  OAI22_X1 U48268 ( .A1(n67869), .A2(n62931), .B1(n68137), .B2(n67861), .ZN(
        n6489) );
  OAI22_X1 U48269 ( .A1(n67869), .A2(n62930), .B1(n68140), .B2(n67861), .ZN(
        n6490) );
  OAI22_X1 U48270 ( .A1(n67869), .A2(n62929), .B1(n68143), .B2(n67861), .ZN(
        n6491) );
  OAI22_X1 U48271 ( .A1(n67869), .A2(n62928), .B1(n68146), .B2(n67861), .ZN(
        n6492) );
  OAI22_X1 U48272 ( .A1(n67869), .A2(n62927), .B1(n68149), .B2(n67861), .ZN(
        n6493) );
  OAI22_X1 U48273 ( .A1(n67869), .A2(n62926), .B1(n68152), .B2(n67861), .ZN(
        n6494) );
  OAI22_X1 U48274 ( .A1(n67869), .A2(n62925), .B1(n68155), .B2(n67861), .ZN(
        n6495) );
  OAI22_X1 U48275 ( .A1(n67869), .A2(n62924), .B1(n68158), .B2(n67861), .ZN(
        n6496) );
  OAI22_X1 U48276 ( .A1(n67869), .A2(n62923), .B1(n68161), .B2(n67861), .ZN(
        n6497) );
  OAI22_X1 U48277 ( .A1(n67869), .A2(n62922), .B1(n68164), .B2(n67861), .ZN(
        n6498) );
  OAI22_X1 U48278 ( .A1(n67869), .A2(n62921), .B1(n68167), .B2(n67862), .ZN(
        n6499) );
  OAI22_X1 U48279 ( .A1(n67869), .A2(n62920), .B1(n68170), .B2(n67862), .ZN(
        n6500) );
  OAI22_X1 U48280 ( .A1(n67870), .A2(n62919), .B1(n68173), .B2(n67862), .ZN(
        n6501) );
  OAI22_X1 U48281 ( .A1(n67870), .A2(n62918), .B1(n68176), .B2(n67862), .ZN(
        n6502) );
  OAI22_X1 U48282 ( .A1(n67870), .A2(n62917), .B1(n68179), .B2(n67862), .ZN(
        n6503) );
  OAI22_X1 U48283 ( .A1(n67870), .A2(n62916), .B1(n68182), .B2(n67862), .ZN(
        n6504) );
  OAI22_X1 U48284 ( .A1(n67870), .A2(n62915), .B1(n68185), .B2(n67862), .ZN(
        n6505) );
  OAI22_X1 U48285 ( .A1(n67870), .A2(n62914), .B1(n68188), .B2(n67862), .ZN(
        n6506) );
  OAI22_X1 U48286 ( .A1(n67870), .A2(n62913), .B1(n68191), .B2(n67862), .ZN(
        n6507) );
  OAI22_X1 U48287 ( .A1(n67870), .A2(n62912), .B1(n68194), .B2(n67862), .ZN(
        n6508) );
  OAI22_X1 U48288 ( .A1(n67870), .A2(n62911), .B1(n68197), .B2(n67862), .ZN(
        n6509) );
  OAI22_X1 U48289 ( .A1(n67870), .A2(n62910), .B1(n68200), .B2(n67862), .ZN(
        n6510) );
  OAI22_X1 U48290 ( .A1(n67870), .A2(n62909), .B1(n68203), .B2(n67863), .ZN(
        n6511) );
  OAI22_X1 U48291 ( .A1(n67870), .A2(n62908), .B1(n68206), .B2(n67863), .ZN(
        n6512) );
  OAI22_X1 U48292 ( .A1(n67870), .A2(n62907), .B1(n68209), .B2(n67863), .ZN(
        n6513) );
  OAI22_X1 U48293 ( .A1(n67871), .A2(n62906), .B1(n68212), .B2(n67863), .ZN(
        n6514) );
  OAI22_X1 U48294 ( .A1(n67871), .A2(n62905), .B1(n68215), .B2(n67863), .ZN(
        n6515) );
  OAI22_X1 U48295 ( .A1(n67871), .A2(n62904), .B1(n68218), .B2(n67863), .ZN(
        n6516) );
  OAI22_X1 U48296 ( .A1(n67871), .A2(n62903), .B1(n68221), .B2(n67863), .ZN(
        n6517) );
  OAI22_X1 U48297 ( .A1(n67871), .A2(n62902), .B1(n68224), .B2(n67863), .ZN(
        n6518) );
  OAI22_X1 U48298 ( .A1(n67871), .A2(n62901), .B1(n68227), .B2(n67863), .ZN(
        n6519) );
  OAI22_X1 U48299 ( .A1(n67871), .A2(n62900), .B1(n68230), .B2(n67863), .ZN(
        n6520) );
  OAI22_X1 U48300 ( .A1(n67871), .A2(n62899), .B1(n68233), .B2(n67863), .ZN(
        n6521) );
  OAI22_X1 U48301 ( .A1(n67871), .A2(n62898), .B1(n68236), .B2(n67863), .ZN(
        n6522) );
  OAI22_X1 U48302 ( .A1(n67918), .A2(n62761), .B1(n68058), .B2(n67910), .ZN(
        n6719) );
  OAI22_X1 U48303 ( .A1(n67918), .A2(n62760), .B1(n68061), .B2(n67910), .ZN(
        n6720) );
  OAI22_X1 U48304 ( .A1(n67918), .A2(n62759), .B1(n68064), .B2(n67910), .ZN(
        n6721) );
  OAI22_X1 U48305 ( .A1(n67918), .A2(n62758), .B1(n68067), .B2(n67910), .ZN(
        n6722) );
  OAI22_X1 U48306 ( .A1(n67918), .A2(n62757), .B1(n68070), .B2(n67910), .ZN(
        n6723) );
  OAI22_X1 U48307 ( .A1(n67918), .A2(n62756), .B1(n68073), .B2(n67910), .ZN(
        n6724) );
  OAI22_X1 U48308 ( .A1(n67918), .A2(n62755), .B1(n68076), .B2(n67910), .ZN(
        n6725) );
  OAI22_X1 U48309 ( .A1(n67918), .A2(n62754), .B1(n68079), .B2(n67910), .ZN(
        n6726) );
  OAI22_X1 U48310 ( .A1(n67918), .A2(n62753), .B1(n68082), .B2(n67910), .ZN(
        n6727) );
  OAI22_X1 U48311 ( .A1(n67918), .A2(n62752), .B1(n68085), .B2(n67910), .ZN(
        n6728) );
  OAI22_X1 U48312 ( .A1(n67918), .A2(n62751), .B1(n68088), .B2(n67910), .ZN(
        n6729) );
  OAI22_X1 U48313 ( .A1(n67918), .A2(n62750), .B1(n68091), .B2(n67910), .ZN(
        n6730) );
  OAI22_X1 U48314 ( .A1(n67919), .A2(n62749), .B1(n68094), .B2(n67911), .ZN(
        n6731) );
  OAI22_X1 U48315 ( .A1(n67919), .A2(n62748), .B1(n68097), .B2(n67911), .ZN(
        n6732) );
  OAI22_X1 U48316 ( .A1(n67919), .A2(n62747), .B1(n68100), .B2(n67911), .ZN(
        n6733) );
  OAI22_X1 U48317 ( .A1(n67919), .A2(n62746), .B1(n68103), .B2(n67911), .ZN(
        n6734) );
  OAI22_X1 U48318 ( .A1(n67919), .A2(n62745), .B1(n68106), .B2(n67911), .ZN(
        n6735) );
  OAI22_X1 U48319 ( .A1(n67919), .A2(n62744), .B1(n68109), .B2(n67911), .ZN(
        n6736) );
  OAI22_X1 U48320 ( .A1(n67919), .A2(n62743), .B1(n68112), .B2(n67911), .ZN(
        n6737) );
  OAI22_X1 U48321 ( .A1(n67919), .A2(n62742), .B1(n68115), .B2(n67911), .ZN(
        n6738) );
  OAI22_X1 U48322 ( .A1(n67919), .A2(n62741), .B1(n68118), .B2(n67911), .ZN(
        n6739) );
  OAI22_X1 U48323 ( .A1(n67919), .A2(n62740), .B1(n68121), .B2(n67911), .ZN(
        n6740) );
  OAI22_X1 U48324 ( .A1(n67919), .A2(n62739), .B1(n68124), .B2(n67911), .ZN(
        n6741) );
  OAI22_X1 U48325 ( .A1(n67919), .A2(n62738), .B1(n68127), .B2(n67911), .ZN(
        n6742) );
  OAI22_X1 U48326 ( .A1(n67919), .A2(n62737), .B1(n68130), .B2(n67912), .ZN(
        n6743) );
  OAI22_X1 U48327 ( .A1(n67920), .A2(n62736), .B1(n68133), .B2(n67912), .ZN(
        n6744) );
  OAI22_X1 U48328 ( .A1(n67920), .A2(n62735), .B1(n68136), .B2(n67912), .ZN(
        n6745) );
  OAI22_X1 U48329 ( .A1(n67920), .A2(n62734), .B1(n68139), .B2(n67912), .ZN(
        n6746) );
  OAI22_X1 U48330 ( .A1(n67920), .A2(n62733), .B1(n68142), .B2(n67912), .ZN(
        n6747) );
  OAI22_X1 U48331 ( .A1(n67920), .A2(n62732), .B1(n68145), .B2(n67912), .ZN(
        n6748) );
  OAI22_X1 U48332 ( .A1(n67920), .A2(n62731), .B1(n68148), .B2(n67912), .ZN(
        n6749) );
  OAI22_X1 U48333 ( .A1(n67920), .A2(n62730), .B1(n68151), .B2(n67912), .ZN(
        n6750) );
  OAI22_X1 U48334 ( .A1(n67920), .A2(n62729), .B1(n68154), .B2(n67912), .ZN(
        n6751) );
  OAI22_X1 U48335 ( .A1(n67920), .A2(n62728), .B1(n68157), .B2(n67912), .ZN(
        n6752) );
  OAI22_X1 U48336 ( .A1(n67920), .A2(n62727), .B1(n68160), .B2(n67912), .ZN(
        n6753) );
  OAI22_X1 U48337 ( .A1(n67920), .A2(n62726), .B1(n68163), .B2(n67912), .ZN(
        n6754) );
  OAI22_X1 U48338 ( .A1(n67920), .A2(n62725), .B1(n68166), .B2(n67913), .ZN(
        n6755) );
  OAI22_X1 U48339 ( .A1(n67920), .A2(n62724), .B1(n68169), .B2(n67913), .ZN(
        n6756) );
  OAI22_X1 U48340 ( .A1(n67921), .A2(n62723), .B1(n68172), .B2(n67913), .ZN(
        n6757) );
  OAI22_X1 U48341 ( .A1(n67921), .A2(n62722), .B1(n68175), .B2(n67913), .ZN(
        n6758) );
  OAI22_X1 U48342 ( .A1(n67921), .A2(n62721), .B1(n68178), .B2(n67913), .ZN(
        n6759) );
  OAI22_X1 U48343 ( .A1(n67921), .A2(n62720), .B1(n68181), .B2(n67913), .ZN(
        n6760) );
  OAI22_X1 U48344 ( .A1(n67921), .A2(n62719), .B1(n68184), .B2(n67913), .ZN(
        n6761) );
  OAI22_X1 U48345 ( .A1(n67921), .A2(n62718), .B1(n68187), .B2(n67913), .ZN(
        n6762) );
  OAI22_X1 U48346 ( .A1(n67921), .A2(n62717), .B1(n68190), .B2(n67913), .ZN(
        n6763) );
  OAI22_X1 U48347 ( .A1(n67921), .A2(n62716), .B1(n68193), .B2(n67913), .ZN(
        n6764) );
  OAI22_X1 U48348 ( .A1(n67921), .A2(n62715), .B1(n68196), .B2(n67913), .ZN(
        n6765) );
  OAI22_X1 U48349 ( .A1(n67921), .A2(n62714), .B1(n68199), .B2(n67913), .ZN(
        n6766) );
  OAI22_X1 U48350 ( .A1(n67921), .A2(n62713), .B1(n68202), .B2(n67914), .ZN(
        n6767) );
  OAI22_X1 U48351 ( .A1(n67921), .A2(n62712), .B1(n68205), .B2(n67914), .ZN(
        n6768) );
  OAI22_X1 U48352 ( .A1(n67921), .A2(n62711), .B1(n68208), .B2(n67914), .ZN(
        n6769) );
  OAI22_X1 U48353 ( .A1(n67922), .A2(n62710), .B1(n68211), .B2(n67914), .ZN(
        n6770) );
  OAI22_X1 U48354 ( .A1(n67922), .A2(n62709), .B1(n68214), .B2(n67914), .ZN(
        n6771) );
  OAI22_X1 U48355 ( .A1(n67922), .A2(n62708), .B1(n68217), .B2(n67914), .ZN(
        n6772) );
  OAI22_X1 U48356 ( .A1(n67922), .A2(n62707), .B1(n68220), .B2(n67914), .ZN(
        n6773) );
  OAI22_X1 U48357 ( .A1(n67922), .A2(n62706), .B1(n68223), .B2(n67914), .ZN(
        n6774) );
  OAI22_X1 U48358 ( .A1(n67922), .A2(n62705), .B1(n68226), .B2(n67914), .ZN(
        n6775) );
  OAI22_X1 U48359 ( .A1(n67922), .A2(n62704), .B1(n68229), .B2(n67914), .ZN(
        n6776) );
  OAI22_X1 U48360 ( .A1(n67922), .A2(n62703), .B1(n68232), .B2(n67914), .ZN(
        n6777) );
  OAI22_X1 U48361 ( .A1(n67922), .A2(n62702), .B1(n68235), .B2(n67914), .ZN(
        n6778) );
  NAND2_X1 U48362 ( .A1(n65076), .A2(n65086), .ZN(n63807) );
  OAI21_X1 U48363 ( .B1(n62156), .B2(n62489), .A(n68052), .ZN(n62493) );
  OAI21_X1 U48364 ( .B1(n62156), .B2(n62223), .A(n68052), .ZN(n62224) );
  OAI21_X1 U48365 ( .B1(n62156), .B2(n62356), .A(n68052), .ZN(n62357) );
  OAI21_X1 U48366 ( .B1(n62088), .B2(n62356), .A(n68052), .ZN(n62290) );
  OAI21_X1 U48367 ( .B1(n62088), .B2(n62223), .A(n68052), .ZN(n62157) );
  OAI21_X1 U48368 ( .B1(n62088), .B2(n62489), .A(n68052), .ZN(n62423) );
  NAND2_X1 U48369 ( .A1(n65087), .A2(n65074), .ZN(n63785) );
  BUF_X1 U48370 ( .A(n62086), .Z(n68060) );
  BUF_X1 U48371 ( .A(n62084), .Z(n68063) );
  BUF_X1 U48372 ( .A(n62082), .Z(n68066) );
  BUF_X1 U48373 ( .A(n62080), .Z(n68069) );
  BUF_X1 U48374 ( .A(n62078), .Z(n68072) );
  BUF_X1 U48375 ( .A(n62076), .Z(n68075) );
  BUF_X1 U48376 ( .A(n62074), .Z(n68078) );
  BUF_X1 U48377 ( .A(n62072), .Z(n68081) );
  BUF_X1 U48378 ( .A(n62070), .Z(n68084) );
  BUF_X1 U48379 ( .A(n62068), .Z(n68087) );
  BUF_X1 U48380 ( .A(n62066), .Z(n68090) );
  BUF_X1 U48381 ( .A(n62064), .Z(n68093) );
  BUF_X1 U48382 ( .A(n62062), .Z(n68096) );
  BUF_X1 U48383 ( .A(n62060), .Z(n68099) );
  BUF_X1 U48384 ( .A(n62058), .Z(n68102) );
  BUF_X1 U48385 ( .A(n62056), .Z(n68105) );
  BUF_X1 U48386 ( .A(n62054), .Z(n68108) );
  BUF_X1 U48387 ( .A(n62052), .Z(n68111) );
  BUF_X1 U48388 ( .A(n62050), .Z(n68114) );
  BUF_X1 U48389 ( .A(n62048), .Z(n68117) );
  BUF_X1 U48390 ( .A(n62046), .Z(n68120) );
  BUF_X1 U48391 ( .A(n62044), .Z(n68123) );
  BUF_X1 U48392 ( .A(n62042), .Z(n68126) );
  BUF_X1 U48393 ( .A(n62040), .Z(n68129) );
  BUF_X1 U48394 ( .A(n62038), .Z(n68132) );
  BUF_X1 U48395 ( .A(n62036), .Z(n68135) );
  BUF_X1 U48396 ( .A(n62034), .Z(n68138) );
  BUF_X1 U48397 ( .A(n62032), .Z(n68141) );
  BUF_X1 U48398 ( .A(n62030), .Z(n68144) );
  BUF_X1 U48399 ( .A(n62028), .Z(n68147) );
  BUF_X1 U48400 ( .A(n62026), .Z(n68150) );
  BUF_X1 U48401 ( .A(n62024), .Z(n68153) );
  BUF_X1 U48402 ( .A(n62022), .Z(n68156) );
  BUF_X1 U48403 ( .A(n62020), .Z(n68159) );
  BUF_X1 U48404 ( .A(n62018), .Z(n68162) );
  BUF_X1 U48405 ( .A(n62016), .Z(n68165) );
  BUF_X1 U48406 ( .A(n62014), .Z(n68168) );
  BUF_X1 U48407 ( .A(n62012), .Z(n68171) );
  BUF_X1 U48408 ( .A(n62010), .Z(n68174) );
  BUF_X1 U48409 ( .A(n62008), .Z(n68177) );
  BUF_X1 U48410 ( .A(n62006), .Z(n68180) );
  BUF_X1 U48411 ( .A(n62004), .Z(n68183) );
  BUF_X1 U48412 ( .A(n62002), .Z(n68186) );
  BUF_X1 U48413 ( .A(n62000), .Z(n68189) );
  BUF_X1 U48414 ( .A(n61998), .Z(n68192) );
  BUF_X1 U48415 ( .A(n61996), .Z(n68195) );
  BUF_X1 U48416 ( .A(n61994), .Z(n68198) );
  BUF_X1 U48417 ( .A(n61992), .Z(n68201) );
  BUF_X1 U48418 ( .A(n61990), .Z(n68204) );
  BUF_X1 U48419 ( .A(n61988), .Z(n68207) );
  BUF_X1 U48420 ( .A(n61986), .Z(n68210) );
  BUF_X1 U48421 ( .A(n61984), .Z(n68213) );
  BUF_X1 U48422 ( .A(n61982), .Z(n68216) );
  BUF_X1 U48423 ( .A(n61980), .Z(n68219) );
  BUF_X1 U48424 ( .A(n61978), .Z(n68222) );
  BUF_X1 U48425 ( .A(n61976), .Z(n68225) );
  BUF_X1 U48426 ( .A(n61974), .Z(n68228) );
  BUF_X1 U48427 ( .A(n61972), .Z(n68231) );
  BUF_X1 U48428 ( .A(n61970), .Z(n68234) );
  BUF_X1 U48429 ( .A(n61968), .Z(n68237) );
  BUF_X1 U48430 ( .A(n61966), .Z(n68240) );
  BUF_X1 U48431 ( .A(n61964), .Z(n68243) );
  BUF_X1 U48432 ( .A(n61962), .Z(n68246) );
  BUF_X1 U48433 ( .A(n61960), .Z(n68249) );
  OAI21_X1 U48434 ( .B1(n62489), .B2(n62625), .A(n68053), .ZN(n62826) );
  OAI21_X1 U48435 ( .B1(n62356), .B2(n63495), .A(n68053), .ZN(n63632) );
  OAI21_X1 U48436 ( .B1(n62089), .B2(n62692), .A(n68052), .ZN(n62626) );
  OAI21_X1 U48437 ( .B1(n62089), .B2(n62625), .A(n68052), .ZN(n62559) );
  OAI21_X1 U48438 ( .B1(n62356), .B2(n63025), .A(n68053), .ZN(n63161) );
  OAI21_X1 U48439 ( .B1(n62089), .B2(n63495), .A(n68054), .ZN(n63429) );
  OAI21_X1 U48440 ( .B1(n62489), .B2(n63495), .A(n68053), .ZN(n63764) );
  OAI21_X1 U48441 ( .B1(n62489), .B2(n63025), .A(n68054), .ZN(n63229) );
  OAI21_X1 U48442 ( .B1(n62223), .B2(n63495), .A(n68054), .ZN(n63500) );
  OAI21_X1 U48443 ( .B1(n62089), .B2(n63092), .A(n68053), .ZN(n63026) );
  OAI21_X1 U48444 ( .B1(n62089), .B2(n63428), .A(n68054), .ZN(n63362) );
  OAI21_X1 U48445 ( .B1(n62223), .B2(n63092), .A(n68053), .ZN(n63095) );
  OAI21_X1 U48446 ( .B1(n62489), .B2(n63428), .A(n68054), .ZN(n63698) );
  OAI21_X1 U48447 ( .B1(n62489), .B2(n63092), .A(n68054), .ZN(n63296) );
  OAI21_X1 U48448 ( .B1(n62356), .B2(n63428), .A(n68054), .ZN(n63566) );
  OAI21_X1 U48449 ( .B1(n62489), .B2(n62692), .A(n68053), .ZN(n62892) );
  OAI21_X1 U48450 ( .B1(n62356), .B2(n62692), .A(n68053), .ZN(n62764) );
  OAI21_X1 U48451 ( .B1(n62223), .B2(n62692), .A(n68052), .ZN(n62696) );
  OAI21_X1 U48452 ( .B1(n62089), .B2(n62156), .A(n68052), .ZN(n62090) );
  NAND2_X1 U48453 ( .A1(n65075), .A2(n65082), .ZN(n63780) );
  NAND2_X1 U48454 ( .A1(n65074), .A2(n65081), .ZN(n63809) );
  NAND2_X1 U48455 ( .A1(n65075), .A2(n65073), .ZN(n63791) );
  AND2_X1 U48456 ( .A1(n66281), .A2(n66279), .ZN(n65117) );
  AND2_X1 U48457 ( .A1(n66281), .A2(n66287), .ZN(n65146) );
  AND2_X1 U48458 ( .A1(n65085), .A2(n65078), .ZN(n63794) );
  AND2_X1 U48459 ( .A1(n65080), .A2(n65086), .ZN(n63795) );
  AND2_X1 U48460 ( .A1(n65073), .A2(n65086), .ZN(n63788) );
  AND2_X1 U48461 ( .A1(n65082), .A2(n65078), .ZN(n63811) );
  AND2_X1 U48462 ( .A1(n65087), .A2(n65078), .ZN(n63815) );
  AND2_X1 U48463 ( .A1(n65087), .A2(n65086), .ZN(n63816) );
  AND2_X1 U48464 ( .A1(n66286), .A2(n66278), .ZN(n65121) );
  AND2_X1 U48465 ( .A1(n66289), .A2(n66278), .ZN(n65126) );
  AND2_X1 U48466 ( .A1(n66285), .A2(n66278), .ZN(n65142) );
  AND2_X1 U48467 ( .A1(n66285), .A2(n66281), .ZN(n65122) );
  AND2_X1 U48468 ( .A1(n66289), .A2(n66281), .ZN(n65127) );
  AND2_X1 U48469 ( .A1(n66280), .A2(n66277), .ZN(n65116) );
  AND2_X1 U48470 ( .A1(n66285), .A2(n66277), .ZN(n65141) );
  AND2_X1 U48471 ( .A1(n66286), .A2(n66277), .ZN(n65147) );
  AND2_X1 U48472 ( .A1(n65077), .A2(n65074), .ZN(n63810) );
  AND2_X1 U48473 ( .A1(n65073), .A2(n65074), .ZN(n63778) );
  AND2_X1 U48474 ( .A1(n65080), .A2(n65074), .ZN(n63783) );
  AND2_X1 U48475 ( .A1(n65074), .A2(n65076), .ZN(n63784) );
  NOR3_X1 U48476 ( .A1(n66297), .A2(ADD_RD2[3]), .A3(n66291), .ZN(n66290) );
  NOR3_X1 U48477 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n65094), .ZN(n65081)
         );
  NOR3_X1 U48478 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n66292), .ZN(n66279)
         );
  NOR3_X1 U48479 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(
        n66287) );
  NOR3_X1 U48480 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n65095), .ZN(n65076)
         );
  NOR3_X1 U48481 ( .A1(n65095), .A2(ADD_RD1[0]), .A3(n65093), .ZN(n65077) );
  NOR3_X1 U48482 ( .A1(n65094), .A2(ADD_RD1[3]), .A3(n65095), .ZN(n65082) );
  NOR3_X1 U48483 ( .A1(n66291), .A2(ADD_RD2[0]), .A3(n66292), .ZN(n66280) );
  NOR3_X1 U48484 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n65093), .ZN(n65073)
         );
  NOR3_X1 U48485 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(
        n65087) );
  NOR3_X1 U48486 ( .A1(n66297), .A2(ADD_RD2[4]), .A3(n66292), .ZN(n66289) );
  NOR3_X1 U48487 ( .A1(n65094), .A2(ADD_RD1[4]), .A3(n65093), .ZN(n65080) );
  NOR3_X1 U48488 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n66297), .ZN(n66286)
         );
  NOR3_X1 U48489 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n66291), .ZN(n66285)
         );
  NOR4_X1 U48490 ( .A1(n66271), .A2(n66272), .A3(n66273), .A4(n66274), .ZN(
        n66270) );
  OAI221_X1 U48491 ( .B1(n63631), .B2(n67380), .C1(n7489), .C2(n67374), .A(
        n66288), .ZN(n66271) );
  OAI221_X1 U48492 ( .B1(n62488), .B2(n67404), .C1(n63697), .C2(n67398), .A(
        n66284), .ZN(n66272) );
  OAI221_X1 U48493 ( .B1(n54670), .B2(n67428), .C1(n63565), .C2(n67422), .A(
        n66282), .ZN(n66273) );
  NOR4_X1 U48494 ( .A1(n66253), .A2(n66254), .A3(n66255), .A4(n66256), .ZN(
        n66252) );
  OAI221_X1 U48495 ( .B1(n63630), .B2(n67380), .C1(n7505), .C2(n67374), .A(
        n66260), .ZN(n66253) );
  OAI221_X1 U48496 ( .B1(n62487), .B2(n67404), .C1(n63696), .C2(n67398), .A(
        n66259), .ZN(n66254) );
  OAI221_X1 U48497 ( .B1(n54669), .B2(n67428), .C1(n63564), .C2(n67422), .A(
        n66258), .ZN(n66255) );
  NOR4_X1 U48498 ( .A1(n66235), .A2(n66236), .A3(n66237), .A4(n66238), .ZN(
        n66234) );
  OAI221_X1 U48499 ( .B1(n63629), .B2(n67380), .C1(n7521), .C2(n67374), .A(
        n66242), .ZN(n66235) );
  OAI221_X1 U48500 ( .B1(n62486), .B2(n67404), .C1(n63695), .C2(n67398), .A(
        n66241), .ZN(n66236) );
  OAI221_X1 U48501 ( .B1(n54668), .B2(n67428), .C1(n63563), .C2(n67422), .A(
        n66240), .ZN(n66237) );
  NOR4_X1 U48502 ( .A1(n66217), .A2(n66218), .A3(n66219), .A4(n66220), .ZN(
        n66216) );
  OAI221_X1 U48503 ( .B1(n63628), .B2(n67380), .C1(n7537), .C2(n67374), .A(
        n66224), .ZN(n66217) );
  OAI221_X1 U48504 ( .B1(n62485), .B2(n67404), .C1(n63694), .C2(n67398), .A(
        n66223), .ZN(n66218) );
  OAI221_X1 U48505 ( .B1(n54667), .B2(n67428), .C1(n63562), .C2(n67422), .A(
        n66222), .ZN(n66219) );
  NOR4_X1 U48506 ( .A1(n66199), .A2(n66200), .A3(n66201), .A4(n66202), .ZN(
        n66198) );
  OAI221_X1 U48507 ( .B1(n63627), .B2(n67380), .C1(n7553), .C2(n67374), .A(
        n66206), .ZN(n66199) );
  OAI221_X1 U48508 ( .B1(n62484), .B2(n67404), .C1(n63693), .C2(n67398), .A(
        n66205), .ZN(n66200) );
  OAI221_X1 U48509 ( .B1(n54666), .B2(n67428), .C1(n63561), .C2(n67422), .A(
        n66204), .ZN(n66201) );
  NOR4_X1 U48510 ( .A1(n66181), .A2(n66182), .A3(n66183), .A4(n66184), .ZN(
        n66180) );
  OAI221_X1 U48511 ( .B1(n63626), .B2(n67380), .C1(n7569), .C2(n67374), .A(
        n66188), .ZN(n66181) );
  OAI221_X1 U48512 ( .B1(n62483), .B2(n67404), .C1(n63692), .C2(n67398), .A(
        n66187), .ZN(n66182) );
  OAI221_X1 U48513 ( .B1(n54665), .B2(n67428), .C1(n63560), .C2(n67422), .A(
        n66186), .ZN(n66183) );
  NOR4_X1 U48514 ( .A1(n66163), .A2(n66164), .A3(n66165), .A4(n66166), .ZN(
        n66162) );
  OAI221_X1 U48515 ( .B1(n63625), .B2(n67380), .C1(n7585), .C2(n67374), .A(
        n66170), .ZN(n66163) );
  OAI221_X1 U48516 ( .B1(n62482), .B2(n67404), .C1(n63691), .C2(n67398), .A(
        n66169), .ZN(n66164) );
  OAI221_X1 U48517 ( .B1(n54664), .B2(n67428), .C1(n63559), .C2(n67422), .A(
        n66168), .ZN(n66165) );
  NOR4_X1 U48518 ( .A1(n66145), .A2(n66146), .A3(n66147), .A4(n66148), .ZN(
        n66144) );
  OAI221_X1 U48519 ( .B1(n63624), .B2(n67380), .C1(n7601), .C2(n67374), .A(
        n66152), .ZN(n66145) );
  OAI221_X1 U48520 ( .B1(n62481), .B2(n67404), .C1(n63690), .C2(n67398), .A(
        n66151), .ZN(n66146) );
  OAI221_X1 U48521 ( .B1(n54663), .B2(n67428), .C1(n63558), .C2(n67422), .A(
        n66150), .ZN(n66147) );
  NOR4_X1 U48522 ( .A1(n66127), .A2(n66128), .A3(n66129), .A4(n66130), .ZN(
        n66126) );
  OAI221_X1 U48523 ( .B1(n63623), .B2(n67380), .C1(n7617), .C2(n67374), .A(
        n66134), .ZN(n66127) );
  OAI221_X1 U48524 ( .B1(n62480), .B2(n67404), .C1(n63689), .C2(n67398), .A(
        n66133), .ZN(n66128) );
  OAI221_X1 U48525 ( .B1(n54662), .B2(n67428), .C1(n63557), .C2(n67422), .A(
        n66132), .ZN(n66129) );
  NOR4_X1 U48526 ( .A1(n66109), .A2(n66110), .A3(n66111), .A4(n66112), .ZN(
        n66108) );
  OAI221_X1 U48527 ( .B1(n63622), .B2(n67380), .C1(n7633), .C2(n67374), .A(
        n66116), .ZN(n66109) );
  OAI221_X1 U48528 ( .B1(n62479), .B2(n67404), .C1(n63688), .C2(n67398), .A(
        n66115), .ZN(n66110) );
  OAI221_X1 U48529 ( .B1(n54661), .B2(n67428), .C1(n63556), .C2(n67422), .A(
        n66114), .ZN(n66111) );
  NOR4_X1 U48530 ( .A1(n66091), .A2(n66092), .A3(n66093), .A4(n66094), .ZN(
        n66090) );
  OAI221_X1 U48531 ( .B1(n63621), .B2(n67380), .C1(n7649), .C2(n67374), .A(
        n66098), .ZN(n66091) );
  OAI221_X1 U48532 ( .B1(n62478), .B2(n67404), .C1(n63687), .C2(n67398), .A(
        n66097), .ZN(n66092) );
  OAI221_X1 U48533 ( .B1(n54660), .B2(n67428), .C1(n63555), .C2(n67422), .A(
        n66096), .ZN(n66093) );
  NOR4_X1 U48534 ( .A1(n66073), .A2(n66074), .A3(n66075), .A4(n66076), .ZN(
        n66072) );
  OAI221_X1 U48535 ( .B1(n63620), .B2(n67380), .C1(n7665), .C2(n67374), .A(
        n66080), .ZN(n66073) );
  OAI221_X1 U48536 ( .B1(n62477), .B2(n67404), .C1(n63686), .C2(n67398), .A(
        n66079), .ZN(n66074) );
  OAI221_X1 U48537 ( .B1(n54659), .B2(n67428), .C1(n63554), .C2(n67422), .A(
        n66078), .ZN(n66075) );
  NOR4_X1 U48538 ( .A1(n66055), .A2(n66056), .A3(n66057), .A4(n66058), .ZN(
        n66054) );
  OAI221_X1 U48539 ( .B1(n63619), .B2(n67381), .C1(n7681), .C2(n67375), .A(
        n66062), .ZN(n66055) );
  OAI221_X1 U48540 ( .B1(n62476), .B2(n67405), .C1(n63685), .C2(n67399), .A(
        n66061), .ZN(n66056) );
  OAI221_X1 U48541 ( .B1(n63415), .B2(n67453), .C1(n49244), .C2(n67447), .A(
        n66059), .ZN(n66058) );
  NOR4_X1 U48542 ( .A1(n66037), .A2(n66038), .A3(n66039), .A4(n66040), .ZN(
        n66036) );
  OAI221_X1 U48543 ( .B1(n63618), .B2(n67381), .C1(n7697), .C2(n67375), .A(
        n66044), .ZN(n66037) );
  OAI221_X1 U48544 ( .B1(n62475), .B2(n67405), .C1(n63684), .C2(n67399), .A(
        n66043), .ZN(n66038) );
  OAI221_X1 U48545 ( .B1(n63414), .B2(n67453), .C1(n49245), .C2(n67447), .A(
        n66041), .ZN(n66040) );
  NOR4_X1 U48546 ( .A1(n66019), .A2(n66020), .A3(n66021), .A4(n66022), .ZN(
        n66018) );
  OAI221_X1 U48547 ( .B1(n63617), .B2(n67381), .C1(n7713), .C2(n67375), .A(
        n66026), .ZN(n66019) );
  OAI221_X1 U48548 ( .B1(n62474), .B2(n67405), .C1(n63683), .C2(n67399), .A(
        n66025), .ZN(n66020) );
  OAI221_X1 U48549 ( .B1(n63413), .B2(n67453), .C1(n49246), .C2(n67447), .A(
        n66023), .ZN(n66022) );
  NOR4_X1 U48550 ( .A1(n66001), .A2(n66002), .A3(n66003), .A4(n66004), .ZN(
        n66000) );
  OAI221_X1 U48551 ( .B1(n63616), .B2(n67381), .C1(n7729), .C2(n67375), .A(
        n66008), .ZN(n66001) );
  OAI221_X1 U48552 ( .B1(n62473), .B2(n67405), .C1(n63682), .C2(n67399), .A(
        n66007), .ZN(n66002) );
  OAI221_X1 U48553 ( .B1(n63412), .B2(n67453), .C1(n49247), .C2(n67447), .A(
        n66005), .ZN(n66004) );
  NOR4_X1 U48554 ( .A1(n65983), .A2(n65984), .A3(n65985), .A4(n65986), .ZN(
        n65982) );
  OAI221_X1 U48555 ( .B1(n63615), .B2(n67381), .C1(n7745), .C2(n67375), .A(
        n65990), .ZN(n65983) );
  OAI221_X1 U48556 ( .B1(n62472), .B2(n67405), .C1(n63681), .C2(n67399), .A(
        n65989), .ZN(n65984) );
  OAI221_X1 U48557 ( .B1(n63411), .B2(n67453), .C1(n49248), .C2(n67447), .A(
        n65987), .ZN(n65986) );
  NOR4_X1 U48558 ( .A1(n65965), .A2(n65966), .A3(n65967), .A4(n65968), .ZN(
        n65964) );
  OAI221_X1 U48559 ( .B1(n63614), .B2(n67381), .C1(n7761), .C2(n67375), .A(
        n65972), .ZN(n65965) );
  OAI221_X1 U48560 ( .B1(n62471), .B2(n67405), .C1(n63680), .C2(n67399), .A(
        n65971), .ZN(n65966) );
  OAI221_X1 U48561 ( .B1(n63410), .B2(n67453), .C1(n49249), .C2(n67447), .A(
        n65969), .ZN(n65968) );
  NOR4_X1 U48562 ( .A1(n65947), .A2(n65948), .A3(n65949), .A4(n65950), .ZN(
        n65946) );
  OAI221_X1 U48563 ( .B1(n63613), .B2(n67381), .C1(n7777), .C2(n67375), .A(
        n65954), .ZN(n65947) );
  OAI221_X1 U48564 ( .B1(n62470), .B2(n67405), .C1(n63679), .C2(n67399), .A(
        n65953), .ZN(n65948) );
  OAI221_X1 U48565 ( .B1(n63409), .B2(n67453), .C1(n49250), .C2(n67447), .A(
        n65951), .ZN(n65950) );
  NOR4_X1 U48566 ( .A1(n65929), .A2(n65930), .A3(n65931), .A4(n65932), .ZN(
        n65928) );
  OAI221_X1 U48567 ( .B1(n63612), .B2(n67381), .C1(n7793), .C2(n67375), .A(
        n65936), .ZN(n65929) );
  OAI221_X1 U48568 ( .B1(n62469), .B2(n67405), .C1(n63678), .C2(n67399), .A(
        n65935), .ZN(n65930) );
  OAI221_X1 U48569 ( .B1(n63408), .B2(n67453), .C1(n49251), .C2(n67447), .A(
        n65933), .ZN(n65932) );
  NOR4_X1 U48570 ( .A1(n65911), .A2(n65912), .A3(n65913), .A4(n65914), .ZN(
        n65910) );
  OAI221_X1 U48571 ( .B1(n63611), .B2(n67381), .C1(n7809), .C2(n67375), .A(
        n65918), .ZN(n65911) );
  OAI221_X1 U48572 ( .B1(n62468), .B2(n67405), .C1(n63677), .C2(n67399), .A(
        n65917), .ZN(n65912) );
  OAI221_X1 U48573 ( .B1(n63407), .B2(n67453), .C1(n49252), .C2(n67447), .A(
        n65915), .ZN(n65914) );
  NOR4_X1 U48574 ( .A1(n65893), .A2(n65894), .A3(n65895), .A4(n65896), .ZN(
        n65892) );
  OAI221_X1 U48575 ( .B1(n63610), .B2(n67381), .C1(n7825), .C2(n67375), .A(
        n65900), .ZN(n65893) );
  OAI221_X1 U48576 ( .B1(n62467), .B2(n67405), .C1(n63676), .C2(n67399), .A(
        n65899), .ZN(n65894) );
  OAI221_X1 U48577 ( .B1(n63406), .B2(n67453), .C1(n49253), .C2(n67447), .A(
        n65897), .ZN(n65896) );
  NOR4_X1 U48578 ( .A1(n65875), .A2(n65876), .A3(n65877), .A4(n65878), .ZN(
        n65874) );
  OAI221_X1 U48579 ( .B1(n63609), .B2(n67381), .C1(n7841), .C2(n67375), .A(
        n65882), .ZN(n65875) );
  OAI221_X1 U48580 ( .B1(n62466), .B2(n67405), .C1(n63675), .C2(n67399), .A(
        n65881), .ZN(n65876) );
  OAI221_X1 U48581 ( .B1(n63405), .B2(n67453), .C1(n49254), .C2(n67447), .A(
        n65879), .ZN(n65878) );
  NOR4_X1 U48582 ( .A1(n65857), .A2(n65858), .A3(n65859), .A4(n65860), .ZN(
        n65856) );
  OAI221_X1 U48583 ( .B1(n63608), .B2(n67381), .C1(n7857), .C2(n67375), .A(
        n65864), .ZN(n65857) );
  OAI221_X1 U48584 ( .B1(n62465), .B2(n67405), .C1(n63674), .C2(n67399), .A(
        n65863), .ZN(n65858) );
  OAI221_X1 U48585 ( .B1(n63404), .B2(n67453), .C1(n49255), .C2(n67447), .A(
        n65861), .ZN(n65860) );
  NOR4_X1 U48586 ( .A1(n65839), .A2(n65840), .A3(n65841), .A4(n65842), .ZN(
        n65838) );
  OAI221_X1 U48587 ( .B1(n63607), .B2(n67382), .C1(n7873), .C2(n67376), .A(
        n65846), .ZN(n65839) );
  OAI221_X1 U48588 ( .B1(n62464), .B2(n67406), .C1(n63673), .C2(n67400), .A(
        n65845), .ZN(n65840) );
  OAI221_X1 U48589 ( .B1(n63403), .B2(n67454), .C1(n49256), .C2(n67448), .A(
        n65843), .ZN(n65842) );
  NOR4_X1 U48590 ( .A1(n65821), .A2(n65822), .A3(n65823), .A4(n65824), .ZN(
        n65820) );
  OAI221_X1 U48591 ( .B1(n63606), .B2(n67382), .C1(n7889), .C2(n67376), .A(
        n65828), .ZN(n65821) );
  OAI221_X1 U48592 ( .B1(n62463), .B2(n67406), .C1(n63672), .C2(n67400), .A(
        n65827), .ZN(n65822) );
  OAI221_X1 U48593 ( .B1(n63402), .B2(n67454), .C1(n49257), .C2(n67448), .A(
        n65825), .ZN(n65824) );
  NOR4_X1 U48594 ( .A1(n65803), .A2(n65804), .A3(n65805), .A4(n65806), .ZN(
        n65802) );
  OAI221_X1 U48595 ( .B1(n63605), .B2(n67382), .C1(n7905), .C2(n67376), .A(
        n65810), .ZN(n65803) );
  OAI221_X1 U48596 ( .B1(n62462), .B2(n67406), .C1(n63671), .C2(n67400), .A(
        n65809), .ZN(n65804) );
  OAI221_X1 U48597 ( .B1(n63401), .B2(n67454), .C1(n49258), .C2(n67448), .A(
        n65807), .ZN(n65806) );
  NOR4_X1 U48598 ( .A1(n65785), .A2(n65786), .A3(n65787), .A4(n65788), .ZN(
        n65784) );
  OAI221_X1 U48599 ( .B1(n63604), .B2(n67382), .C1(n7921), .C2(n67376), .A(
        n65792), .ZN(n65785) );
  OAI221_X1 U48600 ( .B1(n62461), .B2(n67406), .C1(n63670), .C2(n67400), .A(
        n65791), .ZN(n65786) );
  OAI221_X1 U48601 ( .B1(n63400), .B2(n67454), .C1(n49259), .C2(n67448), .A(
        n65789), .ZN(n65788) );
  NOR4_X1 U48602 ( .A1(n65767), .A2(n65768), .A3(n65769), .A4(n65770), .ZN(
        n65766) );
  OAI221_X1 U48603 ( .B1(n63603), .B2(n67382), .C1(n7937), .C2(n67376), .A(
        n65774), .ZN(n65767) );
  OAI221_X1 U48604 ( .B1(n62460), .B2(n67406), .C1(n63669), .C2(n67400), .A(
        n65773), .ZN(n65768) );
  OAI221_X1 U48605 ( .B1(n63399), .B2(n67454), .C1(n49260), .C2(n67448), .A(
        n65771), .ZN(n65770) );
  NOR4_X1 U48606 ( .A1(n65749), .A2(n65750), .A3(n65751), .A4(n65752), .ZN(
        n65748) );
  OAI221_X1 U48607 ( .B1(n63602), .B2(n67382), .C1(n7953), .C2(n67376), .A(
        n65756), .ZN(n65749) );
  OAI221_X1 U48608 ( .B1(n62459), .B2(n67406), .C1(n63668), .C2(n67400), .A(
        n65755), .ZN(n65750) );
  OAI221_X1 U48609 ( .B1(n63398), .B2(n67454), .C1(n49261), .C2(n67448), .A(
        n65753), .ZN(n65752) );
  NOR4_X1 U48610 ( .A1(n65731), .A2(n65732), .A3(n65733), .A4(n65734), .ZN(
        n65730) );
  OAI221_X1 U48611 ( .B1(n63601), .B2(n67382), .C1(n7969), .C2(n67376), .A(
        n65738), .ZN(n65731) );
  OAI221_X1 U48612 ( .B1(n62458), .B2(n67406), .C1(n63667), .C2(n67400), .A(
        n65737), .ZN(n65732) );
  OAI221_X1 U48613 ( .B1(n63397), .B2(n67454), .C1(n49262), .C2(n67448), .A(
        n65735), .ZN(n65734) );
  NOR4_X1 U48614 ( .A1(n65713), .A2(n65714), .A3(n65715), .A4(n65716), .ZN(
        n65712) );
  OAI221_X1 U48615 ( .B1(n63600), .B2(n67382), .C1(n7985), .C2(n67376), .A(
        n65720), .ZN(n65713) );
  OAI221_X1 U48616 ( .B1(n62457), .B2(n67406), .C1(n63666), .C2(n67400), .A(
        n65719), .ZN(n65714) );
  OAI221_X1 U48617 ( .B1(n63396), .B2(n67454), .C1(n49263), .C2(n67448), .A(
        n65717), .ZN(n65716) );
  NOR4_X1 U48618 ( .A1(n65695), .A2(n65696), .A3(n65697), .A4(n65698), .ZN(
        n65694) );
  OAI221_X1 U48619 ( .B1(n63599), .B2(n67382), .C1(n8001), .C2(n67376), .A(
        n65702), .ZN(n65695) );
  OAI221_X1 U48620 ( .B1(n62456), .B2(n67406), .C1(n63665), .C2(n67400), .A(
        n65701), .ZN(n65696) );
  OAI221_X1 U48621 ( .B1(n63395), .B2(n67454), .C1(n49264), .C2(n67448), .A(
        n65699), .ZN(n65698) );
  NOR4_X1 U48622 ( .A1(n65677), .A2(n65678), .A3(n65679), .A4(n65680), .ZN(
        n65676) );
  OAI221_X1 U48623 ( .B1(n63598), .B2(n67382), .C1(n8017), .C2(n67376), .A(
        n65684), .ZN(n65677) );
  OAI221_X1 U48624 ( .B1(n62455), .B2(n67406), .C1(n63664), .C2(n67400), .A(
        n65683), .ZN(n65678) );
  OAI221_X1 U48625 ( .B1(n63394), .B2(n67454), .C1(n49265), .C2(n67448), .A(
        n65681), .ZN(n65680) );
  NOR4_X1 U48626 ( .A1(n65659), .A2(n65660), .A3(n65661), .A4(n65662), .ZN(
        n65658) );
  OAI221_X1 U48627 ( .B1(n63597), .B2(n67382), .C1(n8033), .C2(n67376), .A(
        n65666), .ZN(n65659) );
  OAI221_X1 U48628 ( .B1(n62454), .B2(n67406), .C1(n63663), .C2(n67400), .A(
        n65665), .ZN(n65660) );
  OAI221_X1 U48629 ( .B1(n63393), .B2(n67454), .C1(n49266), .C2(n67448), .A(
        n65663), .ZN(n65662) );
  NOR4_X1 U48630 ( .A1(n65641), .A2(n65642), .A3(n65643), .A4(n65644), .ZN(
        n65640) );
  OAI221_X1 U48631 ( .B1(n63596), .B2(n67382), .C1(n8049), .C2(n67376), .A(
        n65648), .ZN(n65641) );
  OAI221_X1 U48632 ( .B1(n62453), .B2(n67406), .C1(n63662), .C2(n67400), .A(
        n65647), .ZN(n65642) );
  OAI221_X1 U48633 ( .B1(n63392), .B2(n67454), .C1(n49267), .C2(n67448), .A(
        n65645), .ZN(n65644) );
  NOR4_X1 U48634 ( .A1(n65623), .A2(n65624), .A3(n65625), .A4(n65626), .ZN(
        n65622) );
  OAI221_X1 U48635 ( .B1(n63595), .B2(n67383), .C1(n8065), .C2(n67377), .A(
        n65630), .ZN(n65623) );
  OAI221_X1 U48636 ( .B1(n62452), .B2(n67407), .C1(n63661), .C2(n67401), .A(
        n65629), .ZN(n65624) );
  OAI221_X1 U48637 ( .B1(n63391), .B2(n67455), .C1(n49268), .C2(n67449), .A(
        n65627), .ZN(n65626) );
  NOR4_X1 U48638 ( .A1(n65605), .A2(n65606), .A3(n65607), .A4(n65608), .ZN(
        n65604) );
  OAI221_X1 U48639 ( .B1(n63594), .B2(n67383), .C1(n8081), .C2(n67377), .A(
        n65612), .ZN(n65605) );
  OAI221_X1 U48640 ( .B1(n62451), .B2(n67407), .C1(n63660), .C2(n67401), .A(
        n65611), .ZN(n65606) );
  OAI221_X1 U48641 ( .B1(n63390), .B2(n67455), .C1(n49269), .C2(n67449), .A(
        n65609), .ZN(n65608) );
  NOR4_X1 U48642 ( .A1(n65587), .A2(n65588), .A3(n65589), .A4(n65590), .ZN(
        n65586) );
  OAI221_X1 U48643 ( .B1(n63593), .B2(n67383), .C1(n8097), .C2(n67377), .A(
        n65594), .ZN(n65587) );
  OAI221_X1 U48644 ( .B1(n62450), .B2(n67407), .C1(n63659), .C2(n67401), .A(
        n65593), .ZN(n65588) );
  OAI221_X1 U48645 ( .B1(n63389), .B2(n67455), .C1(n49270), .C2(n67449), .A(
        n65591), .ZN(n65590) );
  NOR4_X1 U48646 ( .A1(n65569), .A2(n65570), .A3(n65571), .A4(n65572), .ZN(
        n65568) );
  OAI221_X1 U48647 ( .B1(n63592), .B2(n67383), .C1(n8113), .C2(n67377), .A(
        n65576), .ZN(n65569) );
  OAI221_X1 U48648 ( .B1(n62449), .B2(n67407), .C1(n63658), .C2(n67401), .A(
        n65575), .ZN(n65570) );
  OAI221_X1 U48649 ( .B1(n63388), .B2(n67455), .C1(n49271), .C2(n67449), .A(
        n65573), .ZN(n65572) );
  NOR4_X1 U48650 ( .A1(n65551), .A2(n65552), .A3(n65553), .A4(n65554), .ZN(
        n65550) );
  OAI221_X1 U48651 ( .B1(n63591), .B2(n67383), .C1(n8129), .C2(n67377), .A(
        n65558), .ZN(n65551) );
  OAI221_X1 U48652 ( .B1(n62448), .B2(n67407), .C1(n63657), .C2(n67401), .A(
        n65557), .ZN(n65552) );
  OAI221_X1 U48653 ( .B1(n63387), .B2(n67455), .C1(n49272), .C2(n67449), .A(
        n65555), .ZN(n65554) );
  NOR4_X1 U48654 ( .A1(n65533), .A2(n65534), .A3(n65535), .A4(n65536), .ZN(
        n65532) );
  OAI221_X1 U48655 ( .B1(n63590), .B2(n67383), .C1(n8145), .C2(n67377), .A(
        n65540), .ZN(n65533) );
  OAI221_X1 U48656 ( .B1(n62447), .B2(n67407), .C1(n63656), .C2(n67401), .A(
        n65539), .ZN(n65534) );
  OAI221_X1 U48657 ( .B1(n63386), .B2(n67455), .C1(n49273), .C2(n67449), .A(
        n65537), .ZN(n65536) );
  NOR4_X1 U48658 ( .A1(n65515), .A2(n65516), .A3(n65517), .A4(n65518), .ZN(
        n65514) );
  OAI221_X1 U48659 ( .B1(n63589), .B2(n67383), .C1(n8161), .C2(n67377), .A(
        n65522), .ZN(n65515) );
  OAI221_X1 U48660 ( .B1(n62446), .B2(n67407), .C1(n63655), .C2(n67401), .A(
        n65521), .ZN(n65516) );
  OAI221_X1 U48661 ( .B1(n63385), .B2(n67455), .C1(n49274), .C2(n67449), .A(
        n65519), .ZN(n65518) );
  NOR4_X1 U48662 ( .A1(n65497), .A2(n65498), .A3(n65499), .A4(n65500), .ZN(
        n65496) );
  OAI221_X1 U48663 ( .B1(n63588), .B2(n67383), .C1(n8177), .C2(n67377), .A(
        n65504), .ZN(n65497) );
  OAI221_X1 U48664 ( .B1(n62445), .B2(n67407), .C1(n63654), .C2(n67401), .A(
        n65503), .ZN(n65498) );
  OAI221_X1 U48665 ( .B1(n63384), .B2(n67455), .C1(n49275), .C2(n67449), .A(
        n65501), .ZN(n65500) );
  NOR4_X1 U48666 ( .A1(n65479), .A2(n65480), .A3(n65481), .A4(n65482), .ZN(
        n65478) );
  OAI221_X1 U48667 ( .B1(n63587), .B2(n67383), .C1(n8193), .C2(n67377), .A(
        n65486), .ZN(n65479) );
  OAI221_X1 U48668 ( .B1(n62444), .B2(n67407), .C1(n63653), .C2(n67401), .A(
        n65485), .ZN(n65480) );
  OAI221_X1 U48669 ( .B1(n63383), .B2(n67455), .C1(n49276), .C2(n67449), .A(
        n65483), .ZN(n65482) );
  NOR4_X1 U48670 ( .A1(n65461), .A2(n65462), .A3(n65463), .A4(n65464), .ZN(
        n65460) );
  OAI221_X1 U48671 ( .B1(n63586), .B2(n67383), .C1(n8209), .C2(n67377), .A(
        n65468), .ZN(n65461) );
  OAI221_X1 U48672 ( .B1(n62443), .B2(n67407), .C1(n63652), .C2(n67401), .A(
        n65467), .ZN(n65462) );
  OAI221_X1 U48673 ( .B1(n63382), .B2(n67455), .C1(n49277), .C2(n67449), .A(
        n65465), .ZN(n65464) );
  NOR4_X1 U48674 ( .A1(n65443), .A2(n65444), .A3(n65445), .A4(n65446), .ZN(
        n65442) );
  OAI221_X1 U48675 ( .B1(n63585), .B2(n67383), .C1(n8225), .C2(n67377), .A(
        n65450), .ZN(n65443) );
  OAI221_X1 U48676 ( .B1(n62442), .B2(n67407), .C1(n63651), .C2(n67401), .A(
        n65449), .ZN(n65444) );
  OAI221_X1 U48677 ( .B1(n63381), .B2(n67455), .C1(n49278), .C2(n67449), .A(
        n65447), .ZN(n65446) );
  NOR4_X1 U48678 ( .A1(n65425), .A2(n65426), .A3(n65427), .A4(n65428), .ZN(
        n65424) );
  OAI221_X1 U48679 ( .B1(n63584), .B2(n67383), .C1(n8241), .C2(n67377), .A(
        n65432), .ZN(n65425) );
  OAI221_X1 U48680 ( .B1(n62441), .B2(n67407), .C1(n63650), .C2(n67401), .A(
        n65431), .ZN(n65426) );
  OAI221_X1 U48681 ( .B1(n63380), .B2(n67455), .C1(n49279), .C2(n67449), .A(
        n65429), .ZN(n65428) );
  NOR4_X1 U48682 ( .A1(n65407), .A2(n65408), .A3(n65409), .A4(n65410), .ZN(
        n65406) );
  OAI221_X1 U48683 ( .B1(n63583), .B2(n67384), .C1(n8257), .C2(n67378), .A(
        n65414), .ZN(n65407) );
  OAI221_X1 U48684 ( .B1(n62440), .B2(n67408), .C1(n63649), .C2(n67402), .A(
        n65413), .ZN(n65408) );
  OAI221_X1 U48685 ( .B1(n63379), .B2(n67456), .C1(n49280), .C2(n67450), .A(
        n65411), .ZN(n65410) );
  NOR4_X1 U48686 ( .A1(n65389), .A2(n65390), .A3(n65391), .A4(n65392), .ZN(
        n65388) );
  OAI221_X1 U48687 ( .B1(n63582), .B2(n67384), .C1(n8273), .C2(n67378), .A(
        n65396), .ZN(n65389) );
  OAI221_X1 U48688 ( .B1(n62439), .B2(n67408), .C1(n63648), .C2(n67402), .A(
        n65395), .ZN(n65390) );
  OAI221_X1 U48689 ( .B1(n63378), .B2(n67456), .C1(n49281), .C2(n67450), .A(
        n65393), .ZN(n65392) );
  NOR4_X1 U48690 ( .A1(n65371), .A2(n65372), .A3(n65373), .A4(n65374), .ZN(
        n65370) );
  OAI221_X1 U48691 ( .B1(n63581), .B2(n67384), .C1(n8289), .C2(n67378), .A(
        n65378), .ZN(n65371) );
  OAI221_X1 U48692 ( .B1(n62438), .B2(n67408), .C1(n63647), .C2(n67402), .A(
        n65377), .ZN(n65372) );
  OAI221_X1 U48693 ( .B1(n63377), .B2(n67456), .C1(n49282), .C2(n67450), .A(
        n65375), .ZN(n65374) );
  NOR4_X1 U48694 ( .A1(n65353), .A2(n65354), .A3(n65355), .A4(n65356), .ZN(
        n65352) );
  OAI221_X1 U48695 ( .B1(n63580), .B2(n67384), .C1(n8305), .C2(n67378), .A(
        n65360), .ZN(n65353) );
  OAI221_X1 U48696 ( .B1(n62437), .B2(n67408), .C1(n63646), .C2(n67402), .A(
        n65359), .ZN(n65354) );
  OAI221_X1 U48697 ( .B1(n63376), .B2(n67456), .C1(n49283), .C2(n67450), .A(
        n65357), .ZN(n65356) );
  NOR4_X1 U48698 ( .A1(n65335), .A2(n65336), .A3(n65337), .A4(n65338), .ZN(
        n65334) );
  OAI221_X1 U48699 ( .B1(n63579), .B2(n67384), .C1(n8321), .C2(n67378), .A(
        n65342), .ZN(n65335) );
  OAI221_X1 U48700 ( .B1(n62436), .B2(n67408), .C1(n63645), .C2(n67402), .A(
        n65341), .ZN(n65336) );
  OAI221_X1 U48701 ( .B1(n63375), .B2(n67456), .C1(n49284), .C2(n67450), .A(
        n65339), .ZN(n65338) );
  NOR4_X1 U48702 ( .A1(n65317), .A2(n65318), .A3(n65319), .A4(n65320), .ZN(
        n65316) );
  OAI221_X1 U48703 ( .B1(n63578), .B2(n67384), .C1(n8337), .C2(n67378), .A(
        n65324), .ZN(n65317) );
  OAI221_X1 U48704 ( .B1(n62435), .B2(n67408), .C1(n63644), .C2(n67402), .A(
        n65323), .ZN(n65318) );
  OAI221_X1 U48705 ( .B1(n63374), .B2(n67456), .C1(n49285), .C2(n67450), .A(
        n65321), .ZN(n65320) );
  NOR4_X1 U48706 ( .A1(n65299), .A2(n65300), .A3(n65301), .A4(n65302), .ZN(
        n65298) );
  OAI221_X1 U48707 ( .B1(n63577), .B2(n67384), .C1(n8353), .C2(n67378), .A(
        n65306), .ZN(n65299) );
  OAI221_X1 U48708 ( .B1(n62434), .B2(n67408), .C1(n63643), .C2(n67402), .A(
        n65305), .ZN(n65300) );
  OAI221_X1 U48709 ( .B1(n63373), .B2(n67456), .C1(n49286), .C2(n67450), .A(
        n65303), .ZN(n65302) );
  NOR4_X1 U48710 ( .A1(n65281), .A2(n65282), .A3(n65283), .A4(n65284), .ZN(
        n65280) );
  OAI221_X1 U48711 ( .B1(n63576), .B2(n67384), .C1(n8369), .C2(n67378), .A(
        n65288), .ZN(n65281) );
  OAI221_X1 U48712 ( .B1(n62433), .B2(n67408), .C1(n63642), .C2(n67402), .A(
        n65287), .ZN(n65282) );
  OAI221_X1 U48713 ( .B1(n63372), .B2(n67456), .C1(n49287), .C2(n67450), .A(
        n65285), .ZN(n65284) );
  NOR4_X1 U48714 ( .A1(n65263), .A2(n65264), .A3(n65265), .A4(n65266), .ZN(
        n65262) );
  OAI221_X1 U48715 ( .B1(n63575), .B2(n67384), .C1(n8385), .C2(n67378), .A(
        n65270), .ZN(n65263) );
  OAI221_X1 U48716 ( .B1(n62432), .B2(n67408), .C1(n63641), .C2(n67402), .A(
        n65269), .ZN(n65264) );
  OAI221_X1 U48717 ( .B1(n63371), .B2(n67456), .C1(n49288), .C2(n67450), .A(
        n65267), .ZN(n65266) );
  NOR4_X1 U48718 ( .A1(n65245), .A2(n65246), .A3(n65247), .A4(n65248), .ZN(
        n65244) );
  OAI221_X1 U48719 ( .B1(n63574), .B2(n67384), .C1(n8401), .C2(n67378), .A(
        n65252), .ZN(n65245) );
  OAI221_X1 U48720 ( .B1(n62431), .B2(n67408), .C1(n63640), .C2(n67402), .A(
        n65251), .ZN(n65246) );
  OAI221_X1 U48721 ( .B1(n63370), .B2(n67456), .C1(n49289), .C2(n67450), .A(
        n65249), .ZN(n65248) );
  NOR4_X1 U48722 ( .A1(n65227), .A2(n65228), .A3(n65229), .A4(n65230), .ZN(
        n65226) );
  OAI221_X1 U48723 ( .B1(n63573), .B2(n67384), .C1(n8417), .C2(n67378), .A(
        n65234), .ZN(n65227) );
  OAI221_X1 U48724 ( .B1(n62430), .B2(n67408), .C1(n63639), .C2(n67402), .A(
        n65233), .ZN(n65228) );
  OAI221_X1 U48725 ( .B1(n63369), .B2(n67456), .C1(n49290), .C2(n67450), .A(
        n65231), .ZN(n65230) );
  NOR4_X1 U48726 ( .A1(n65209), .A2(n65210), .A3(n65211), .A4(n65212), .ZN(
        n65208) );
  OAI221_X1 U48727 ( .B1(n63572), .B2(n67384), .C1(n8433), .C2(n67378), .A(
        n65216), .ZN(n65209) );
  OAI221_X1 U48728 ( .B1(n62429), .B2(n67408), .C1(n63638), .C2(n67402), .A(
        n65215), .ZN(n65210) );
  OAI221_X1 U48729 ( .B1(n63368), .B2(n67456), .C1(n49291), .C2(n67450), .A(
        n65213), .ZN(n65212) );
  NOR4_X1 U48730 ( .A1(n65068), .A2(n65069), .A3(n65070), .A4(n65071), .ZN(
        n65067) );
  OAI221_X1 U48731 ( .B1(n63160), .B2(n67626), .C1(n62289), .C2(n67620), .A(
        n65079), .ZN(n65070) );
  OAI221_X1 U48732 ( .B1(n63427), .B2(n67648), .C1(n49420), .C2(n67642), .A(
        n65072), .ZN(n65071) );
  OAI221_X1 U48733 ( .B1(n62488), .B2(n67602), .C1(n63565), .C2(n67596), .A(
        n65083), .ZN(n65069) );
  NOR4_X1 U48734 ( .A1(n65048), .A2(n65049), .A3(n65050), .A4(n65051), .ZN(
        n65047) );
  OAI221_X1 U48735 ( .B1(n63159), .B2(n67626), .C1(n62288), .C2(n67620), .A(
        n65053), .ZN(n65050) );
  OAI221_X1 U48736 ( .B1(n63426), .B2(n67648), .C1(n49421), .C2(n67642), .A(
        n65052), .ZN(n65051) );
  OAI221_X1 U48737 ( .B1(n62487), .B2(n67602), .C1(n63564), .C2(n67596), .A(
        n65054), .ZN(n65049) );
  NOR4_X1 U48738 ( .A1(n65028), .A2(n65029), .A3(n65030), .A4(n65031), .ZN(
        n65027) );
  OAI221_X1 U48739 ( .B1(n63158), .B2(n67626), .C1(n62287), .C2(n67620), .A(
        n65033), .ZN(n65030) );
  OAI221_X1 U48740 ( .B1(n63425), .B2(n67648), .C1(n49422), .C2(n67642), .A(
        n65032), .ZN(n65031) );
  OAI221_X1 U48741 ( .B1(n62486), .B2(n67602), .C1(n63563), .C2(n67596), .A(
        n65034), .ZN(n65029) );
  NOR4_X1 U48742 ( .A1(n65008), .A2(n65009), .A3(n65010), .A4(n65011), .ZN(
        n65007) );
  OAI221_X1 U48743 ( .B1(n63157), .B2(n67626), .C1(n62286), .C2(n67620), .A(
        n65013), .ZN(n65010) );
  OAI221_X1 U48744 ( .B1(n63424), .B2(n67648), .C1(n49423), .C2(n67642), .A(
        n65012), .ZN(n65011) );
  OAI221_X1 U48745 ( .B1(n62485), .B2(n67602), .C1(n63562), .C2(n67596), .A(
        n65014), .ZN(n65009) );
  NOR4_X1 U48746 ( .A1(n64988), .A2(n64989), .A3(n64990), .A4(n64991), .ZN(
        n64987) );
  OAI221_X1 U48747 ( .B1(n63156), .B2(n67626), .C1(n62285), .C2(n67620), .A(
        n64993), .ZN(n64990) );
  OAI221_X1 U48748 ( .B1(n63423), .B2(n67648), .C1(n49424), .C2(n67642), .A(
        n64992), .ZN(n64991) );
  OAI221_X1 U48749 ( .B1(n62484), .B2(n67602), .C1(n63561), .C2(n67596), .A(
        n64994), .ZN(n64989) );
  NOR4_X1 U48750 ( .A1(n64968), .A2(n64969), .A3(n64970), .A4(n64971), .ZN(
        n64967) );
  OAI221_X1 U48751 ( .B1(n63155), .B2(n67626), .C1(n62284), .C2(n67620), .A(
        n64973), .ZN(n64970) );
  OAI221_X1 U48752 ( .B1(n63422), .B2(n67648), .C1(n49425), .C2(n67642), .A(
        n64972), .ZN(n64971) );
  OAI221_X1 U48753 ( .B1(n62483), .B2(n67602), .C1(n63560), .C2(n67596), .A(
        n64974), .ZN(n64969) );
  NOR4_X1 U48754 ( .A1(n64948), .A2(n64949), .A3(n64950), .A4(n64951), .ZN(
        n64947) );
  OAI221_X1 U48755 ( .B1(n63154), .B2(n67626), .C1(n62283), .C2(n67620), .A(
        n64953), .ZN(n64950) );
  OAI221_X1 U48756 ( .B1(n63421), .B2(n67648), .C1(n49426), .C2(n67642), .A(
        n64952), .ZN(n64951) );
  OAI221_X1 U48757 ( .B1(n62482), .B2(n67602), .C1(n63559), .C2(n67596), .A(
        n64954), .ZN(n64949) );
  NOR4_X1 U48758 ( .A1(n64928), .A2(n64929), .A3(n64930), .A4(n64931), .ZN(
        n64927) );
  OAI221_X1 U48759 ( .B1(n63153), .B2(n67626), .C1(n62282), .C2(n67620), .A(
        n64933), .ZN(n64930) );
  OAI221_X1 U48760 ( .B1(n63420), .B2(n67648), .C1(n49427), .C2(n67642), .A(
        n64932), .ZN(n64931) );
  OAI221_X1 U48761 ( .B1(n62481), .B2(n67602), .C1(n63558), .C2(n67596), .A(
        n64934), .ZN(n64929) );
  NOR4_X1 U48762 ( .A1(n64908), .A2(n64909), .A3(n64910), .A4(n64911), .ZN(
        n64907) );
  OAI221_X1 U48763 ( .B1(n63152), .B2(n67626), .C1(n62281), .C2(n67620), .A(
        n64913), .ZN(n64910) );
  OAI221_X1 U48764 ( .B1(n63419), .B2(n67648), .C1(n49428), .C2(n67642), .A(
        n64912), .ZN(n64911) );
  OAI221_X1 U48765 ( .B1(n62480), .B2(n67602), .C1(n63557), .C2(n67596), .A(
        n64914), .ZN(n64909) );
  NOR4_X1 U48766 ( .A1(n64888), .A2(n64889), .A3(n64890), .A4(n64891), .ZN(
        n64887) );
  OAI221_X1 U48767 ( .B1(n63151), .B2(n67626), .C1(n62280), .C2(n67620), .A(
        n64893), .ZN(n64890) );
  OAI221_X1 U48768 ( .B1(n63418), .B2(n67648), .C1(n49429), .C2(n67642), .A(
        n64892), .ZN(n64891) );
  OAI221_X1 U48769 ( .B1(n62479), .B2(n67602), .C1(n63556), .C2(n67596), .A(
        n64894), .ZN(n64889) );
  NOR4_X1 U48770 ( .A1(n64868), .A2(n64869), .A3(n64870), .A4(n64871), .ZN(
        n64867) );
  OAI221_X1 U48771 ( .B1(n63150), .B2(n67626), .C1(n62279), .C2(n67620), .A(
        n64873), .ZN(n64870) );
  OAI221_X1 U48772 ( .B1(n63417), .B2(n67648), .C1(n49430), .C2(n67642), .A(
        n64872), .ZN(n64871) );
  OAI221_X1 U48773 ( .B1(n62478), .B2(n67602), .C1(n63555), .C2(n67596), .A(
        n64874), .ZN(n64869) );
  NOR4_X1 U48774 ( .A1(n64848), .A2(n64849), .A3(n64850), .A4(n64851), .ZN(
        n64847) );
  OAI221_X1 U48775 ( .B1(n63149), .B2(n67626), .C1(n62278), .C2(n67620), .A(
        n64853), .ZN(n64850) );
  OAI221_X1 U48776 ( .B1(n63416), .B2(n67648), .C1(n49431), .C2(n67642), .A(
        n64852), .ZN(n64851) );
  OAI221_X1 U48777 ( .B1(n62477), .B2(n67602), .C1(n63554), .C2(n67596), .A(
        n64854), .ZN(n64849) );
  NOR4_X1 U48778 ( .A1(n64828), .A2(n64829), .A3(n64830), .A4(n64831), .ZN(
        n64827) );
  OAI221_X1 U48779 ( .B1(n63148), .B2(n67627), .C1(n62277), .C2(n67621), .A(
        n64833), .ZN(n64830) );
  OAI221_X1 U48780 ( .B1(n62476), .B2(n67603), .C1(n63553), .C2(n67597), .A(
        n64834), .ZN(n64829) );
  OAI221_X1 U48781 ( .B1(n54234), .B2(n67579), .C1(n63619), .C2(n67573), .A(
        n64836), .ZN(n64828) );
  NOR4_X1 U48782 ( .A1(n64808), .A2(n64809), .A3(n64810), .A4(n64811), .ZN(
        n64807) );
  OAI221_X1 U48783 ( .B1(n63147), .B2(n67627), .C1(n62276), .C2(n67621), .A(
        n64813), .ZN(n64810) );
  OAI221_X1 U48784 ( .B1(n62475), .B2(n67603), .C1(n63552), .C2(n67597), .A(
        n64814), .ZN(n64809) );
  OAI221_X1 U48785 ( .B1(n54233), .B2(n67579), .C1(n63618), .C2(n67573), .A(
        n64816), .ZN(n64808) );
  NOR4_X1 U48786 ( .A1(n64788), .A2(n64789), .A3(n64790), .A4(n64791), .ZN(
        n64787) );
  OAI221_X1 U48787 ( .B1(n63146), .B2(n67627), .C1(n62275), .C2(n67621), .A(
        n64793), .ZN(n64790) );
  OAI221_X1 U48788 ( .B1(n62474), .B2(n67603), .C1(n63551), .C2(n67597), .A(
        n64794), .ZN(n64789) );
  OAI221_X1 U48789 ( .B1(n54232), .B2(n67579), .C1(n63617), .C2(n67573), .A(
        n64796), .ZN(n64788) );
  NOR4_X1 U48790 ( .A1(n64768), .A2(n64769), .A3(n64770), .A4(n64771), .ZN(
        n64767) );
  OAI221_X1 U48791 ( .B1(n63145), .B2(n67627), .C1(n62274), .C2(n67621), .A(
        n64773), .ZN(n64770) );
  OAI221_X1 U48792 ( .B1(n62473), .B2(n67603), .C1(n63550), .C2(n67597), .A(
        n64774), .ZN(n64769) );
  OAI221_X1 U48793 ( .B1(n54231), .B2(n67579), .C1(n63616), .C2(n67573), .A(
        n64776), .ZN(n64768) );
  NOR4_X1 U48794 ( .A1(n64748), .A2(n64749), .A3(n64750), .A4(n64751), .ZN(
        n64747) );
  OAI221_X1 U48795 ( .B1(n63144), .B2(n67627), .C1(n62273), .C2(n67621), .A(
        n64753), .ZN(n64750) );
  OAI221_X1 U48796 ( .B1(n62472), .B2(n67603), .C1(n63549), .C2(n67597), .A(
        n64754), .ZN(n64749) );
  OAI221_X1 U48797 ( .B1(n54230), .B2(n67579), .C1(n63615), .C2(n67573), .A(
        n64756), .ZN(n64748) );
  NOR4_X1 U48798 ( .A1(n64728), .A2(n64729), .A3(n64730), .A4(n64731), .ZN(
        n64727) );
  OAI221_X1 U48799 ( .B1(n63143), .B2(n67627), .C1(n62272), .C2(n67621), .A(
        n64733), .ZN(n64730) );
  OAI221_X1 U48800 ( .B1(n62471), .B2(n67603), .C1(n63548), .C2(n67597), .A(
        n64734), .ZN(n64729) );
  OAI221_X1 U48801 ( .B1(n54229), .B2(n67579), .C1(n63614), .C2(n67573), .A(
        n64736), .ZN(n64728) );
  NOR4_X1 U48802 ( .A1(n64708), .A2(n64709), .A3(n64710), .A4(n64711), .ZN(
        n64707) );
  OAI221_X1 U48803 ( .B1(n63142), .B2(n67627), .C1(n62271), .C2(n67621), .A(
        n64713), .ZN(n64710) );
  OAI221_X1 U48804 ( .B1(n62470), .B2(n67603), .C1(n63547), .C2(n67597), .A(
        n64714), .ZN(n64709) );
  OAI221_X1 U48805 ( .B1(n54228), .B2(n67579), .C1(n63613), .C2(n67573), .A(
        n64716), .ZN(n64708) );
  NOR4_X1 U48806 ( .A1(n64688), .A2(n64689), .A3(n64690), .A4(n64691), .ZN(
        n64687) );
  OAI221_X1 U48807 ( .B1(n63141), .B2(n67627), .C1(n62270), .C2(n67621), .A(
        n64693), .ZN(n64690) );
  OAI221_X1 U48808 ( .B1(n62469), .B2(n67603), .C1(n63546), .C2(n67597), .A(
        n64694), .ZN(n64689) );
  OAI221_X1 U48809 ( .B1(n54227), .B2(n67579), .C1(n63612), .C2(n67573), .A(
        n64696), .ZN(n64688) );
  NOR4_X1 U48810 ( .A1(n64668), .A2(n64669), .A3(n64670), .A4(n64671), .ZN(
        n64667) );
  OAI221_X1 U48811 ( .B1(n63140), .B2(n67627), .C1(n62269), .C2(n67621), .A(
        n64673), .ZN(n64670) );
  OAI221_X1 U48812 ( .B1(n62468), .B2(n67603), .C1(n63545), .C2(n67597), .A(
        n64674), .ZN(n64669) );
  OAI221_X1 U48813 ( .B1(n54226), .B2(n67579), .C1(n63611), .C2(n67573), .A(
        n64676), .ZN(n64668) );
  NOR4_X1 U48814 ( .A1(n64648), .A2(n64649), .A3(n64650), .A4(n64651), .ZN(
        n64647) );
  OAI221_X1 U48815 ( .B1(n63139), .B2(n67627), .C1(n62268), .C2(n67621), .A(
        n64653), .ZN(n64650) );
  OAI221_X1 U48816 ( .B1(n62467), .B2(n67603), .C1(n63544), .C2(n67597), .A(
        n64654), .ZN(n64649) );
  OAI221_X1 U48817 ( .B1(n54225), .B2(n67579), .C1(n63610), .C2(n67573), .A(
        n64656), .ZN(n64648) );
  NOR4_X1 U48818 ( .A1(n64628), .A2(n64629), .A3(n64630), .A4(n64631), .ZN(
        n64627) );
  OAI221_X1 U48819 ( .B1(n63138), .B2(n67627), .C1(n62267), .C2(n67621), .A(
        n64633), .ZN(n64630) );
  OAI221_X1 U48820 ( .B1(n62466), .B2(n67603), .C1(n63543), .C2(n67597), .A(
        n64634), .ZN(n64629) );
  OAI221_X1 U48821 ( .B1(n54224), .B2(n67579), .C1(n63609), .C2(n67573), .A(
        n64636), .ZN(n64628) );
  NOR4_X1 U48822 ( .A1(n64608), .A2(n64609), .A3(n64610), .A4(n64611), .ZN(
        n64607) );
  OAI221_X1 U48823 ( .B1(n63137), .B2(n67627), .C1(n62266), .C2(n67621), .A(
        n64613), .ZN(n64610) );
  OAI221_X1 U48824 ( .B1(n62465), .B2(n67603), .C1(n63542), .C2(n67597), .A(
        n64614), .ZN(n64609) );
  OAI221_X1 U48825 ( .B1(n54223), .B2(n67579), .C1(n63608), .C2(n67573), .A(
        n64616), .ZN(n64608) );
  NOR4_X1 U48826 ( .A1(n64588), .A2(n64589), .A3(n64590), .A4(n64591), .ZN(
        n64587) );
  OAI221_X1 U48827 ( .B1(n63136), .B2(n67628), .C1(n62265), .C2(n67622), .A(
        n64593), .ZN(n64590) );
  OAI221_X1 U48828 ( .B1(n62464), .B2(n67604), .C1(n63541), .C2(n67598), .A(
        n64594), .ZN(n64589) );
  OAI221_X1 U48829 ( .B1(n54222), .B2(n67580), .C1(n63607), .C2(n67574), .A(
        n64596), .ZN(n64588) );
  NOR4_X1 U48830 ( .A1(n64568), .A2(n64569), .A3(n64570), .A4(n64571), .ZN(
        n64567) );
  OAI221_X1 U48831 ( .B1(n63135), .B2(n67628), .C1(n62264), .C2(n67622), .A(
        n64573), .ZN(n64570) );
  OAI221_X1 U48832 ( .B1(n62463), .B2(n67604), .C1(n63540), .C2(n67598), .A(
        n64574), .ZN(n64569) );
  OAI221_X1 U48833 ( .B1(n54221), .B2(n67580), .C1(n63606), .C2(n67574), .A(
        n64576), .ZN(n64568) );
  NOR4_X1 U48834 ( .A1(n64548), .A2(n64549), .A3(n64550), .A4(n64551), .ZN(
        n64547) );
  OAI221_X1 U48835 ( .B1(n63134), .B2(n67628), .C1(n62263), .C2(n67622), .A(
        n64553), .ZN(n64550) );
  OAI221_X1 U48836 ( .B1(n62462), .B2(n67604), .C1(n63539), .C2(n67598), .A(
        n64554), .ZN(n64549) );
  OAI221_X1 U48837 ( .B1(n54220), .B2(n67580), .C1(n63605), .C2(n67574), .A(
        n64556), .ZN(n64548) );
  NOR4_X1 U48838 ( .A1(n64528), .A2(n64529), .A3(n64530), .A4(n64531), .ZN(
        n64527) );
  OAI221_X1 U48839 ( .B1(n63133), .B2(n67628), .C1(n62262), .C2(n67622), .A(
        n64533), .ZN(n64530) );
  OAI221_X1 U48840 ( .B1(n62461), .B2(n67604), .C1(n63538), .C2(n67598), .A(
        n64534), .ZN(n64529) );
  OAI221_X1 U48841 ( .B1(n54219), .B2(n67580), .C1(n63604), .C2(n67574), .A(
        n64536), .ZN(n64528) );
  NOR4_X1 U48842 ( .A1(n64508), .A2(n64509), .A3(n64510), .A4(n64511), .ZN(
        n64507) );
  OAI221_X1 U48843 ( .B1(n63132), .B2(n67628), .C1(n62261), .C2(n67622), .A(
        n64513), .ZN(n64510) );
  OAI221_X1 U48844 ( .B1(n62460), .B2(n67604), .C1(n63537), .C2(n67598), .A(
        n64514), .ZN(n64509) );
  OAI221_X1 U48845 ( .B1(n54218), .B2(n67580), .C1(n63603), .C2(n67574), .A(
        n64516), .ZN(n64508) );
  NOR4_X1 U48846 ( .A1(n64488), .A2(n64489), .A3(n64490), .A4(n64491), .ZN(
        n64487) );
  OAI221_X1 U48847 ( .B1(n63131), .B2(n67628), .C1(n62260), .C2(n67622), .A(
        n64493), .ZN(n64490) );
  OAI221_X1 U48848 ( .B1(n62459), .B2(n67604), .C1(n63536), .C2(n67598), .A(
        n64494), .ZN(n64489) );
  OAI221_X1 U48849 ( .B1(n54217), .B2(n67580), .C1(n63602), .C2(n67574), .A(
        n64496), .ZN(n64488) );
  NOR4_X1 U48850 ( .A1(n64468), .A2(n64469), .A3(n64470), .A4(n64471), .ZN(
        n64467) );
  OAI221_X1 U48851 ( .B1(n63130), .B2(n67628), .C1(n62259), .C2(n67622), .A(
        n64473), .ZN(n64470) );
  OAI221_X1 U48852 ( .B1(n62458), .B2(n67604), .C1(n63535), .C2(n67598), .A(
        n64474), .ZN(n64469) );
  OAI221_X1 U48853 ( .B1(n54216), .B2(n67580), .C1(n63601), .C2(n67574), .A(
        n64476), .ZN(n64468) );
  NOR4_X1 U48854 ( .A1(n64448), .A2(n64449), .A3(n64450), .A4(n64451), .ZN(
        n64447) );
  OAI221_X1 U48855 ( .B1(n63129), .B2(n67628), .C1(n62258), .C2(n67622), .A(
        n64453), .ZN(n64450) );
  OAI221_X1 U48856 ( .B1(n62457), .B2(n67604), .C1(n63534), .C2(n67598), .A(
        n64454), .ZN(n64449) );
  OAI221_X1 U48857 ( .B1(n54215), .B2(n67580), .C1(n63600), .C2(n67574), .A(
        n64456), .ZN(n64448) );
  NOR4_X1 U48858 ( .A1(n64428), .A2(n64429), .A3(n64430), .A4(n64431), .ZN(
        n64427) );
  OAI221_X1 U48859 ( .B1(n63128), .B2(n67628), .C1(n62257), .C2(n67622), .A(
        n64433), .ZN(n64430) );
  OAI221_X1 U48860 ( .B1(n62456), .B2(n67604), .C1(n63533), .C2(n67598), .A(
        n64434), .ZN(n64429) );
  OAI221_X1 U48861 ( .B1(n54214), .B2(n67580), .C1(n63599), .C2(n67574), .A(
        n64436), .ZN(n64428) );
  NOR4_X1 U48862 ( .A1(n64408), .A2(n64409), .A3(n64410), .A4(n64411), .ZN(
        n64407) );
  OAI221_X1 U48863 ( .B1(n63127), .B2(n67628), .C1(n62256), .C2(n67622), .A(
        n64413), .ZN(n64410) );
  OAI221_X1 U48864 ( .B1(n62455), .B2(n67604), .C1(n63532), .C2(n67598), .A(
        n64414), .ZN(n64409) );
  OAI221_X1 U48865 ( .B1(n54213), .B2(n67580), .C1(n63598), .C2(n67574), .A(
        n64416), .ZN(n64408) );
  NOR4_X1 U48866 ( .A1(n64388), .A2(n64389), .A3(n64390), .A4(n64391), .ZN(
        n64387) );
  OAI221_X1 U48867 ( .B1(n63126), .B2(n67628), .C1(n62255), .C2(n67622), .A(
        n64393), .ZN(n64390) );
  OAI221_X1 U48868 ( .B1(n62454), .B2(n67604), .C1(n63531), .C2(n67598), .A(
        n64394), .ZN(n64389) );
  OAI221_X1 U48869 ( .B1(n54212), .B2(n67580), .C1(n63597), .C2(n67574), .A(
        n64396), .ZN(n64388) );
  NOR4_X1 U48870 ( .A1(n64368), .A2(n64369), .A3(n64370), .A4(n64371), .ZN(
        n64367) );
  OAI221_X1 U48871 ( .B1(n63125), .B2(n67628), .C1(n62254), .C2(n67622), .A(
        n64373), .ZN(n64370) );
  OAI221_X1 U48872 ( .B1(n62453), .B2(n67604), .C1(n63530), .C2(n67598), .A(
        n64374), .ZN(n64369) );
  OAI221_X1 U48873 ( .B1(n54211), .B2(n67580), .C1(n63596), .C2(n67574), .A(
        n64376), .ZN(n64368) );
  NOR4_X1 U48874 ( .A1(n64348), .A2(n64349), .A3(n64350), .A4(n64351), .ZN(
        n64347) );
  OAI221_X1 U48875 ( .B1(n63124), .B2(n67629), .C1(n62253), .C2(n67623), .A(
        n64353), .ZN(n64350) );
  OAI221_X1 U48876 ( .B1(n62452), .B2(n67605), .C1(n63529), .C2(n67599), .A(
        n64354), .ZN(n64349) );
  OAI221_X1 U48877 ( .B1(n54210), .B2(n67581), .C1(n63595), .C2(n67575), .A(
        n64356), .ZN(n64348) );
  NOR4_X1 U48878 ( .A1(n64328), .A2(n64329), .A3(n64330), .A4(n64331), .ZN(
        n64327) );
  OAI221_X1 U48879 ( .B1(n63123), .B2(n67629), .C1(n62252), .C2(n67623), .A(
        n64333), .ZN(n64330) );
  OAI221_X1 U48880 ( .B1(n62451), .B2(n67605), .C1(n63528), .C2(n67599), .A(
        n64334), .ZN(n64329) );
  OAI221_X1 U48881 ( .B1(n54209), .B2(n67581), .C1(n63594), .C2(n67575), .A(
        n64336), .ZN(n64328) );
  NOR4_X1 U48882 ( .A1(n64308), .A2(n64309), .A3(n64310), .A4(n64311), .ZN(
        n64307) );
  OAI221_X1 U48883 ( .B1(n63122), .B2(n67629), .C1(n62251), .C2(n67623), .A(
        n64313), .ZN(n64310) );
  OAI221_X1 U48884 ( .B1(n62450), .B2(n67605), .C1(n63527), .C2(n67599), .A(
        n64314), .ZN(n64309) );
  OAI221_X1 U48885 ( .B1(n54208), .B2(n67581), .C1(n63593), .C2(n67575), .A(
        n64316), .ZN(n64308) );
  NOR4_X1 U48886 ( .A1(n64288), .A2(n64289), .A3(n64290), .A4(n64291), .ZN(
        n64287) );
  OAI221_X1 U48887 ( .B1(n63121), .B2(n67629), .C1(n62250), .C2(n67623), .A(
        n64293), .ZN(n64290) );
  OAI221_X1 U48888 ( .B1(n62449), .B2(n67605), .C1(n63526), .C2(n67599), .A(
        n64294), .ZN(n64289) );
  OAI221_X1 U48889 ( .B1(n54207), .B2(n67581), .C1(n63592), .C2(n67575), .A(
        n64296), .ZN(n64288) );
  NOR4_X1 U48890 ( .A1(n64268), .A2(n64269), .A3(n64270), .A4(n64271), .ZN(
        n64267) );
  OAI221_X1 U48891 ( .B1(n63120), .B2(n67629), .C1(n62249), .C2(n67623), .A(
        n64273), .ZN(n64270) );
  OAI221_X1 U48892 ( .B1(n62448), .B2(n67605), .C1(n63525), .C2(n67599), .A(
        n64274), .ZN(n64269) );
  OAI221_X1 U48893 ( .B1(n54206), .B2(n67581), .C1(n63591), .C2(n67575), .A(
        n64276), .ZN(n64268) );
  NOR4_X1 U48894 ( .A1(n64248), .A2(n64249), .A3(n64250), .A4(n64251), .ZN(
        n64247) );
  OAI221_X1 U48895 ( .B1(n63119), .B2(n67629), .C1(n62248), .C2(n67623), .A(
        n64253), .ZN(n64250) );
  OAI221_X1 U48896 ( .B1(n62447), .B2(n67605), .C1(n63524), .C2(n67599), .A(
        n64254), .ZN(n64249) );
  OAI221_X1 U48897 ( .B1(n54205), .B2(n67581), .C1(n63590), .C2(n67575), .A(
        n64256), .ZN(n64248) );
  NOR4_X1 U48898 ( .A1(n64228), .A2(n64229), .A3(n64230), .A4(n64231), .ZN(
        n64227) );
  OAI221_X1 U48899 ( .B1(n63118), .B2(n67629), .C1(n62247), .C2(n67623), .A(
        n64233), .ZN(n64230) );
  OAI221_X1 U48900 ( .B1(n62446), .B2(n67605), .C1(n63523), .C2(n67599), .A(
        n64234), .ZN(n64229) );
  OAI221_X1 U48901 ( .B1(n54204), .B2(n67581), .C1(n63589), .C2(n67575), .A(
        n64236), .ZN(n64228) );
  NOR4_X1 U48902 ( .A1(n64208), .A2(n64209), .A3(n64210), .A4(n64211), .ZN(
        n64207) );
  OAI221_X1 U48903 ( .B1(n63117), .B2(n67629), .C1(n62246), .C2(n67623), .A(
        n64213), .ZN(n64210) );
  OAI221_X1 U48904 ( .B1(n62445), .B2(n67605), .C1(n63522), .C2(n67599), .A(
        n64214), .ZN(n64209) );
  OAI221_X1 U48905 ( .B1(n54203), .B2(n67581), .C1(n63588), .C2(n67575), .A(
        n64216), .ZN(n64208) );
  NOR4_X1 U48906 ( .A1(n64188), .A2(n64189), .A3(n64190), .A4(n64191), .ZN(
        n64187) );
  OAI221_X1 U48907 ( .B1(n63116), .B2(n67629), .C1(n62245), .C2(n67623), .A(
        n64193), .ZN(n64190) );
  OAI221_X1 U48908 ( .B1(n62444), .B2(n67605), .C1(n63521), .C2(n67599), .A(
        n64194), .ZN(n64189) );
  OAI221_X1 U48909 ( .B1(n54202), .B2(n67581), .C1(n63587), .C2(n67575), .A(
        n64196), .ZN(n64188) );
  NOR4_X1 U48910 ( .A1(n64168), .A2(n64169), .A3(n64170), .A4(n64171), .ZN(
        n64167) );
  OAI221_X1 U48911 ( .B1(n63115), .B2(n67629), .C1(n62244), .C2(n67623), .A(
        n64173), .ZN(n64170) );
  OAI221_X1 U48912 ( .B1(n62443), .B2(n67605), .C1(n63520), .C2(n67599), .A(
        n64174), .ZN(n64169) );
  OAI221_X1 U48913 ( .B1(n54201), .B2(n67581), .C1(n63586), .C2(n67575), .A(
        n64176), .ZN(n64168) );
  NOR4_X1 U48914 ( .A1(n64148), .A2(n64149), .A3(n64150), .A4(n64151), .ZN(
        n64147) );
  OAI221_X1 U48915 ( .B1(n63114), .B2(n67629), .C1(n62243), .C2(n67623), .A(
        n64153), .ZN(n64150) );
  OAI221_X1 U48916 ( .B1(n62442), .B2(n67605), .C1(n63519), .C2(n67599), .A(
        n64154), .ZN(n64149) );
  OAI221_X1 U48917 ( .B1(n54200), .B2(n67581), .C1(n63585), .C2(n67575), .A(
        n64156), .ZN(n64148) );
  NOR4_X1 U48918 ( .A1(n64128), .A2(n64129), .A3(n64130), .A4(n64131), .ZN(
        n64127) );
  OAI221_X1 U48919 ( .B1(n63113), .B2(n67629), .C1(n62242), .C2(n67623), .A(
        n64133), .ZN(n64130) );
  OAI221_X1 U48920 ( .B1(n62441), .B2(n67605), .C1(n63518), .C2(n67599), .A(
        n64134), .ZN(n64129) );
  OAI221_X1 U48921 ( .B1(n54199), .B2(n67581), .C1(n63584), .C2(n67575), .A(
        n64136), .ZN(n64128) );
  NOR4_X1 U48922 ( .A1(n64108), .A2(n64109), .A3(n64110), .A4(n64111), .ZN(
        n64107) );
  OAI221_X1 U48923 ( .B1(n63112), .B2(n67630), .C1(n62241), .C2(n67624), .A(
        n64113), .ZN(n64110) );
  OAI221_X1 U48924 ( .B1(n62440), .B2(n67606), .C1(n63517), .C2(n67600), .A(
        n64114), .ZN(n64109) );
  OAI221_X1 U48925 ( .B1(n54198), .B2(n67582), .C1(n63583), .C2(n67576), .A(
        n64116), .ZN(n64108) );
  NOR4_X1 U48926 ( .A1(n64088), .A2(n64089), .A3(n64090), .A4(n64091), .ZN(
        n64087) );
  OAI221_X1 U48927 ( .B1(n63111), .B2(n67630), .C1(n62240), .C2(n67624), .A(
        n64093), .ZN(n64090) );
  OAI221_X1 U48928 ( .B1(n62439), .B2(n67606), .C1(n63516), .C2(n67600), .A(
        n64094), .ZN(n64089) );
  OAI221_X1 U48929 ( .B1(n54197), .B2(n67582), .C1(n63582), .C2(n67576), .A(
        n64096), .ZN(n64088) );
  NOR4_X1 U48930 ( .A1(n64068), .A2(n64069), .A3(n64070), .A4(n64071), .ZN(
        n64067) );
  OAI221_X1 U48931 ( .B1(n63110), .B2(n67630), .C1(n62239), .C2(n67624), .A(
        n64073), .ZN(n64070) );
  OAI221_X1 U48932 ( .B1(n62438), .B2(n67606), .C1(n63515), .C2(n67600), .A(
        n64074), .ZN(n64069) );
  OAI221_X1 U48933 ( .B1(n54196), .B2(n67582), .C1(n63581), .C2(n67576), .A(
        n64076), .ZN(n64068) );
  NOR4_X1 U48934 ( .A1(n64048), .A2(n64049), .A3(n64050), .A4(n64051), .ZN(
        n64047) );
  OAI221_X1 U48935 ( .B1(n63109), .B2(n67630), .C1(n62238), .C2(n67624), .A(
        n64053), .ZN(n64050) );
  OAI221_X1 U48936 ( .B1(n62437), .B2(n67606), .C1(n63514), .C2(n67600), .A(
        n64054), .ZN(n64049) );
  OAI221_X1 U48937 ( .B1(n54195), .B2(n67582), .C1(n63580), .C2(n67576), .A(
        n64056), .ZN(n64048) );
  NOR4_X1 U48938 ( .A1(n64028), .A2(n64029), .A3(n64030), .A4(n64031), .ZN(
        n64027) );
  OAI221_X1 U48939 ( .B1(n63108), .B2(n67630), .C1(n62237), .C2(n67624), .A(
        n64033), .ZN(n64030) );
  OAI221_X1 U48940 ( .B1(n62436), .B2(n67606), .C1(n63513), .C2(n67600), .A(
        n64034), .ZN(n64029) );
  OAI221_X1 U48941 ( .B1(n54194), .B2(n67582), .C1(n63579), .C2(n67576), .A(
        n64036), .ZN(n64028) );
  NOR4_X1 U48942 ( .A1(n64008), .A2(n64009), .A3(n64010), .A4(n64011), .ZN(
        n64007) );
  OAI221_X1 U48943 ( .B1(n63107), .B2(n67630), .C1(n62236), .C2(n67624), .A(
        n64013), .ZN(n64010) );
  OAI221_X1 U48944 ( .B1(n62435), .B2(n67606), .C1(n63512), .C2(n67600), .A(
        n64014), .ZN(n64009) );
  OAI221_X1 U48945 ( .B1(n54193), .B2(n67582), .C1(n63578), .C2(n67576), .A(
        n64016), .ZN(n64008) );
  NOR4_X1 U48946 ( .A1(n63988), .A2(n63989), .A3(n63990), .A4(n63991), .ZN(
        n63987) );
  OAI221_X1 U48947 ( .B1(n63106), .B2(n67630), .C1(n62235), .C2(n67624), .A(
        n63993), .ZN(n63990) );
  OAI221_X1 U48948 ( .B1(n62434), .B2(n67606), .C1(n63511), .C2(n67600), .A(
        n63994), .ZN(n63989) );
  OAI221_X1 U48949 ( .B1(n54192), .B2(n67582), .C1(n63577), .C2(n67576), .A(
        n63996), .ZN(n63988) );
  NOR4_X1 U48950 ( .A1(n63968), .A2(n63969), .A3(n63970), .A4(n63971), .ZN(
        n63967) );
  OAI221_X1 U48951 ( .B1(n63105), .B2(n67630), .C1(n62234), .C2(n67624), .A(
        n63973), .ZN(n63970) );
  OAI221_X1 U48952 ( .B1(n62433), .B2(n67606), .C1(n63510), .C2(n67600), .A(
        n63974), .ZN(n63969) );
  OAI221_X1 U48953 ( .B1(n54191), .B2(n67582), .C1(n63576), .C2(n67576), .A(
        n63976), .ZN(n63968) );
  NOR4_X1 U48954 ( .A1(n63948), .A2(n63949), .A3(n63950), .A4(n63951), .ZN(
        n63947) );
  OAI221_X1 U48955 ( .B1(n63104), .B2(n67630), .C1(n62233), .C2(n67624), .A(
        n63953), .ZN(n63950) );
  OAI221_X1 U48956 ( .B1(n62432), .B2(n67606), .C1(n63509), .C2(n67600), .A(
        n63954), .ZN(n63949) );
  OAI221_X1 U48957 ( .B1(n54190), .B2(n67582), .C1(n63575), .C2(n67576), .A(
        n63956), .ZN(n63948) );
  NOR4_X1 U48958 ( .A1(n63928), .A2(n63929), .A3(n63930), .A4(n63931), .ZN(
        n63927) );
  OAI221_X1 U48959 ( .B1(n63103), .B2(n67630), .C1(n62232), .C2(n67624), .A(
        n63933), .ZN(n63930) );
  OAI221_X1 U48960 ( .B1(n62431), .B2(n67606), .C1(n63508), .C2(n67600), .A(
        n63934), .ZN(n63929) );
  OAI221_X1 U48961 ( .B1(n54189), .B2(n67582), .C1(n63574), .C2(n67576), .A(
        n63936), .ZN(n63928) );
  NOR4_X1 U48962 ( .A1(n63908), .A2(n63909), .A3(n63910), .A4(n63911), .ZN(
        n63907) );
  OAI221_X1 U48963 ( .B1(n63102), .B2(n67630), .C1(n62231), .C2(n67624), .A(
        n63913), .ZN(n63910) );
  OAI221_X1 U48964 ( .B1(n62430), .B2(n67606), .C1(n63507), .C2(n67600), .A(
        n63914), .ZN(n63909) );
  OAI221_X1 U48965 ( .B1(n54188), .B2(n67582), .C1(n63573), .C2(n67576), .A(
        n63916), .ZN(n63908) );
  NOR4_X1 U48966 ( .A1(n63888), .A2(n63889), .A3(n63890), .A4(n63891), .ZN(
        n63887) );
  OAI221_X1 U48967 ( .B1(n63101), .B2(n67630), .C1(n62230), .C2(n67624), .A(
        n63893), .ZN(n63890) );
  OAI221_X1 U48968 ( .B1(n62429), .B2(n67606), .C1(n63506), .C2(n67600), .A(
        n63894), .ZN(n63889) );
  OAI221_X1 U48969 ( .B1(n54187), .B2(n67582), .C1(n63572), .C2(n67576), .A(
        n63896), .ZN(n63888) );
  NOR4_X1 U48970 ( .A1(n63877), .A2(n63878), .A3(n63879), .A4(n63880), .ZN(
        n63865) );
  OAI222_X1 U48971 ( .A1(n63166), .A2(n67523), .B1(n62095), .B2(n67517), .C1(
        n62498), .C2(n67511), .ZN(n63877) );
  OAI22_X1 U48972 ( .A1(n8449), .A2(n67547), .B1(n62362), .B2(n67541), .ZN(
        n63879) );
  OAI22_X1 U48973 ( .A1(n62631), .A2(n67559), .B1(n54610), .B2(n67553), .ZN(
        n63880) );
  NOR4_X1 U48974 ( .A1(n63856), .A2(n63857), .A3(n63858), .A4(n63859), .ZN(
        n63844) );
  OAI222_X1 U48975 ( .A1(n63165), .A2(n67523), .B1(n62094), .B2(n67517), .C1(
        n62497), .C2(n67511), .ZN(n63856) );
  OAI22_X1 U48976 ( .A1(n8465), .A2(n67547), .B1(n62361), .B2(n67541), .ZN(
        n63858) );
  OAI22_X1 U48977 ( .A1(n62630), .A2(n67559), .B1(n54609), .B2(n67553), .ZN(
        n63859) );
  NOR4_X1 U48978 ( .A1(n63835), .A2(n63836), .A3(n63837), .A4(n63838), .ZN(
        n63823) );
  OAI222_X1 U48979 ( .A1(n63164), .A2(n67523), .B1(n62093), .B2(n67517), .C1(
        n62496), .C2(n67511), .ZN(n63835) );
  OAI22_X1 U48980 ( .A1(n8481), .A2(n67547), .B1(n62360), .B2(n67541), .ZN(
        n63837) );
  OAI22_X1 U48981 ( .A1(n62629), .A2(n67559), .B1(n54608), .B2(n67553), .ZN(
        n63838) );
  NOR4_X1 U48982 ( .A1(n63797), .A2(n63798), .A3(n63799), .A4(n63800), .ZN(
        n63769) );
  OAI222_X1 U48983 ( .A1(n63162), .A2(n67523), .B1(n62091), .B2(n67517), .C1(
        n62494), .C2(n67511), .ZN(n63797) );
  OAI22_X1 U48984 ( .A1(n8497), .A2(n67547), .B1(n62358), .B2(n67541), .ZN(
        n63799) );
  OAI22_X1 U48985 ( .A1(n62627), .A2(n67559), .B1(n54606), .B2(n67553), .ZN(
        n63800) );
  AOI221_X1 U48986 ( .B1(n67307), .B2(n58717), .C1(n67301), .C2(n58299), .A(
        n65167), .ZN(n65152) );
  OAI22_X1 U48987 ( .A1(n62093), .A2(n67295), .B1(n62160), .B2(n67289), .ZN(
        n65167) );
  AOI221_X1 U48988 ( .B1(n67307), .B2(n58718), .C1(n67301), .C2(n58301), .A(
        n65143), .ZN(n65101) );
  OAI22_X1 U48989 ( .A1(n62091), .A2(n67295), .B1(n62158), .B2(n67289), .ZN(
        n65143) );
  AOI221_X1 U48990 ( .B1(n67307), .B2(n58715), .C1(n67301), .C2(n58295), .A(
        n65203), .ZN(n65188) );
  OAI22_X1 U48991 ( .A1(n62095), .A2(n67295), .B1(n62162), .B2(n67289), .ZN(
        n65203) );
  AOI221_X1 U48992 ( .B1(n67307), .B2(n58716), .C1(n67301), .C2(n58297), .A(
        n65185), .ZN(n65170) );
  OAI22_X1 U48993 ( .A1(n62094), .A2(n67295), .B1(n62161), .B2(n67289), .ZN(
        n65185) );
  NAND2_X1 U48994 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .ZN(n62489) );
  NAND2_X1 U48995 ( .A1(ADD_WR[2]), .A2(n63497), .ZN(n62356) );
  NAND2_X1 U48996 ( .A1(ADD_WR[1]), .A2(n63496), .ZN(n62223) );
  AND3_X1 U48997 ( .A1(n66494), .A2(n65099), .A3(ADD_RD1[1]), .ZN(n65075) );
  OAI221_X1 U48998 ( .B1(n63415), .B2(n67649), .C1(n49432), .C2(n67643), .A(
        n64832), .ZN(n64831) );
  AOI22_X1 U48999 ( .A1(n67637), .A2(n57725), .B1(n67633), .B2(OUT1[12]), .ZN(
        n64832) );
  OAI221_X1 U49000 ( .B1(n63414), .B2(n67649), .C1(n49433), .C2(n67643), .A(
        n64812), .ZN(n64811) );
  AOI22_X1 U49001 ( .A1(n67637), .A2(n57701), .B1(n67635), .B2(OUT1[13]), .ZN(
        n64812) );
  OAI221_X1 U49002 ( .B1(n63413), .B2(n67649), .C1(n49434), .C2(n67643), .A(
        n64792), .ZN(n64791) );
  AOI22_X1 U49003 ( .A1(n67637), .A2(n57677), .B1(n67634), .B2(OUT1[14]), .ZN(
        n64792) );
  OAI221_X1 U49004 ( .B1(n63412), .B2(n67649), .C1(n49435), .C2(n67643), .A(
        n64772), .ZN(n64771) );
  AOI22_X1 U49005 ( .A1(n67637), .A2(n57653), .B1(n67633), .B2(OUT1[15]), .ZN(
        n64772) );
  OAI221_X1 U49006 ( .B1(n63411), .B2(n67649), .C1(n49436), .C2(n67643), .A(
        n64752), .ZN(n64751) );
  AOI22_X1 U49007 ( .A1(n67637), .A2(n57629), .B1(n67635), .B2(OUT1[16]), .ZN(
        n64752) );
  OAI221_X1 U49008 ( .B1(n63410), .B2(n67649), .C1(n49437), .C2(n67643), .A(
        n64732), .ZN(n64731) );
  AOI22_X1 U49009 ( .A1(n67637), .A2(n57605), .B1(n67634), .B2(OUT1[17]), .ZN(
        n64732) );
  OAI221_X1 U49010 ( .B1(n63409), .B2(n67649), .C1(n49438), .C2(n67643), .A(
        n64712), .ZN(n64711) );
  AOI22_X1 U49011 ( .A1(n67637), .A2(n57581), .B1(n67633), .B2(OUT1[18]), .ZN(
        n64712) );
  OAI221_X1 U49012 ( .B1(n63408), .B2(n67649), .C1(n49439), .C2(n67643), .A(
        n64692), .ZN(n64691) );
  AOI22_X1 U49013 ( .A1(n67637), .A2(n57557), .B1(n67635), .B2(OUT1[19]), .ZN(
        n64692) );
  OAI221_X1 U49014 ( .B1(n63407), .B2(n67649), .C1(n49440), .C2(n67643), .A(
        n64672), .ZN(n64671) );
  AOI22_X1 U49015 ( .A1(n67637), .A2(n57533), .B1(n67634), .B2(OUT1[20]), .ZN(
        n64672) );
  OAI221_X1 U49016 ( .B1(n63406), .B2(n67649), .C1(n49441), .C2(n67643), .A(
        n64652), .ZN(n64651) );
  AOI22_X1 U49017 ( .A1(n67637), .A2(n57509), .B1(n67633), .B2(OUT1[21]), .ZN(
        n64652) );
  OAI221_X1 U49018 ( .B1(n63405), .B2(n67649), .C1(n49442), .C2(n67643), .A(
        n64632), .ZN(n64631) );
  AOI22_X1 U49019 ( .A1(n67637), .A2(n57485), .B1(n67634), .B2(OUT1[22]), .ZN(
        n64632) );
  OAI221_X1 U49020 ( .B1(n63404), .B2(n67649), .C1(n49443), .C2(n67643), .A(
        n64612), .ZN(n64611) );
  AOI22_X1 U49021 ( .A1(n67637), .A2(n57461), .B1(n67633), .B2(OUT1[23]), .ZN(
        n64612) );
  OAI221_X1 U49022 ( .B1(n63403), .B2(n67650), .C1(n49444), .C2(n67644), .A(
        n64592), .ZN(n64591) );
  AOI22_X1 U49023 ( .A1(n67638), .A2(n57437), .B1(n67633), .B2(OUT1[24]), .ZN(
        n64592) );
  OAI221_X1 U49024 ( .B1(n63402), .B2(n67650), .C1(n49445), .C2(n67644), .A(
        n64572), .ZN(n64571) );
  AOI22_X1 U49025 ( .A1(n67638), .A2(n57413), .B1(n67633), .B2(OUT1[25]), .ZN(
        n64572) );
  OAI221_X1 U49026 ( .B1(n63401), .B2(n67650), .C1(n49446), .C2(n67644), .A(
        n64552), .ZN(n64551) );
  AOI22_X1 U49027 ( .A1(n67638), .A2(n57389), .B1(n67633), .B2(OUT1[26]), .ZN(
        n64552) );
  OAI221_X1 U49028 ( .B1(n63400), .B2(n67650), .C1(n49447), .C2(n67644), .A(
        n64532), .ZN(n64531) );
  AOI22_X1 U49029 ( .A1(n67638), .A2(n57365), .B1(n67633), .B2(OUT1[27]), .ZN(
        n64532) );
  OAI221_X1 U49030 ( .B1(n63399), .B2(n67650), .C1(n49448), .C2(n67644), .A(
        n64512), .ZN(n64511) );
  AOI22_X1 U49031 ( .A1(n67638), .A2(n57341), .B1(n67633), .B2(OUT1[28]), .ZN(
        n64512) );
  OAI221_X1 U49032 ( .B1(n63398), .B2(n67650), .C1(n49449), .C2(n67644), .A(
        n64492), .ZN(n64491) );
  AOI22_X1 U49033 ( .A1(n67638), .A2(n57317), .B1(n67633), .B2(OUT1[29]), .ZN(
        n64492) );
  OAI221_X1 U49034 ( .B1(n63397), .B2(n67650), .C1(n49450), .C2(n67644), .A(
        n64472), .ZN(n64471) );
  AOI22_X1 U49035 ( .A1(n67638), .A2(n57293), .B1(n67633), .B2(OUT1[30]), .ZN(
        n64472) );
  OAI221_X1 U49036 ( .B1(n63396), .B2(n67650), .C1(n49451), .C2(n67644), .A(
        n64452), .ZN(n64451) );
  AOI22_X1 U49037 ( .A1(n67638), .A2(n57269), .B1(n67633), .B2(OUT1[31]), .ZN(
        n64452) );
  OAI221_X1 U49038 ( .B1(n63395), .B2(n67650), .C1(n49452), .C2(n67644), .A(
        n64432), .ZN(n64431) );
  AOI22_X1 U49039 ( .A1(n67638), .A2(n57245), .B1(n67633), .B2(OUT1[32]), .ZN(
        n64432) );
  OAI221_X1 U49040 ( .B1(n63394), .B2(n67650), .C1(n49453), .C2(n67644), .A(
        n64412), .ZN(n64411) );
  AOI22_X1 U49041 ( .A1(n67638), .A2(n57221), .B1(n67633), .B2(OUT1[33]), .ZN(
        n64412) );
  OAI221_X1 U49042 ( .B1(n63393), .B2(n67650), .C1(n49454), .C2(n67644), .A(
        n64392), .ZN(n64391) );
  AOI22_X1 U49043 ( .A1(n67638), .A2(n57197), .B1(n67633), .B2(OUT1[34]), .ZN(
        n64392) );
  OAI221_X1 U49044 ( .B1(n63392), .B2(n67650), .C1(n49455), .C2(n67644), .A(
        n64372), .ZN(n64371) );
  AOI22_X1 U49045 ( .A1(n67638), .A2(n57173), .B1(n67633), .B2(OUT1[35]), .ZN(
        n64372) );
  OAI221_X1 U49046 ( .B1(n63391), .B2(n67651), .C1(n49456), .C2(n67645), .A(
        n64352), .ZN(n64351) );
  AOI22_X1 U49047 ( .A1(n67639), .A2(n57149), .B1(n67633), .B2(OUT1[36]), .ZN(
        n64352) );
  OAI221_X1 U49048 ( .B1(n63390), .B2(n67651), .C1(n49457), .C2(n67645), .A(
        n64332), .ZN(n64331) );
  AOI22_X1 U49049 ( .A1(n67639), .A2(n57125), .B1(n67634), .B2(OUT1[37]), .ZN(
        n64332) );
  OAI221_X1 U49050 ( .B1(n63389), .B2(n67651), .C1(n49458), .C2(n67645), .A(
        n64312), .ZN(n64311) );
  AOI22_X1 U49051 ( .A1(n67639), .A2(n57101), .B1(n67634), .B2(OUT1[38]), .ZN(
        n64312) );
  OAI221_X1 U49052 ( .B1(n63388), .B2(n67651), .C1(n49459), .C2(n67645), .A(
        n64292), .ZN(n64291) );
  AOI22_X1 U49053 ( .A1(n67639), .A2(n57077), .B1(n67634), .B2(OUT1[39]), .ZN(
        n64292) );
  OAI221_X1 U49054 ( .B1(n63387), .B2(n67651), .C1(n49460), .C2(n67645), .A(
        n64272), .ZN(n64271) );
  AOI22_X1 U49055 ( .A1(n67639), .A2(n57053), .B1(n67634), .B2(OUT1[40]), .ZN(
        n64272) );
  OAI221_X1 U49056 ( .B1(n63386), .B2(n67651), .C1(n49461), .C2(n67645), .A(
        n64252), .ZN(n64251) );
  AOI22_X1 U49057 ( .A1(n67639), .A2(n57029), .B1(n67634), .B2(OUT1[41]), .ZN(
        n64252) );
  OAI221_X1 U49058 ( .B1(n63385), .B2(n67651), .C1(n49462), .C2(n67645), .A(
        n64232), .ZN(n64231) );
  AOI22_X1 U49059 ( .A1(n67639), .A2(n57005), .B1(n67634), .B2(OUT1[42]), .ZN(
        n64232) );
  OAI221_X1 U49060 ( .B1(n63384), .B2(n67651), .C1(n49463), .C2(n67645), .A(
        n64212), .ZN(n64211) );
  AOI22_X1 U49061 ( .A1(n67639), .A2(n56981), .B1(n67634), .B2(OUT1[43]), .ZN(
        n64212) );
  OAI221_X1 U49062 ( .B1(n63383), .B2(n67651), .C1(n49464), .C2(n67645), .A(
        n64192), .ZN(n64191) );
  AOI22_X1 U49063 ( .A1(n67639), .A2(n56957), .B1(n67634), .B2(OUT1[44]), .ZN(
        n64192) );
  OAI221_X1 U49064 ( .B1(n63382), .B2(n67651), .C1(n49465), .C2(n67645), .A(
        n64172), .ZN(n64171) );
  AOI22_X1 U49065 ( .A1(n67639), .A2(n56933), .B1(n67634), .B2(OUT1[45]), .ZN(
        n64172) );
  OAI221_X1 U49066 ( .B1(n63381), .B2(n67651), .C1(n49466), .C2(n67645), .A(
        n64152), .ZN(n64151) );
  AOI22_X1 U49067 ( .A1(n67639), .A2(n56909), .B1(n67634), .B2(OUT1[46]), .ZN(
        n64152) );
  OAI221_X1 U49068 ( .B1(n63380), .B2(n67651), .C1(n49467), .C2(n67645), .A(
        n64132), .ZN(n64131) );
  AOI22_X1 U49069 ( .A1(n67639), .A2(n56885), .B1(n67634), .B2(OUT1[47]), .ZN(
        n64132) );
  OAI221_X1 U49070 ( .B1(n63379), .B2(n67652), .C1(n49468), .C2(n67646), .A(
        n64112), .ZN(n64111) );
  AOI22_X1 U49071 ( .A1(n67640), .A2(n56861), .B1(n67634), .B2(OUT1[48]), .ZN(
        n64112) );
  OAI221_X1 U49072 ( .B1(n63378), .B2(n67652), .C1(n49469), .C2(n67646), .A(
        n64092), .ZN(n64091) );
  AOI22_X1 U49073 ( .A1(n67640), .A2(n56837), .B1(n67634), .B2(OUT1[49]), .ZN(
        n64092) );
  OAI221_X1 U49074 ( .B1(n63377), .B2(n67652), .C1(n49470), .C2(n67646), .A(
        n64072), .ZN(n64071) );
  AOI22_X1 U49075 ( .A1(n67640), .A2(n56813), .B1(n67635), .B2(OUT1[50]), .ZN(
        n64072) );
  OAI221_X1 U49076 ( .B1(n63376), .B2(n67652), .C1(n49471), .C2(n67646), .A(
        n64052), .ZN(n64051) );
  AOI22_X1 U49077 ( .A1(n67640), .A2(n56789), .B1(n67635), .B2(OUT1[51]), .ZN(
        n64052) );
  OAI221_X1 U49078 ( .B1(n63375), .B2(n67652), .C1(n49472), .C2(n67646), .A(
        n64032), .ZN(n64031) );
  AOI22_X1 U49079 ( .A1(n67640), .A2(n56765), .B1(n67635), .B2(OUT1[52]), .ZN(
        n64032) );
  OAI221_X1 U49080 ( .B1(n63374), .B2(n67652), .C1(n49473), .C2(n67646), .A(
        n64012), .ZN(n64011) );
  AOI22_X1 U49081 ( .A1(n67640), .A2(n56741), .B1(n67635), .B2(OUT1[53]), .ZN(
        n64012) );
  OAI221_X1 U49082 ( .B1(n63373), .B2(n67652), .C1(n49474), .C2(n67646), .A(
        n63992), .ZN(n63991) );
  AOI22_X1 U49083 ( .A1(n67640), .A2(n56717), .B1(n67635), .B2(OUT1[54]), .ZN(
        n63992) );
  OAI221_X1 U49084 ( .B1(n63372), .B2(n67652), .C1(n49475), .C2(n67646), .A(
        n63972), .ZN(n63971) );
  AOI22_X1 U49085 ( .A1(n67640), .A2(n56693), .B1(n67635), .B2(OUT1[55]), .ZN(
        n63972) );
  OAI221_X1 U49086 ( .B1(n63371), .B2(n67652), .C1(n49476), .C2(n67646), .A(
        n63952), .ZN(n63951) );
  AOI22_X1 U49087 ( .A1(n67640), .A2(n56669), .B1(n67635), .B2(OUT1[56]), .ZN(
        n63952) );
  OAI221_X1 U49088 ( .B1(n63370), .B2(n67652), .C1(n49477), .C2(n67646), .A(
        n63932), .ZN(n63931) );
  AOI22_X1 U49089 ( .A1(n67640), .A2(n56645), .B1(n67635), .B2(OUT1[57]), .ZN(
        n63932) );
  OAI221_X1 U49090 ( .B1(n63369), .B2(n67652), .C1(n49478), .C2(n67646), .A(
        n63912), .ZN(n63911) );
  AOI22_X1 U49091 ( .A1(n67640), .A2(n56621), .B1(n67635), .B2(OUT1[58]), .ZN(
        n63912) );
  OAI221_X1 U49092 ( .B1(n63368), .B2(n67652), .C1(n49479), .C2(n67646), .A(
        n63892), .ZN(n63891) );
  AOI22_X1 U49093 ( .A1(n67640), .A2(n56597), .B1(n67635), .B2(OUT1[59]), .ZN(
        n63892) );
  OAI221_X1 U49094 ( .B1(n63365), .B2(n67457), .C1(n49231), .C2(n67451), .A(
        n65159), .ZN(n65158) );
  AOI22_X1 U49095 ( .A1(n67445), .A2(n58377), .B1(n67439), .B2(OUT2[62]), .ZN(
        n65159) );
  OAI221_X1 U49096 ( .B1(n63363), .B2(n67457), .C1(n49228), .C2(n67451), .A(
        n65110), .ZN(n65107) );
  AOI22_X1 U49097 ( .A1(n67445), .A2(n58378), .B1(n67439), .B2(OUT2[63]), .ZN(
        n65110) );
  OAI221_X1 U49098 ( .B1(n63367), .B2(n67457), .C1(n49229), .C2(n67451), .A(
        n65195), .ZN(n65194) );
  AOI22_X1 U49099 ( .A1(n67445), .A2(n58375), .B1(n67438), .B2(OUT2[60]), .ZN(
        n65195) );
  OAI221_X1 U49100 ( .B1(n63366), .B2(n67457), .C1(n49230), .C2(n67451), .A(
        n65177), .ZN(n65176) );
  AOI22_X1 U49101 ( .A1(n67445), .A2(n58376), .B1(n67439), .B2(OUT2[61]), .ZN(
        n65177) );
  OAI221_X1 U49102 ( .B1(n63367), .B2(n67653), .C1(n49480), .C2(n67647), .A(
        n63871), .ZN(n63870) );
  AOI22_X1 U49103 ( .A1(n67641), .A2(n58784), .B1(n67635), .B2(OUT1[60]), .ZN(
        n63871) );
  OAI221_X1 U49104 ( .B1(n63366), .B2(n67653), .C1(n49481), .C2(n67647), .A(
        n63850), .ZN(n63849) );
  AOI22_X1 U49105 ( .A1(n67641), .A2(n58785), .B1(n67635), .B2(OUT1[61]), .ZN(
        n63850) );
  OAI221_X1 U49106 ( .B1(n63365), .B2(n67653), .C1(n49482), .C2(n67647), .A(
        n63829), .ZN(n63828) );
  AOI22_X1 U49107 ( .A1(n67641), .A2(n58786), .B1(n67635), .B2(OUT1[62]), .ZN(
        n63829) );
  OAI221_X1 U49108 ( .B1(n63363), .B2(n67653), .C1(n49483), .C2(n67647), .A(
        n63777), .ZN(n63774) );
  AOI22_X1 U49109 ( .A1(n67641), .A2(n58783), .B1(n67635), .B2(OUT1[63]), .ZN(
        n63777) );
  OAI221_X1 U49110 ( .B1(n54658), .B2(n67429), .C1(n63553), .C2(n67423), .A(
        n66060), .ZN(n66057) );
  AOI22_X1 U49111 ( .A1(n67417), .A2(n66325), .B1(n67411), .B2(n58319), .ZN(
        n66060) );
  OAI221_X1 U49112 ( .B1(n54657), .B2(n67429), .C1(n63552), .C2(n67423), .A(
        n66042), .ZN(n66039) );
  AOI22_X1 U49113 ( .A1(n67417), .A2(n66326), .B1(n67411), .B2(n58320), .ZN(
        n66042) );
  OAI221_X1 U49114 ( .B1(n54656), .B2(n67429), .C1(n63551), .C2(n67423), .A(
        n66024), .ZN(n66021) );
  AOI22_X1 U49115 ( .A1(n67417), .A2(n66327), .B1(n67411), .B2(n58321), .ZN(
        n66024) );
  OAI221_X1 U49116 ( .B1(n54655), .B2(n67429), .C1(n63550), .C2(n67423), .A(
        n66006), .ZN(n66003) );
  AOI22_X1 U49117 ( .A1(n67417), .A2(n66328), .B1(n67411), .B2(n58322), .ZN(
        n66006) );
  OAI221_X1 U49118 ( .B1(n54654), .B2(n67429), .C1(n63549), .C2(n67423), .A(
        n65988), .ZN(n65985) );
  AOI22_X1 U49119 ( .A1(n67417), .A2(n66329), .B1(n67411), .B2(n58323), .ZN(
        n65988) );
  OAI221_X1 U49120 ( .B1(n54653), .B2(n67429), .C1(n63548), .C2(n67423), .A(
        n65970), .ZN(n65967) );
  AOI22_X1 U49121 ( .A1(n67417), .A2(n66330), .B1(n67411), .B2(n58324), .ZN(
        n65970) );
  OAI221_X1 U49122 ( .B1(n54652), .B2(n67429), .C1(n63547), .C2(n67423), .A(
        n65952), .ZN(n65949) );
  AOI22_X1 U49123 ( .A1(n67417), .A2(n66331), .B1(n67411), .B2(n58325), .ZN(
        n65952) );
  OAI221_X1 U49124 ( .B1(n54651), .B2(n67429), .C1(n63546), .C2(n67423), .A(
        n65934), .ZN(n65931) );
  AOI22_X1 U49125 ( .A1(n67417), .A2(n66332), .B1(n67411), .B2(n58326), .ZN(
        n65934) );
  OAI221_X1 U49126 ( .B1(n54650), .B2(n67429), .C1(n63545), .C2(n67423), .A(
        n65916), .ZN(n65913) );
  AOI22_X1 U49127 ( .A1(n67417), .A2(n66333), .B1(n67411), .B2(n58327), .ZN(
        n65916) );
  OAI221_X1 U49128 ( .B1(n54649), .B2(n67429), .C1(n63544), .C2(n67423), .A(
        n65898), .ZN(n65895) );
  AOI22_X1 U49129 ( .A1(n67417), .A2(n66334), .B1(n67411), .B2(n58328), .ZN(
        n65898) );
  OAI221_X1 U49130 ( .B1(n54648), .B2(n67429), .C1(n63543), .C2(n67423), .A(
        n65880), .ZN(n65877) );
  AOI22_X1 U49131 ( .A1(n67417), .A2(n66335), .B1(n67411), .B2(n58329), .ZN(
        n65880) );
  OAI221_X1 U49132 ( .B1(n54647), .B2(n67429), .C1(n63542), .C2(n67423), .A(
        n65862), .ZN(n65859) );
  AOI22_X1 U49133 ( .A1(n67417), .A2(n66336), .B1(n67411), .B2(n58330), .ZN(
        n65862) );
  OAI221_X1 U49134 ( .B1(n54646), .B2(n67430), .C1(n63541), .C2(n67424), .A(
        n65844), .ZN(n65841) );
  AOI22_X1 U49135 ( .A1(n67418), .A2(n66337), .B1(n67412), .B2(n58331), .ZN(
        n65844) );
  OAI221_X1 U49136 ( .B1(n54645), .B2(n67430), .C1(n63540), .C2(n67424), .A(
        n65826), .ZN(n65823) );
  AOI22_X1 U49137 ( .A1(n67418), .A2(n66338), .B1(n67412), .B2(n58332), .ZN(
        n65826) );
  OAI221_X1 U49138 ( .B1(n54644), .B2(n67430), .C1(n63539), .C2(n67424), .A(
        n65808), .ZN(n65805) );
  AOI22_X1 U49139 ( .A1(n67418), .A2(n66339), .B1(n67412), .B2(n58333), .ZN(
        n65808) );
  OAI221_X1 U49140 ( .B1(n54643), .B2(n67430), .C1(n63538), .C2(n67424), .A(
        n65790), .ZN(n65787) );
  AOI22_X1 U49141 ( .A1(n67418), .A2(n66340), .B1(n67412), .B2(n58334), .ZN(
        n65790) );
  OAI221_X1 U49142 ( .B1(n54642), .B2(n67430), .C1(n63537), .C2(n67424), .A(
        n65772), .ZN(n65769) );
  AOI22_X1 U49143 ( .A1(n67418), .A2(n66341), .B1(n67412), .B2(n58335), .ZN(
        n65772) );
  OAI221_X1 U49144 ( .B1(n54641), .B2(n67430), .C1(n63536), .C2(n67424), .A(
        n65754), .ZN(n65751) );
  AOI22_X1 U49145 ( .A1(n67418), .A2(n66342), .B1(n67412), .B2(n58336), .ZN(
        n65754) );
  OAI221_X1 U49146 ( .B1(n54640), .B2(n67430), .C1(n63535), .C2(n67424), .A(
        n65736), .ZN(n65733) );
  AOI22_X1 U49147 ( .A1(n67418), .A2(n66343), .B1(n67412), .B2(n58337), .ZN(
        n65736) );
  OAI221_X1 U49148 ( .B1(n54639), .B2(n67430), .C1(n63534), .C2(n67424), .A(
        n65718), .ZN(n65715) );
  AOI22_X1 U49149 ( .A1(n67418), .A2(n66344), .B1(n67412), .B2(n58338), .ZN(
        n65718) );
  OAI221_X1 U49150 ( .B1(n54638), .B2(n67430), .C1(n63533), .C2(n67424), .A(
        n65700), .ZN(n65697) );
  AOI22_X1 U49151 ( .A1(n67418), .A2(n66345), .B1(n67412), .B2(n58339), .ZN(
        n65700) );
  OAI221_X1 U49152 ( .B1(n54637), .B2(n67430), .C1(n63532), .C2(n67424), .A(
        n65682), .ZN(n65679) );
  AOI22_X1 U49153 ( .A1(n67418), .A2(n66346), .B1(n67412), .B2(n58340), .ZN(
        n65682) );
  OAI221_X1 U49154 ( .B1(n54636), .B2(n67430), .C1(n63531), .C2(n67424), .A(
        n65664), .ZN(n65661) );
  AOI22_X1 U49155 ( .A1(n67418), .A2(n66347), .B1(n67412), .B2(n58341), .ZN(
        n65664) );
  OAI221_X1 U49156 ( .B1(n54635), .B2(n67430), .C1(n63530), .C2(n67424), .A(
        n65646), .ZN(n65643) );
  AOI22_X1 U49157 ( .A1(n67418), .A2(n66348), .B1(n67412), .B2(n58342), .ZN(
        n65646) );
  OAI221_X1 U49158 ( .B1(n54634), .B2(n67431), .C1(n63529), .C2(n67425), .A(
        n65628), .ZN(n65625) );
  AOI22_X1 U49159 ( .A1(n67419), .A2(n66349), .B1(n67413), .B2(n58343), .ZN(
        n65628) );
  OAI221_X1 U49160 ( .B1(n54633), .B2(n67431), .C1(n63528), .C2(n67425), .A(
        n65610), .ZN(n65607) );
  AOI22_X1 U49161 ( .A1(n67419), .A2(n66350), .B1(n67413), .B2(n58344), .ZN(
        n65610) );
  OAI221_X1 U49162 ( .B1(n54632), .B2(n67431), .C1(n63527), .C2(n67425), .A(
        n65592), .ZN(n65589) );
  AOI22_X1 U49163 ( .A1(n67419), .A2(n66351), .B1(n67413), .B2(n58345), .ZN(
        n65592) );
  OAI221_X1 U49164 ( .B1(n54631), .B2(n67431), .C1(n63526), .C2(n67425), .A(
        n65574), .ZN(n65571) );
  AOI22_X1 U49165 ( .A1(n67419), .A2(n66352), .B1(n67413), .B2(n58346), .ZN(
        n65574) );
  OAI221_X1 U49166 ( .B1(n54630), .B2(n67431), .C1(n63525), .C2(n67425), .A(
        n65556), .ZN(n65553) );
  AOI22_X1 U49167 ( .A1(n67419), .A2(n66353), .B1(n67413), .B2(n58347), .ZN(
        n65556) );
  OAI221_X1 U49168 ( .B1(n54629), .B2(n67431), .C1(n63524), .C2(n67425), .A(
        n65538), .ZN(n65535) );
  AOI22_X1 U49169 ( .A1(n67419), .A2(n66354), .B1(n67413), .B2(n58348), .ZN(
        n65538) );
  OAI221_X1 U49170 ( .B1(n54628), .B2(n67431), .C1(n63523), .C2(n67425), .A(
        n65520), .ZN(n65517) );
  AOI22_X1 U49171 ( .A1(n67419), .A2(n66355), .B1(n67413), .B2(n58349), .ZN(
        n65520) );
  OAI221_X1 U49172 ( .B1(n54627), .B2(n67431), .C1(n63522), .C2(n67425), .A(
        n65502), .ZN(n65499) );
  AOI22_X1 U49173 ( .A1(n67419), .A2(n66356), .B1(n67413), .B2(n58350), .ZN(
        n65502) );
  OAI221_X1 U49174 ( .B1(n54626), .B2(n67431), .C1(n63521), .C2(n67425), .A(
        n65484), .ZN(n65481) );
  AOI22_X1 U49175 ( .A1(n67419), .A2(n66357), .B1(n67413), .B2(n58351), .ZN(
        n65484) );
  OAI221_X1 U49176 ( .B1(n54625), .B2(n67431), .C1(n63520), .C2(n67425), .A(
        n65466), .ZN(n65463) );
  AOI22_X1 U49177 ( .A1(n67419), .A2(n66358), .B1(n67413), .B2(n58352), .ZN(
        n65466) );
  OAI221_X1 U49178 ( .B1(n54624), .B2(n67431), .C1(n63519), .C2(n67425), .A(
        n65448), .ZN(n65445) );
  AOI22_X1 U49179 ( .A1(n67419), .A2(n66359), .B1(n67413), .B2(n58353), .ZN(
        n65448) );
  OAI221_X1 U49180 ( .B1(n54623), .B2(n67431), .C1(n63518), .C2(n67425), .A(
        n65430), .ZN(n65427) );
  AOI22_X1 U49181 ( .A1(n67419), .A2(n66360), .B1(n67413), .B2(n58354), .ZN(
        n65430) );
  OAI221_X1 U49182 ( .B1(n54622), .B2(n67432), .C1(n63517), .C2(n67426), .A(
        n65412), .ZN(n65409) );
  AOI22_X1 U49183 ( .A1(n67420), .A2(n66361), .B1(n67414), .B2(n58355), .ZN(
        n65412) );
  OAI221_X1 U49184 ( .B1(n54621), .B2(n67432), .C1(n63516), .C2(n67426), .A(
        n65394), .ZN(n65391) );
  AOI22_X1 U49185 ( .A1(n67420), .A2(n66362), .B1(n67414), .B2(n58356), .ZN(
        n65394) );
  OAI221_X1 U49186 ( .B1(n54620), .B2(n67432), .C1(n63515), .C2(n67426), .A(
        n65376), .ZN(n65373) );
  AOI22_X1 U49187 ( .A1(n67420), .A2(n66363), .B1(n67414), .B2(n58357), .ZN(
        n65376) );
  OAI221_X1 U49188 ( .B1(n54619), .B2(n67432), .C1(n63514), .C2(n67426), .A(
        n65358), .ZN(n65355) );
  AOI22_X1 U49189 ( .A1(n67420), .A2(n66364), .B1(n67414), .B2(n58358), .ZN(
        n65358) );
  OAI221_X1 U49190 ( .B1(n54618), .B2(n67432), .C1(n63513), .C2(n67426), .A(
        n65340), .ZN(n65337) );
  AOI22_X1 U49191 ( .A1(n67420), .A2(n66365), .B1(n67414), .B2(n58359), .ZN(
        n65340) );
  OAI221_X1 U49192 ( .B1(n54617), .B2(n67432), .C1(n63512), .C2(n67426), .A(
        n65322), .ZN(n65319) );
  AOI22_X1 U49193 ( .A1(n67420), .A2(n66366), .B1(n67414), .B2(n58360), .ZN(
        n65322) );
  OAI221_X1 U49194 ( .B1(n54616), .B2(n67432), .C1(n63511), .C2(n67426), .A(
        n65304), .ZN(n65301) );
  AOI22_X1 U49195 ( .A1(n67420), .A2(n66367), .B1(n67414), .B2(n58361), .ZN(
        n65304) );
  OAI221_X1 U49196 ( .B1(n54615), .B2(n67432), .C1(n63510), .C2(n67426), .A(
        n65286), .ZN(n65283) );
  AOI22_X1 U49197 ( .A1(n67420), .A2(n66368), .B1(n67414), .B2(n58362), .ZN(
        n65286) );
  OAI221_X1 U49198 ( .B1(n54614), .B2(n67432), .C1(n63509), .C2(n67426), .A(
        n65268), .ZN(n65265) );
  AOI22_X1 U49199 ( .A1(n67420), .A2(n66369), .B1(n67414), .B2(n58363), .ZN(
        n65268) );
  OAI221_X1 U49200 ( .B1(n54613), .B2(n67432), .C1(n63508), .C2(n67426), .A(
        n65250), .ZN(n65247) );
  AOI22_X1 U49201 ( .A1(n67420), .A2(n66370), .B1(n67414), .B2(n58364), .ZN(
        n65250) );
  OAI221_X1 U49202 ( .B1(n54612), .B2(n67432), .C1(n63507), .C2(n67426), .A(
        n65232), .ZN(n65229) );
  AOI22_X1 U49203 ( .A1(n67420), .A2(n66371), .B1(n67414), .B2(n58365), .ZN(
        n65232) );
  OAI221_X1 U49204 ( .B1(n54611), .B2(n67432), .C1(n63506), .C2(n67426), .A(
        n65214), .ZN(n65211) );
  AOI22_X1 U49205 ( .A1(n67420), .A2(n66372), .B1(n67414), .B2(n58366), .ZN(
        n65214) );
  OAI221_X1 U49206 ( .B1(n54608), .B2(n67433), .C1(n63503), .C2(n67427), .A(
        n65160), .ZN(n65157) );
  AOI22_X1 U49207 ( .A1(n67421), .A2(n66307), .B1(n67415), .B2(n58306), .ZN(
        n65160) );
  OAI221_X1 U49208 ( .B1(n54606), .B2(n67433), .C1(n63501), .C2(n67427), .A(
        n65115), .ZN(n65106) );
  AOI22_X1 U49209 ( .A1(n67421), .A2(n66308), .B1(n67415), .B2(n58303), .ZN(
        n65115) );
  OAI221_X1 U49210 ( .B1(n54610), .B2(n67433), .C1(n63505), .C2(n67427), .A(
        n65196), .ZN(n65193) );
  AOI22_X1 U49211 ( .A1(n67421), .A2(n66305), .B1(n67415), .B2(n58304), .ZN(
        n65196) );
  OAI221_X1 U49212 ( .B1(n54609), .B2(n67433), .C1(n63504), .C2(n67427), .A(
        n65178), .ZN(n65175) );
  AOI22_X1 U49213 ( .A1(n67421), .A2(n66306), .B1(n67415), .B2(n58305), .ZN(
        n65178) );
  OAI221_X1 U49214 ( .B1(n62426), .B2(n67409), .C1(n63635), .C2(n67403), .A(
        n65161), .ZN(n65156) );
  AOI22_X1 U49215 ( .A1(n67397), .A2(n58781), .B1(n67391), .B2(n58369), .ZN(
        n65161) );
  OAI221_X1 U49216 ( .B1(n62424), .B2(n67409), .C1(n63633), .C2(n67403), .A(
        n65120), .ZN(n65105) );
  AOI22_X1 U49217 ( .A1(n67397), .A2(n58782), .B1(n67391), .B2(n58370), .ZN(
        n65120) );
  OAI221_X1 U49218 ( .B1(n62428), .B2(n67409), .C1(n63637), .C2(n67403), .A(
        n65197), .ZN(n65192) );
  AOI22_X1 U49219 ( .A1(n67397), .A2(n58779), .B1(n67391), .B2(n58367), .ZN(
        n65197) );
  OAI221_X1 U49220 ( .B1(n62427), .B2(n67409), .C1(n63636), .C2(n67403), .A(
        n65179), .ZN(n65174) );
  AOI22_X1 U49221 ( .A1(n67397), .A2(n58780), .B1(n67391), .B2(n58368), .ZN(
        n65179) );
  OAI221_X1 U49222 ( .B1(n62428), .B2(n67607), .C1(n63505), .C2(n67601), .A(
        n63873), .ZN(n63868) );
  AOI22_X1 U49223 ( .A1(n67595), .A2(n66499), .B1(n58375), .B2(n67589), .ZN(
        n63873) );
  OAI221_X1 U49224 ( .B1(n62427), .B2(n67607), .C1(n63504), .C2(n67601), .A(
        n63852), .ZN(n63847) );
  AOI22_X1 U49225 ( .A1(n67595), .A2(n66500), .B1(n58376), .B2(n67589), .ZN(
        n63852) );
  OAI221_X1 U49226 ( .B1(n62426), .B2(n67607), .C1(n63503), .C2(n67601), .A(
        n63831), .ZN(n63826) );
  AOI22_X1 U49227 ( .A1(n67595), .A2(n66501), .B1(n58377), .B2(n67589), .ZN(
        n63831) );
  OAI221_X1 U49228 ( .B1(n63569), .B2(n67385), .C1(n8481), .C2(n67379), .A(
        n65162), .ZN(n65155) );
  AOI22_X1 U49229 ( .A1(n67373), .A2(n66497), .B1(n67367), .B2(n8896), .ZN(
        n65162) );
  OAI221_X1 U49230 ( .B1(n63567), .B2(n67385), .C1(n8497), .C2(n67379), .A(
        n65125), .ZN(n65104) );
  AOI22_X1 U49231 ( .A1(n67373), .A2(n66498), .B1(n67367), .B2(n8895), .ZN(
        n65125) );
  OAI221_X1 U49232 ( .B1(n63571), .B2(n67385), .C1(n8449), .C2(n67379), .A(
        n65198), .ZN(n65191) );
  AOI22_X1 U49233 ( .A1(n67373), .A2(n66495), .B1(n67367), .B2(n8898), .ZN(
        n65198) );
  OAI221_X1 U49234 ( .B1(n63570), .B2(n67385), .C1(n8465), .C2(n67379), .A(
        n65180), .ZN(n65173) );
  AOI22_X1 U49235 ( .A1(n67373), .A2(n66496), .B1(n67367), .B2(n8897), .ZN(
        n65180) );
  OAI221_X1 U49236 ( .B1(n54186), .B2(n67583), .C1(n63571), .C2(n67577), .A(
        n63875), .ZN(n63867) );
  AOI22_X1 U49237 ( .A1(n67571), .A2(n8965), .B1(n67565), .B2(n66495), .ZN(
        n63875) );
  OAI221_X1 U49238 ( .B1(n54185), .B2(n67583), .C1(n63570), .C2(n67577), .A(
        n63854), .ZN(n63846) );
  AOI22_X1 U49239 ( .A1(n67571), .A2(n8963), .B1(n67565), .B2(n66496), .ZN(
        n63854) );
  OAI221_X1 U49240 ( .B1(n54184), .B2(n67583), .C1(n63569), .C2(n67577), .A(
        n63833), .ZN(n63825) );
  AOI22_X1 U49241 ( .A1(n67571), .A2(n8961), .B1(n67565), .B2(n66497), .ZN(
        n63833) );
  OAI221_X1 U49242 ( .B1(n62694), .B2(n67583), .C1(n63567), .C2(n67577), .A(
        n63793), .ZN(n63771) );
  AOI22_X1 U49243 ( .A1(n67571), .A2(n8959), .B1(n67565), .B2(n66498), .ZN(
        n63793) );
  OAI221_X1 U49244 ( .B1(n54246), .B2(n67578), .C1(n63631), .C2(n67572), .A(
        n65088), .ZN(n65068) );
  AOI22_X1 U49245 ( .A1(n67566), .A2(n9085), .B1(n67560), .B2(n58036), .ZN(
        n65088) );
  OAI221_X1 U49246 ( .B1(n54245), .B2(n67578), .C1(n63630), .C2(n67572), .A(
        n65056), .ZN(n65048) );
  AOI22_X1 U49247 ( .A1(n67566), .A2(n9083), .B1(n67560), .B2(n58001), .ZN(
        n65056) );
  OAI221_X1 U49248 ( .B1(n54244), .B2(n67578), .C1(n63629), .C2(n67572), .A(
        n65036), .ZN(n65028) );
  AOI22_X1 U49249 ( .A1(n67566), .A2(n9081), .B1(n67560), .B2(n57977), .ZN(
        n65036) );
  OAI221_X1 U49250 ( .B1(n54243), .B2(n67578), .C1(n63628), .C2(n67572), .A(
        n65016), .ZN(n65008) );
  AOI22_X1 U49251 ( .A1(n67566), .A2(n9079), .B1(n67560), .B2(n57953), .ZN(
        n65016) );
  OAI221_X1 U49252 ( .B1(n54242), .B2(n67578), .C1(n63627), .C2(n67572), .A(
        n64996), .ZN(n64988) );
  AOI22_X1 U49253 ( .A1(n67566), .A2(n9077), .B1(n67560), .B2(n57929), .ZN(
        n64996) );
  OAI221_X1 U49254 ( .B1(n54241), .B2(n67578), .C1(n63626), .C2(n67572), .A(
        n64976), .ZN(n64968) );
  AOI22_X1 U49255 ( .A1(n67566), .A2(n9075), .B1(n67560), .B2(n57905), .ZN(
        n64976) );
  OAI221_X1 U49256 ( .B1(n54240), .B2(n67578), .C1(n63625), .C2(n67572), .A(
        n64956), .ZN(n64948) );
  AOI22_X1 U49257 ( .A1(n67566), .A2(n9073), .B1(n67560), .B2(n57881), .ZN(
        n64956) );
  OAI221_X1 U49258 ( .B1(n54239), .B2(n67578), .C1(n63624), .C2(n67572), .A(
        n64936), .ZN(n64928) );
  AOI22_X1 U49259 ( .A1(n67566), .A2(n9071), .B1(n67560), .B2(n57857), .ZN(
        n64936) );
  OAI221_X1 U49260 ( .B1(n54238), .B2(n67578), .C1(n63623), .C2(n67572), .A(
        n64916), .ZN(n64908) );
  AOI22_X1 U49261 ( .A1(n67566), .A2(n9069), .B1(n67560), .B2(n57833), .ZN(
        n64916) );
  OAI221_X1 U49262 ( .B1(n54237), .B2(n67578), .C1(n63622), .C2(n67572), .A(
        n64896), .ZN(n64888) );
  AOI22_X1 U49263 ( .A1(n67566), .A2(n9067), .B1(n67560), .B2(n57809), .ZN(
        n64896) );
  OAI221_X1 U49264 ( .B1(n54236), .B2(n67578), .C1(n63621), .C2(n67572), .A(
        n64876), .ZN(n64868) );
  AOI22_X1 U49265 ( .A1(n67566), .A2(n9065), .B1(n67560), .B2(n57785), .ZN(
        n64876) );
  OAI221_X1 U49266 ( .B1(n54235), .B2(n67578), .C1(n63620), .C2(n67572), .A(
        n64856), .ZN(n64848) );
  AOI22_X1 U49267 ( .A1(n67566), .A2(n9063), .B1(n67560), .B2(n57761), .ZN(
        n64856) );
  OAI22_X1 U49268 ( .A1(n54184), .A2(n67361), .B1(n49482), .B2(n67355), .ZN(
        n65166) );
  OAI22_X1 U49269 ( .A1(n62694), .A2(n67361), .B1(n49483), .B2(n67355), .ZN(
        n65131) );
  OAI22_X1 U49270 ( .A1(n54186), .A2(n67361), .B1(n49480), .B2(n67355), .ZN(
        n65202) );
  OAI22_X1 U49271 ( .A1(n54185), .A2(n67361), .B1(n49481), .B2(n67355), .ZN(
        n65184) );
  OAI22_X1 U49272 ( .A1(n62691), .A2(n67554), .B1(n54670), .B2(n67548), .ZN(
        n65092) );
  OAI22_X1 U49273 ( .A1(n62690), .A2(n67554), .B1(n54669), .B2(n67548), .ZN(
        n65060) );
  OAI22_X1 U49274 ( .A1(n62689), .A2(n67554), .B1(n54668), .B2(n67548), .ZN(
        n65040) );
  OAI22_X1 U49275 ( .A1(n62688), .A2(n67554), .B1(n54667), .B2(n67548), .ZN(
        n65020) );
  OAI22_X1 U49276 ( .A1(n62687), .A2(n67554), .B1(n54666), .B2(n67548), .ZN(
        n65000) );
  OAI22_X1 U49277 ( .A1(n62686), .A2(n67554), .B1(n54665), .B2(n67548), .ZN(
        n64980) );
  OAI22_X1 U49278 ( .A1(n62685), .A2(n67554), .B1(n54664), .B2(n67548), .ZN(
        n64960) );
  OAI22_X1 U49279 ( .A1(n62684), .A2(n67554), .B1(n54663), .B2(n67548), .ZN(
        n64940) );
  OAI22_X1 U49280 ( .A1(n62683), .A2(n67554), .B1(n54662), .B2(n67548), .ZN(
        n64920) );
  OAI22_X1 U49281 ( .A1(n62682), .A2(n67554), .B1(n54661), .B2(n67548), .ZN(
        n64900) );
  OAI22_X1 U49282 ( .A1(n62681), .A2(n67554), .B1(n54660), .B2(n67548), .ZN(
        n64880) );
  OAI22_X1 U49283 ( .A1(n62680), .A2(n67554), .B1(n54659), .B2(n67548), .ZN(
        n64860) );
  OAI22_X1 U49284 ( .A1(n62679), .A2(n67555), .B1(n54658), .B2(n67549), .ZN(
        n64840) );
  OAI22_X1 U49285 ( .A1(n62678), .A2(n67555), .B1(n54657), .B2(n67549), .ZN(
        n64820) );
  OAI22_X1 U49286 ( .A1(n62677), .A2(n67555), .B1(n54656), .B2(n67549), .ZN(
        n64800) );
  OAI22_X1 U49287 ( .A1(n62676), .A2(n67555), .B1(n54655), .B2(n67549), .ZN(
        n64780) );
  OAI22_X1 U49288 ( .A1(n62675), .A2(n67555), .B1(n54654), .B2(n67549), .ZN(
        n64760) );
  OAI22_X1 U49289 ( .A1(n62674), .A2(n67555), .B1(n54653), .B2(n67549), .ZN(
        n64740) );
  OAI22_X1 U49290 ( .A1(n62673), .A2(n67555), .B1(n54652), .B2(n67549), .ZN(
        n64720) );
  OAI22_X1 U49291 ( .A1(n62672), .A2(n67555), .B1(n54651), .B2(n67549), .ZN(
        n64700) );
  OAI22_X1 U49292 ( .A1(n62671), .A2(n67555), .B1(n54650), .B2(n67549), .ZN(
        n64680) );
  OAI22_X1 U49293 ( .A1(n62670), .A2(n67555), .B1(n54649), .B2(n67549), .ZN(
        n64660) );
  OAI22_X1 U49294 ( .A1(n62669), .A2(n67555), .B1(n54648), .B2(n67549), .ZN(
        n64640) );
  OAI22_X1 U49295 ( .A1(n62668), .A2(n67555), .B1(n54647), .B2(n67549), .ZN(
        n64620) );
  OAI22_X1 U49296 ( .A1(n62667), .A2(n67556), .B1(n54646), .B2(n67550), .ZN(
        n64600) );
  OAI22_X1 U49297 ( .A1(n62666), .A2(n67556), .B1(n54645), .B2(n67550), .ZN(
        n64580) );
  OAI22_X1 U49298 ( .A1(n62665), .A2(n67556), .B1(n54644), .B2(n67550), .ZN(
        n64560) );
  OAI22_X1 U49299 ( .A1(n62664), .A2(n67556), .B1(n54643), .B2(n67550), .ZN(
        n64540) );
  OAI22_X1 U49300 ( .A1(n62663), .A2(n67556), .B1(n54642), .B2(n67550), .ZN(
        n64520) );
  OAI22_X1 U49301 ( .A1(n62662), .A2(n67556), .B1(n54641), .B2(n67550), .ZN(
        n64500) );
  OAI22_X1 U49302 ( .A1(n62661), .A2(n67556), .B1(n54640), .B2(n67550), .ZN(
        n64480) );
  OAI22_X1 U49303 ( .A1(n62660), .A2(n67556), .B1(n54639), .B2(n67550), .ZN(
        n64460) );
  OAI22_X1 U49304 ( .A1(n62659), .A2(n67556), .B1(n54638), .B2(n67550), .ZN(
        n64440) );
  OAI22_X1 U49305 ( .A1(n62658), .A2(n67556), .B1(n54637), .B2(n67550), .ZN(
        n64420) );
  OAI22_X1 U49306 ( .A1(n62657), .A2(n67556), .B1(n54636), .B2(n67550), .ZN(
        n64400) );
  OAI22_X1 U49307 ( .A1(n62656), .A2(n67556), .B1(n54635), .B2(n67550), .ZN(
        n64380) );
  OAI22_X1 U49308 ( .A1(n62655), .A2(n67557), .B1(n54634), .B2(n67551), .ZN(
        n64360) );
  OAI22_X1 U49309 ( .A1(n62654), .A2(n67557), .B1(n54633), .B2(n67551), .ZN(
        n64340) );
  OAI22_X1 U49310 ( .A1(n62653), .A2(n67557), .B1(n54632), .B2(n67551), .ZN(
        n64320) );
  OAI22_X1 U49311 ( .A1(n62652), .A2(n67557), .B1(n54631), .B2(n67551), .ZN(
        n64300) );
  OAI22_X1 U49312 ( .A1(n62651), .A2(n67557), .B1(n54630), .B2(n67551), .ZN(
        n64280) );
  OAI22_X1 U49313 ( .A1(n62650), .A2(n67557), .B1(n54629), .B2(n67551), .ZN(
        n64260) );
  OAI22_X1 U49314 ( .A1(n62649), .A2(n67557), .B1(n54628), .B2(n67551), .ZN(
        n64240) );
  OAI22_X1 U49315 ( .A1(n62648), .A2(n67557), .B1(n54627), .B2(n67551), .ZN(
        n64220) );
  OAI22_X1 U49316 ( .A1(n62647), .A2(n67557), .B1(n54626), .B2(n67551), .ZN(
        n64200) );
  OAI22_X1 U49317 ( .A1(n62646), .A2(n67557), .B1(n54625), .B2(n67551), .ZN(
        n64180) );
  OAI22_X1 U49318 ( .A1(n62645), .A2(n67557), .B1(n54624), .B2(n67551), .ZN(
        n64160) );
  OAI22_X1 U49319 ( .A1(n62644), .A2(n67557), .B1(n54623), .B2(n67551), .ZN(
        n64140) );
  OAI22_X1 U49320 ( .A1(n62643), .A2(n67558), .B1(n54622), .B2(n67552), .ZN(
        n64120) );
  OAI22_X1 U49321 ( .A1(n62642), .A2(n67558), .B1(n54621), .B2(n67552), .ZN(
        n64100) );
  OAI22_X1 U49322 ( .A1(n62641), .A2(n67558), .B1(n54620), .B2(n67552), .ZN(
        n64080) );
  OAI22_X1 U49323 ( .A1(n62640), .A2(n67558), .B1(n54619), .B2(n67552), .ZN(
        n64060) );
  OAI22_X1 U49324 ( .A1(n62639), .A2(n67558), .B1(n54618), .B2(n67552), .ZN(
        n64040) );
  OAI22_X1 U49325 ( .A1(n62638), .A2(n67558), .B1(n54617), .B2(n67552), .ZN(
        n64020) );
  OAI22_X1 U49326 ( .A1(n62637), .A2(n67558), .B1(n54616), .B2(n67552), .ZN(
        n64000) );
  OAI22_X1 U49327 ( .A1(n62636), .A2(n67558), .B1(n54615), .B2(n67552), .ZN(
        n63980) );
  OAI22_X1 U49328 ( .A1(n62635), .A2(n67558), .B1(n54614), .B2(n67552), .ZN(
        n63960) );
  OAI22_X1 U49329 ( .A1(n62634), .A2(n67558), .B1(n54613), .B2(n67552), .ZN(
        n63940) );
  OAI22_X1 U49330 ( .A1(n62633), .A2(n67558), .B1(n54612), .B2(n67552), .ZN(
        n63920) );
  OAI22_X1 U49331 ( .A1(n62632), .A2(n67558), .B1(n54611), .B2(n67552), .ZN(
        n63900) );
  OAI22_X1 U49332 ( .A1(n54246), .A2(n67356), .B1(n49420), .B2(n67350), .ZN(
        n66296) );
  OAI22_X1 U49333 ( .A1(n54245), .A2(n67356), .B1(n49421), .B2(n67350), .ZN(
        n66264) );
  OAI22_X1 U49334 ( .A1(n54244), .A2(n67356), .B1(n49422), .B2(n67350), .ZN(
        n66246) );
  OAI22_X1 U49335 ( .A1(n54243), .A2(n67356), .B1(n49423), .B2(n67350), .ZN(
        n66228) );
  OAI22_X1 U49336 ( .A1(n54242), .A2(n67356), .B1(n49424), .B2(n67350), .ZN(
        n66210) );
  OAI22_X1 U49337 ( .A1(n54241), .A2(n67356), .B1(n49425), .B2(n67350), .ZN(
        n66192) );
  OAI22_X1 U49338 ( .A1(n54240), .A2(n67356), .B1(n49426), .B2(n67350), .ZN(
        n66174) );
  OAI22_X1 U49339 ( .A1(n54239), .A2(n67356), .B1(n49427), .B2(n67350), .ZN(
        n66156) );
  OAI22_X1 U49340 ( .A1(n54238), .A2(n67356), .B1(n49428), .B2(n67350), .ZN(
        n66138) );
  OAI22_X1 U49341 ( .A1(n54237), .A2(n67356), .B1(n49429), .B2(n67350), .ZN(
        n66120) );
  OAI22_X1 U49342 ( .A1(n54236), .A2(n67356), .B1(n49430), .B2(n67350), .ZN(
        n66102) );
  OAI22_X1 U49343 ( .A1(n54235), .A2(n67356), .B1(n49431), .B2(n67350), .ZN(
        n66084) );
  OAI22_X1 U49344 ( .A1(n54234), .A2(n67357), .B1(n49432), .B2(n67351), .ZN(
        n66066) );
  OAI22_X1 U49345 ( .A1(n54233), .A2(n67357), .B1(n49433), .B2(n67351), .ZN(
        n66048) );
  OAI22_X1 U49346 ( .A1(n54232), .A2(n67357), .B1(n49434), .B2(n67351), .ZN(
        n66030) );
  OAI22_X1 U49347 ( .A1(n54231), .A2(n67357), .B1(n49435), .B2(n67351), .ZN(
        n66012) );
  OAI22_X1 U49348 ( .A1(n54230), .A2(n67357), .B1(n49436), .B2(n67351), .ZN(
        n65994) );
  OAI22_X1 U49349 ( .A1(n54229), .A2(n67357), .B1(n49437), .B2(n67351), .ZN(
        n65976) );
  OAI22_X1 U49350 ( .A1(n54228), .A2(n67357), .B1(n49438), .B2(n67351), .ZN(
        n65958) );
  OAI22_X1 U49351 ( .A1(n54227), .A2(n67357), .B1(n49439), .B2(n67351), .ZN(
        n65940) );
  OAI22_X1 U49352 ( .A1(n54226), .A2(n67357), .B1(n49440), .B2(n67351), .ZN(
        n65922) );
  OAI22_X1 U49353 ( .A1(n54225), .A2(n67357), .B1(n49441), .B2(n67351), .ZN(
        n65904) );
  OAI22_X1 U49354 ( .A1(n54224), .A2(n67357), .B1(n49442), .B2(n67351), .ZN(
        n65886) );
  OAI22_X1 U49355 ( .A1(n54223), .A2(n67357), .B1(n49443), .B2(n67351), .ZN(
        n65868) );
  OAI22_X1 U49356 ( .A1(n54222), .A2(n67358), .B1(n49444), .B2(n67352), .ZN(
        n65850) );
  OAI22_X1 U49357 ( .A1(n54221), .A2(n67358), .B1(n49445), .B2(n67352), .ZN(
        n65832) );
  OAI22_X1 U49358 ( .A1(n54220), .A2(n67358), .B1(n49446), .B2(n67352), .ZN(
        n65814) );
  OAI22_X1 U49359 ( .A1(n54219), .A2(n67358), .B1(n49447), .B2(n67352), .ZN(
        n65796) );
  OAI22_X1 U49360 ( .A1(n54218), .A2(n67358), .B1(n49448), .B2(n67352), .ZN(
        n65778) );
  OAI22_X1 U49361 ( .A1(n54217), .A2(n67358), .B1(n49449), .B2(n67352), .ZN(
        n65760) );
  OAI22_X1 U49362 ( .A1(n54216), .A2(n67358), .B1(n49450), .B2(n67352), .ZN(
        n65742) );
  OAI22_X1 U49363 ( .A1(n54215), .A2(n67358), .B1(n49451), .B2(n67352), .ZN(
        n65724) );
  OAI22_X1 U49364 ( .A1(n54214), .A2(n67358), .B1(n49452), .B2(n67352), .ZN(
        n65706) );
  OAI22_X1 U49365 ( .A1(n54213), .A2(n67358), .B1(n49453), .B2(n67352), .ZN(
        n65688) );
  OAI22_X1 U49366 ( .A1(n54212), .A2(n67358), .B1(n49454), .B2(n67352), .ZN(
        n65670) );
  OAI22_X1 U49367 ( .A1(n54211), .A2(n67358), .B1(n49455), .B2(n67352), .ZN(
        n65652) );
  OAI22_X1 U49368 ( .A1(n54210), .A2(n67359), .B1(n49456), .B2(n67353), .ZN(
        n65634) );
  OAI22_X1 U49369 ( .A1(n54209), .A2(n67359), .B1(n49457), .B2(n67353), .ZN(
        n65616) );
  OAI22_X1 U49370 ( .A1(n54208), .A2(n67359), .B1(n49458), .B2(n67353), .ZN(
        n65598) );
  OAI22_X1 U49371 ( .A1(n54207), .A2(n67359), .B1(n49459), .B2(n67353), .ZN(
        n65580) );
  OAI22_X1 U49372 ( .A1(n54206), .A2(n67359), .B1(n49460), .B2(n67353), .ZN(
        n65562) );
  OAI22_X1 U49373 ( .A1(n54205), .A2(n67359), .B1(n49461), .B2(n67353), .ZN(
        n65544) );
  OAI22_X1 U49374 ( .A1(n54204), .A2(n67359), .B1(n49462), .B2(n67353), .ZN(
        n65526) );
  OAI22_X1 U49375 ( .A1(n54203), .A2(n67359), .B1(n49463), .B2(n67353), .ZN(
        n65508) );
  OAI22_X1 U49376 ( .A1(n54202), .A2(n67359), .B1(n49464), .B2(n67353), .ZN(
        n65490) );
  OAI22_X1 U49377 ( .A1(n54201), .A2(n67359), .B1(n49465), .B2(n67353), .ZN(
        n65472) );
  OAI22_X1 U49378 ( .A1(n54200), .A2(n67359), .B1(n49466), .B2(n67353), .ZN(
        n65454) );
  OAI22_X1 U49379 ( .A1(n54199), .A2(n67359), .B1(n49467), .B2(n67353), .ZN(
        n65436) );
  OAI22_X1 U49380 ( .A1(n54198), .A2(n67360), .B1(n49468), .B2(n67354), .ZN(
        n65418) );
  OAI22_X1 U49381 ( .A1(n54197), .A2(n67360), .B1(n49469), .B2(n67354), .ZN(
        n65400) );
  OAI22_X1 U49382 ( .A1(n54196), .A2(n67360), .B1(n49470), .B2(n67354), .ZN(
        n65382) );
  OAI22_X1 U49383 ( .A1(n54195), .A2(n67360), .B1(n49471), .B2(n67354), .ZN(
        n65364) );
  OAI22_X1 U49384 ( .A1(n54194), .A2(n67360), .B1(n49472), .B2(n67354), .ZN(
        n65346) );
  OAI22_X1 U49385 ( .A1(n54193), .A2(n67360), .B1(n49473), .B2(n67354), .ZN(
        n65328) );
  OAI22_X1 U49386 ( .A1(n54192), .A2(n67360), .B1(n49474), .B2(n67354), .ZN(
        n65310) );
  OAI22_X1 U49387 ( .A1(n54191), .A2(n67360), .B1(n49475), .B2(n67354), .ZN(
        n65292) );
  OAI22_X1 U49388 ( .A1(n54190), .A2(n67360), .B1(n49476), .B2(n67354), .ZN(
        n65274) );
  OAI22_X1 U49389 ( .A1(n54189), .A2(n67360), .B1(n49477), .B2(n67354), .ZN(
        n65256) );
  OAI22_X1 U49390 ( .A1(n54188), .A2(n67360), .B1(n49478), .B2(n67354), .ZN(
        n65238) );
  OAI22_X1 U49391 ( .A1(n54187), .A2(n67360), .B1(n49479), .B2(n67354), .ZN(
        n65220) );
  OAI22_X1 U49392 ( .A1(n7489), .A2(n67542), .B1(n62422), .B2(n67536), .ZN(
        n65091) );
  OAI22_X1 U49393 ( .A1(n7505), .A2(n67542), .B1(n62421), .B2(n67536), .ZN(
        n65059) );
  OAI22_X1 U49394 ( .A1(n7521), .A2(n67542), .B1(n62420), .B2(n67536), .ZN(
        n65039) );
  OAI22_X1 U49395 ( .A1(n7537), .A2(n67542), .B1(n62419), .B2(n67536), .ZN(
        n65019) );
  OAI22_X1 U49396 ( .A1(n7553), .A2(n67542), .B1(n62418), .B2(n67536), .ZN(
        n64999) );
  OAI22_X1 U49397 ( .A1(n7569), .A2(n67542), .B1(n62417), .B2(n67536), .ZN(
        n64979) );
  OAI22_X1 U49398 ( .A1(n7585), .A2(n67542), .B1(n62416), .B2(n67536), .ZN(
        n64959) );
  OAI22_X1 U49399 ( .A1(n7601), .A2(n67542), .B1(n62415), .B2(n67536), .ZN(
        n64939) );
  OAI22_X1 U49400 ( .A1(n7617), .A2(n67542), .B1(n62414), .B2(n67536), .ZN(
        n64919) );
  OAI22_X1 U49401 ( .A1(n7633), .A2(n67542), .B1(n62413), .B2(n67536), .ZN(
        n64899) );
  OAI22_X1 U49402 ( .A1(n7649), .A2(n67542), .B1(n62412), .B2(n67536), .ZN(
        n64879) );
  OAI22_X1 U49403 ( .A1(n7665), .A2(n67542), .B1(n62411), .B2(n67536), .ZN(
        n64859) );
  OAI22_X1 U49404 ( .A1(n7681), .A2(n67543), .B1(n62410), .B2(n67537), .ZN(
        n64839) );
  OAI22_X1 U49405 ( .A1(n7697), .A2(n67543), .B1(n62409), .B2(n67537), .ZN(
        n64819) );
  OAI22_X1 U49406 ( .A1(n7713), .A2(n67543), .B1(n62408), .B2(n67537), .ZN(
        n64799) );
  OAI22_X1 U49407 ( .A1(n7729), .A2(n67543), .B1(n62407), .B2(n67537), .ZN(
        n64779) );
  OAI22_X1 U49408 ( .A1(n7745), .A2(n67543), .B1(n62406), .B2(n67537), .ZN(
        n64759) );
  OAI22_X1 U49409 ( .A1(n7761), .A2(n67543), .B1(n62405), .B2(n67537), .ZN(
        n64739) );
  OAI22_X1 U49410 ( .A1(n7777), .A2(n67543), .B1(n62404), .B2(n67537), .ZN(
        n64719) );
  OAI22_X1 U49411 ( .A1(n7793), .A2(n67543), .B1(n62403), .B2(n67537), .ZN(
        n64699) );
  OAI22_X1 U49412 ( .A1(n7809), .A2(n67543), .B1(n62402), .B2(n67537), .ZN(
        n64679) );
  OAI22_X1 U49413 ( .A1(n7825), .A2(n67543), .B1(n62401), .B2(n67537), .ZN(
        n64659) );
  OAI22_X1 U49414 ( .A1(n7841), .A2(n67543), .B1(n62400), .B2(n67537), .ZN(
        n64639) );
  OAI22_X1 U49415 ( .A1(n7857), .A2(n67543), .B1(n62399), .B2(n67537), .ZN(
        n64619) );
  OAI22_X1 U49416 ( .A1(n7873), .A2(n67544), .B1(n62398), .B2(n67538), .ZN(
        n64599) );
  OAI22_X1 U49417 ( .A1(n7889), .A2(n67544), .B1(n62397), .B2(n67538), .ZN(
        n64579) );
  OAI22_X1 U49418 ( .A1(n7905), .A2(n67544), .B1(n62396), .B2(n67538), .ZN(
        n64559) );
  OAI22_X1 U49419 ( .A1(n7921), .A2(n67544), .B1(n62395), .B2(n67538), .ZN(
        n64539) );
  OAI22_X1 U49420 ( .A1(n7937), .A2(n67544), .B1(n62394), .B2(n67538), .ZN(
        n64519) );
  OAI22_X1 U49421 ( .A1(n7953), .A2(n67544), .B1(n62393), .B2(n67538), .ZN(
        n64499) );
  OAI22_X1 U49422 ( .A1(n7969), .A2(n67544), .B1(n62392), .B2(n67538), .ZN(
        n64479) );
  OAI22_X1 U49423 ( .A1(n7985), .A2(n67544), .B1(n62391), .B2(n67538), .ZN(
        n64459) );
  OAI22_X1 U49424 ( .A1(n8001), .A2(n67544), .B1(n62390), .B2(n67538), .ZN(
        n64439) );
  OAI22_X1 U49425 ( .A1(n8017), .A2(n67544), .B1(n62389), .B2(n67538), .ZN(
        n64419) );
  OAI22_X1 U49426 ( .A1(n8033), .A2(n67544), .B1(n62388), .B2(n67538), .ZN(
        n64399) );
  OAI22_X1 U49427 ( .A1(n8049), .A2(n67544), .B1(n62387), .B2(n67538), .ZN(
        n64379) );
  OAI22_X1 U49428 ( .A1(n8065), .A2(n67545), .B1(n62386), .B2(n67539), .ZN(
        n64359) );
  OAI22_X1 U49429 ( .A1(n8081), .A2(n67545), .B1(n62385), .B2(n67539), .ZN(
        n64339) );
  OAI22_X1 U49430 ( .A1(n8097), .A2(n67545), .B1(n62384), .B2(n67539), .ZN(
        n64319) );
  OAI22_X1 U49431 ( .A1(n8113), .A2(n67545), .B1(n62383), .B2(n67539), .ZN(
        n64299) );
  OAI22_X1 U49432 ( .A1(n8129), .A2(n67545), .B1(n62382), .B2(n67539), .ZN(
        n64279) );
  OAI22_X1 U49433 ( .A1(n8145), .A2(n67545), .B1(n62381), .B2(n67539), .ZN(
        n64259) );
  OAI22_X1 U49434 ( .A1(n8161), .A2(n67545), .B1(n62380), .B2(n67539), .ZN(
        n64239) );
  OAI22_X1 U49435 ( .A1(n8177), .A2(n67545), .B1(n62379), .B2(n67539), .ZN(
        n64219) );
  OAI22_X1 U49436 ( .A1(n8193), .A2(n67545), .B1(n62378), .B2(n67539), .ZN(
        n64199) );
  OAI22_X1 U49437 ( .A1(n8209), .A2(n67545), .B1(n62377), .B2(n67539), .ZN(
        n64179) );
  OAI22_X1 U49438 ( .A1(n8225), .A2(n67545), .B1(n62376), .B2(n67539), .ZN(
        n64159) );
  OAI22_X1 U49439 ( .A1(n8241), .A2(n67545), .B1(n62375), .B2(n67539), .ZN(
        n64139) );
  OAI22_X1 U49440 ( .A1(n8257), .A2(n67546), .B1(n62374), .B2(n67540), .ZN(
        n64119) );
  OAI22_X1 U49441 ( .A1(n8273), .A2(n67546), .B1(n62373), .B2(n67540), .ZN(
        n64099) );
  OAI22_X1 U49442 ( .A1(n8289), .A2(n67546), .B1(n62372), .B2(n67540), .ZN(
        n64079) );
  OAI22_X1 U49443 ( .A1(n8305), .A2(n67546), .B1(n62371), .B2(n67540), .ZN(
        n64059) );
  OAI22_X1 U49444 ( .A1(n8321), .A2(n67546), .B1(n62370), .B2(n67540), .ZN(
        n64039) );
  OAI22_X1 U49445 ( .A1(n8337), .A2(n67546), .B1(n62369), .B2(n67540), .ZN(
        n64019) );
  OAI22_X1 U49446 ( .A1(n8353), .A2(n67546), .B1(n62368), .B2(n67540), .ZN(
        n63999) );
  OAI22_X1 U49447 ( .A1(n8369), .A2(n67546), .B1(n62367), .B2(n67540), .ZN(
        n63979) );
  OAI22_X1 U49448 ( .A1(n8385), .A2(n67546), .B1(n62366), .B2(n67540), .ZN(
        n63959) );
  OAI22_X1 U49449 ( .A1(n8401), .A2(n67546), .B1(n62365), .B2(n67540), .ZN(
        n63939) );
  OAI22_X1 U49450 ( .A1(n8417), .A2(n67546), .B1(n62364), .B2(n67540), .ZN(
        n63919) );
  OAI22_X1 U49451 ( .A1(n8433), .A2(n67546), .B1(n62363), .B2(n67540), .ZN(
        n63899) );
  AND3_X1 U49452 ( .A1(ADD_RD1[2]), .A2(n66494), .A3(ADD_RD1[1]), .ZN(n65074)
         );
  OAI22_X1 U49453 ( .A1(n68259), .A2(n62061), .B1(n68251), .B2(n68094), .ZN(
        n7435) );
  OAI22_X1 U49454 ( .A1(n68259), .A2(n62059), .B1(n68251), .B2(n68097), .ZN(
        n7436) );
  OAI22_X1 U49455 ( .A1(n68259), .A2(n62057), .B1(n68251), .B2(n68100), .ZN(
        n7437) );
  OAI22_X1 U49456 ( .A1(n68259), .A2(n62055), .B1(n68251), .B2(n68103), .ZN(
        n7438) );
  OAI22_X1 U49457 ( .A1(n68259), .A2(n62053), .B1(n68251), .B2(n68106), .ZN(
        n7439) );
  OAI22_X1 U49458 ( .A1(n68259), .A2(n62051), .B1(n68251), .B2(n68109), .ZN(
        n7440) );
  OAI22_X1 U49459 ( .A1(n68259), .A2(n62049), .B1(n68251), .B2(n68112), .ZN(
        n7441) );
  OAI22_X1 U49460 ( .A1(n68259), .A2(n62047), .B1(n68251), .B2(n68115), .ZN(
        n7442) );
  OAI22_X1 U49461 ( .A1(n68259), .A2(n62045), .B1(n68251), .B2(n68118), .ZN(
        n7443) );
  OAI22_X1 U49462 ( .A1(n68259), .A2(n62043), .B1(n68251), .B2(n68121), .ZN(
        n7444) );
  OAI22_X1 U49463 ( .A1(n68259), .A2(n62041), .B1(n68251), .B2(n68124), .ZN(
        n7445) );
  OAI22_X1 U49464 ( .A1(n68259), .A2(n62039), .B1(n68251), .B2(n68127), .ZN(
        n7446) );
  OAI22_X1 U49465 ( .A1(n68259), .A2(n62037), .B1(n68252), .B2(n68130), .ZN(
        n7447) );
  OAI22_X1 U49466 ( .A1(n68260), .A2(n62035), .B1(n68252), .B2(n68133), .ZN(
        n7448) );
  OAI22_X1 U49467 ( .A1(n68260), .A2(n62033), .B1(n68252), .B2(n68136), .ZN(
        n7449) );
  OAI22_X1 U49468 ( .A1(n68260), .A2(n62031), .B1(n68252), .B2(n68139), .ZN(
        n7450) );
  OAI22_X1 U49469 ( .A1(n68260), .A2(n62029), .B1(n68252), .B2(n68142), .ZN(
        n7451) );
  OAI22_X1 U49470 ( .A1(n68260), .A2(n62027), .B1(n68252), .B2(n68145), .ZN(
        n7452) );
  OAI22_X1 U49471 ( .A1(n68260), .A2(n62025), .B1(n68252), .B2(n68148), .ZN(
        n7453) );
  OAI22_X1 U49472 ( .A1(n68260), .A2(n62023), .B1(n68252), .B2(n68151), .ZN(
        n7454) );
  OAI22_X1 U49473 ( .A1(n68260), .A2(n62021), .B1(n68252), .B2(n68154), .ZN(
        n7455) );
  OAI22_X1 U49474 ( .A1(n68260), .A2(n62019), .B1(n68252), .B2(n68157), .ZN(
        n7456) );
  OAI22_X1 U49475 ( .A1(n68260), .A2(n62017), .B1(n68252), .B2(n68160), .ZN(
        n7457) );
  OAI22_X1 U49476 ( .A1(n68260), .A2(n62015), .B1(n68252), .B2(n68163), .ZN(
        n7458) );
  OAI22_X1 U49477 ( .A1(n68260), .A2(n62013), .B1(n68253), .B2(n68166), .ZN(
        n7459) );
  OAI22_X1 U49478 ( .A1(n68260), .A2(n62011), .B1(n68253), .B2(n68169), .ZN(
        n7460) );
  OAI22_X1 U49479 ( .A1(n68261), .A2(n62009), .B1(n68253), .B2(n68172), .ZN(
        n7461) );
  OAI22_X1 U49480 ( .A1(n68261), .A2(n62007), .B1(n68253), .B2(n68175), .ZN(
        n7462) );
  OAI22_X1 U49481 ( .A1(n68261), .A2(n62005), .B1(n68253), .B2(n68178), .ZN(
        n7463) );
  OAI22_X1 U49482 ( .A1(n68261), .A2(n62003), .B1(n68253), .B2(n68181), .ZN(
        n7464) );
  OAI22_X1 U49483 ( .A1(n68261), .A2(n62001), .B1(n68253), .B2(n68184), .ZN(
        n7465) );
  OAI22_X1 U49484 ( .A1(n68261), .A2(n61999), .B1(n68253), .B2(n68187), .ZN(
        n7466) );
  OAI22_X1 U49485 ( .A1(n68261), .A2(n61997), .B1(n68253), .B2(n68190), .ZN(
        n7467) );
  OAI22_X1 U49486 ( .A1(n68261), .A2(n61995), .B1(n68253), .B2(n68193), .ZN(
        n7468) );
  OAI22_X1 U49487 ( .A1(n68261), .A2(n61993), .B1(n68253), .B2(n68196), .ZN(
        n7469) );
  OAI22_X1 U49488 ( .A1(n68261), .A2(n61991), .B1(n68253), .B2(n68199), .ZN(
        n7470) );
  OAI22_X1 U49489 ( .A1(n68261), .A2(n61989), .B1(n68254), .B2(n68202), .ZN(
        n7471) );
  OAI22_X1 U49490 ( .A1(n68261), .A2(n61987), .B1(n68254), .B2(n68205), .ZN(
        n7472) );
  OAI22_X1 U49491 ( .A1(n68261), .A2(n61985), .B1(n68254), .B2(n68208), .ZN(
        n7473) );
  OAI22_X1 U49492 ( .A1(n68262), .A2(n61983), .B1(n68254), .B2(n68211), .ZN(
        n7474) );
  OAI22_X1 U49493 ( .A1(n68262), .A2(n61981), .B1(n68254), .B2(n68214), .ZN(
        n7475) );
  OAI22_X1 U49494 ( .A1(n68262), .A2(n61979), .B1(n68254), .B2(n68217), .ZN(
        n7476) );
  OAI22_X1 U49495 ( .A1(n68262), .A2(n61977), .B1(n68254), .B2(n68220), .ZN(
        n7477) );
  OAI22_X1 U49496 ( .A1(n68262), .A2(n61975), .B1(n68254), .B2(n68223), .ZN(
        n7478) );
  OAI22_X1 U49497 ( .A1(n68262), .A2(n61973), .B1(n68254), .B2(n68226), .ZN(
        n7479) );
  OAI22_X1 U49498 ( .A1(n68262), .A2(n61971), .B1(n68254), .B2(n68229), .ZN(
        n7480) );
  OAI22_X1 U49499 ( .A1(n68262), .A2(n61969), .B1(n68254), .B2(n68232), .ZN(
        n7481) );
  OAI22_X1 U49500 ( .A1(n68262), .A2(n61967), .B1(n68254), .B2(n68235), .ZN(
        n7482) );
  OAI22_X1 U49501 ( .A1(n68262), .A2(n61965), .B1(n68255), .B2(n68238), .ZN(
        n7483) );
  OAI22_X1 U49502 ( .A1(n68262), .A2(n61963), .B1(n68255), .B2(n68241), .ZN(
        n7484) );
  OAI22_X1 U49503 ( .A1(n68262), .A2(n61961), .B1(n68255), .B2(n68244), .ZN(
        n7485) );
  OAI22_X1 U49504 ( .A1(n68262), .A2(n61958), .B1(n68255), .B2(n68247), .ZN(
        n7486) );
  AOI22_X1 U49505 ( .A1(n67594), .A2(n66502), .B1(n58427), .B2(n67588), .ZN(
        n64114) );
  AOI22_X1 U49506 ( .A1(n67594), .A2(n66503), .B1(n58428), .B2(n67588), .ZN(
        n64094) );
  AOI22_X1 U49507 ( .A1(n67594), .A2(n66504), .B1(n58429), .B2(n67588), .ZN(
        n64074) );
  AOI22_X1 U49508 ( .A1(n67594), .A2(n66505), .B1(n58430), .B2(n67588), .ZN(
        n64054) );
  AOI22_X1 U49509 ( .A1(n67594), .A2(n66506), .B1(n58431), .B2(n67588), .ZN(
        n64034) );
  AOI22_X1 U49510 ( .A1(n67594), .A2(n66507), .B1(n58432), .B2(n67588), .ZN(
        n64014) );
  AOI22_X1 U49511 ( .A1(n67594), .A2(n66508), .B1(n58433), .B2(n67588), .ZN(
        n63994) );
  AOI22_X1 U49512 ( .A1(n67594), .A2(n66509), .B1(n58434), .B2(n67588), .ZN(
        n63974) );
  AOI22_X1 U49513 ( .A1(n67594), .A2(n66510), .B1(n58435), .B2(n67588), .ZN(
        n63954) );
  AOI22_X1 U49514 ( .A1(n67594), .A2(n66511), .B1(n58436), .B2(n67588), .ZN(
        n63934) );
  AOI22_X1 U49515 ( .A1(n67594), .A2(n66512), .B1(n58437), .B2(n67588), .ZN(
        n63914) );
  AOI22_X1 U49516 ( .A1(n67594), .A2(n66513), .B1(n58438), .B2(n67588), .ZN(
        n63894) );
  OAI22_X1 U49517 ( .A1(n54186), .A2(n67934), .B1(n68238), .B2(n67928), .ZN(
        n6843) );
  OAI22_X1 U49518 ( .A1(n54185), .A2(n67934), .B1(n68241), .B2(n67928), .ZN(
        n6844) );
  OAI22_X1 U49519 ( .A1(n54184), .A2(n67934), .B1(n68244), .B2(n67928), .ZN(
        n6845) );
  OAI22_X1 U49520 ( .A1(n54610), .A2(n67730), .B1(n68240), .B2(n67724), .ZN(
        n5819) );
  OAI22_X1 U49521 ( .A1(n54609), .A2(n67730), .B1(n68243), .B2(n67724), .ZN(
        n5820) );
  OAI22_X1 U49522 ( .A1(n54608), .A2(n67730), .B1(n68246), .B2(n67724), .ZN(
        n5821) );
  OAI22_X1 U49523 ( .A1(n54606), .A2(n67730), .B1(n68249), .B2(n67724), .ZN(
        n5822) );
  OAI22_X1 U49524 ( .A1(n67666), .A2(n63862), .B1(n68240), .B2(n67659), .ZN(
        n5496) );
  OAI22_X1 U49525 ( .A1(n67666), .A2(n63841), .B1(n68243), .B2(n67659), .ZN(
        n5498) );
  OAI22_X1 U49526 ( .A1(n67666), .A2(n63820), .B1(n68246), .B2(n67659), .ZN(
        n5500) );
  OAI22_X1 U49527 ( .A1(n67666), .A2(n63765), .B1(n68249), .B2(n67659), .ZN(
        n5502) );
  OAI22_X1 U49528 ( .A1(n49229), .A2(n67909), .B1(n68239), .B2(n67903), .ZN(
        n6715) );
  OAI22_X1 U49529 ( .A1(n49230), .A2(n67909), .B1(n68242), .B2(n67903), .ZN(
        n6716) );
  OAI22_X1 U49530 ( .A1(n49231), .A2(n67909), .B1(n68245), .B2(n67903), .ZN(
        n6717) );
  OAI22_X1 U49531 ( .A1(n49228), .A2(n67909), .B1(n68248), .B2(n67903), .ZN(
        n6718) );
  OAI22_X1 U49532 ( .A1(n67679), .A2(n63703), .B1(n68240), .B2(n67672), .ZN(
        n5563) );
  OAI22_X1 U49533 ( .A1(n67679), .A2(n63702), .B1(n68243), .B2(n67672), .ZN(
        n5564) );
  OAI22_X1 U49534 ( .A1(n67679), .A2(n63701), .B1(n68246), .B2(n67672), .ZN(
        n5565) );
  OAI22_X1 U49535 ( .A1(n67679), .A2(n63699), .B1(n68249), .B2(n67672), .ZN(
        n5566) );
  OAI22_X1 U49536 ( .A1(n8461), .A2(n67893), .B1(n68239), .B2(n67890), .ZN(
        n6651) );
  OAI22_X1 U49537 ( .A1(n8477), .A2(n67893), .B1(n68242), .B2(n67890), .ZN(
        n6652) );
  OAI22_X1 U49538 ( .A1(n8493), .A2(n67893), .B1(n68245), .B2(n67890), .ZN(
        n6653) );
  OAI22_X1 U49539 ( .A1(n8509), .A2(n67893), .B1(n68248), .B2(n67890), .ZN(
        n6654) );
  OAI22_X1 U49540 ( .A1(n49480), .A2(n67832), .B1(n68239), .B2(n67826), .ZN(
        n6331) );
  OAI22_X1 U49541 ( .A1(n49481), .A2(n67832), .B1(n68242), .B2(n67826), .ZN(
        n6332) );
  OAI22_X1 U49542 ( .A1(n49482), .A2(n67832), .B1(n68245), .B2(n67826), .ZN(
        n6333) );
  OAI22_X1 U49543 ( .A1(n49483), .A2(n67832), .B1(n68248), .B2(n67826), .ZN(
        n6334) );
  OAI22_X1 U49544 ( .A1(n67782), .A2(n63234), .B1(n68239), .B2(n67775), .ZN(
        n6075) );
  OAI22_X1 U49545 ( .A1(n67782), .A2(n63233), .B1(n68242), .B2(n67775), .ZN(
        n6076) );
  OAI22_X1 U49546 ( .A1(n67782), .A2(n63232), .B1(n68245), .B2(n67775), .ZN(
        n6077) );
  OAI22_X1 U49547 ( .A1(n67782), .A2(n63230), .B1(n68248), .B2(n67775), .ZN(
        n6078) );
  OAI22_X1 U49548 ( .A1(n8449), .A2(n67794), .B1(n68239), .B2(n67788), .ZN(
        n6139) );
  OAI22_X1 U49549 ( .A1(n8465), .A2(n67794), .B1(n68242), .B2(n67788), .ZN(
        n6140) );
  OAI22_X1 U49550 ( .A1(n8481), .A2(n67794), .B1(n68245), .B2(n67788), .ZN(
        n6141) );
  OAI22_X1 U49551 ( .A1(n8497), .A2(n67794), .B1(n68248), .B2(n67788), .ZN(
        n6142) );
  AOI22_X1 U49552 ( .A1(n67416), .A2(n66313), .B1(n67410), .B2(n58307), .ZN(
        n66282) );
  AOI22_X1 U49553 ( .A1(n67392), .A2(n58787), .B1(n67386), .B2(n58439), .ZN(
        n66284) );
  AOI22_X1 U49554 ( .A1(n67368), .A2(n58036), .B1(n67362), .B2(n8958), .ZN(
        n66288) );
  AOI22_X1 U49555 ( .A1(n67416), .A2(n66314), .B1(n67410), .B2(n58308), .ZN(
        n66258) );
  AOI22_X1 U49556 ( .A1(n67392), .A2(n58788), .B1(n67386), .B2(n58440), .ZN(
        n66259) );
  AOI22_X1 U49557 ( .A1(n67368), .A2(n58001), .B1(n67362), .B2(n8957), .ZN(
        n66260) );
  AOI22_X1 U49558 ( .A1(n67416), .A2(n66315), .B1(n67410), .B2(n58309), .ZN(
        n66240) );
  AOI22_X1 U49559 ( .A1(n67392), .A2(n58789), .B1(n67386), .B2(n58441), .ZN(
        n66241) );
  AOI22_X1 U49560 ( .A1(n67368), .A2(n57977), .B1(n67362), .B2(n8956), .ZN(
        n66242) );
  AOI22_X1 U49561 ( .A1(n67416), .A2(n66316), .B1(n67410), .B2(n58310), .ZN(
        n66222) );
  AOI22_X1 U49562 ( .A1(n67392), .A2(n58790), .B1(n67386), .B2(n58442), .ZN(
        n66223) );
  AOI22_X1 U49563 ( .A1(n67368), .A2(n57953), .B1(n67362), .B2(n8955), .ZN(
        n66224) );
  AOI22_X1 U49564 ( .A1(n67416), .A2(n66317), .B1(n67410), .B2(n58311), .ZN(
        n66204) );
  AOI22_X1 U49565 ( .A1(n67392), .A2(n58791), .B1(n67386), .B2(n58443), .ZN(
        n66205) );
  AOI22_X1 U49566 ( .A1(n67368), .A2(n57929), .B1(n67362), .B2(n8954), .ZN(
        n66206) );
  AOI22_X1 U49567 ( .A1(n67416), .A2(n66318), .B1(n67410), .B2(n58312), .ZN(
        n66186) );
  AOI22_X1 U49568 ( .A1(n67392), .A2(n58792), .B1(n67386), .B2(n58444), .ZN(
        n66187) );
  AOI22_X1 U49569 ( .A1(n67368), .A2(n57905), .B1(n67362), .B2(n8953), .ZN(
        n66188) );
  AOI22_X1 U49570 ( .A1(n67416), .A2(n66319), .B1(n67410), .B2(n58313), .ZN(
        n66168) );
  AOI22_X1 U49571 ( .A1(n67392), .A2(n58793), .B1(n67386), .B2(n58445), .ZN(
        n66169) );
  AOI22_X1 U49572 ( .A1(n67368), .A2(n57881), .B1(n67362), .B2(n8952), .ZN(
        n66170) );
  AOI22_X1 U49573 ( .A1(n67416), .A2(n66320), .B1(n67410), .B2(n58314), .ZN(
        n66150) );
  AOI22_X1 U49574 ( .A1(n67392), .A2(n58794), .B1(n67386), .B2(n58446), .ZN(
        n66151) );
  AOI22_X1 U49575 ( .A1(n67368), .A2(n57857), .B1(n67362), .B2(n8951), .ZN(
        n66152) );
  AOI22_X1 U49576 ( .A1(n67416), .A2(n66321), .B1(n67410), .B2(n58315), .ZN(
        n66132) );
  AOI22_X1 U49577 ( .A1(n67392), .A2(n58795), .B1(n67386), .B2(n58447), .ZN(
        n66133) );
  AOI22_X1 U49578 ( .A1(n67368), .A2(n57833), .B1(n67362), .B2(n8950), .ZN(
        n66134) );
  AOI22_X1 U49579 ( .A1(n67416), .A2(n66322), .B1(n67410), .B2(n58316), .ZN(
        n66114) );
  AOI22_X1 U49580 ( .A1(n67392), .A2(n58796), .B1(n67386), .B2(n58448), .ZN(
        n66115) );
  AOI22_X1 U49581 ( .A1(n67368), .A2(n57809), .B1(n67362), .B2(n8949), .ZN(
        n66116) );
  AOI22_X1 U49582 ( .A1(n67416), .A2(n66323), .B1(n67410), .B2(n58317), .ZN(
        n66096) );
  AOI22_X1 U49583 ( .A1(n67392), .A2(n58797), .B1(n67386), .B2(n58449), .ZN(
        n66097) );
  AOI22_X1 U49584 ( .A1(n67368), .A2(n57785), .B1(n67362), .B2(n8948), .ZN(
        n66098) );
  AOI22_X1 U49585 ( .A1(n67416), .A2(n66324), .B1(n67410), .B2(n58318), .ZN(
        n66078) );
  AOI22_X1 U49586 ( .A1(n67392), .A2(n58798), .B1(n67386), .B2(n58450), .ZN(
        n66079) );
  AOI22_X1 U49587 ( .A1(n67368), .A2(n57761), .B1(n67362), .B2(n8947), .ZN(
        n66080) );
  AOI22_X1 U49588 ( .A1(n67441), .A2(n58391), .B1(n67435), .B2(OUT2[12]), .ZN(
        n66059) );
  AOI22_X1 U49589 ( .A1(n67393), .A2(n56101), .B1(n67387), .B2(n58451), .ZN(
        n66061) );
  AOI22_X1 U49590 ( .A1(n67369), .A2(n57737), .B1(n67363), .B2(n8946), .ZN(
        n66062) );
  AOI22_X1 U49591 ( .A1(n67441), .A2(n58392), .B1(n67435), .B2(OUT2[13]), .ZN(
        n66041) );
  AOI22_X1 U49592 ( .A1(n67393), .A2(n56074), .B1(n67387), .B2(n58452), .ZN(
        n66043) );
  AOI22_X1 U49593 ( .A1(n67369), .A2(n57713), .B1(n67363), .B2(n8945), .ZN(
        n66044) );
  AOI22_X1 U49594 ( .A1(n67441), .A2(n58393), .B1(n67435), .B2(OUT2[14]), .ZN(
        n66023) );
  AOI22_X1 U49595 ( .A1(n67393), .A2(n56047), .B1(n67387), .B2(n58453), .ZN(
        n66025) );
  AOI22_X1 U49596 ( .A1(n67369), .A2(n57689), .B1(n67363), .B2(n8944), .ZN(
        n66026) );
  AOI22_X1 U49597 ( .A1(n67441), .A2(n58394), .B1(n67435), .B2(OUT2[15]), .ZN(
        n66005) );
  AOI22_X1 U49598 ( .A1(n67393), .A2(n56020), .B1(n67387), .B2(n58454), .ZN(
        n66007) );
  AOI22_X1 U49599 ( .A1(n67369), .A2(n57665), .B1(n67363), .B2(n8943), .ZN(
        n66008) );
  AOI22_X1 U49600 ( .A1(n67441), .A2(n58395), .B1(n67435), .B2(OUT2[16]), .ZN(
        n65987) );
  AOI22_X1 U49601 ( .A1(n67393), .A2(n58799), .B1(n67387), .B2(n58455), .ZN(
        n65989) );
  AOI22_X1 U49602 ( .A1(n67369), .A2(n57641), .B1(n67363), .B2(n8942), .ZN(
        n65990) );
  AOI22_X1 U49603 ( .A1(n67441), .A2(n58396), .B1(n67435), .B2(OUT2[17]), .ZN(
        n65969) );
  AOI22_X1 U49604 ( .A1(n67393), .A2(n58800), .B1(n67387), .B2(n58456), .ZN(
        n65971) );
  AOI22_X1 U49605 ( .A1(n67369), .A2(n57617), .B1(n67363), .B2(n8941), .ZN(
        n65972) );
  AOI22_X1 U49606 ( .A1(n67441), .A2(n58397), .B1(n67435), .B2(OUT2[18]), .ZN(
        n65951) );
  AOI22_X1 U49607 ( .A1(n67393), .A2(n58801), .B1(n67387), .B2(n58457), .ZN(
        n65953) );
  AOI22_X1 U49608 ( .A1(n67369), .A2(n57593), .B1(n67363), .B2(n8940), .ZN(
        n65954) );
  AOI22_X1 U49609 ( .A1(n67441), .A2(n58398), .B1(n67435), .B2(OUT2[19]), .ZN(
        n65933) );
  AOI22_X1 U49610 ( .A1(n67393), .A2(n58802), .B1(n67387), .B2(n58458), .ZN(
        n65935) );
  AOI22_X1 U49611 ( .A1(n67369), .A2(n57569), .B1(n67363), .B2(n8939), .ZN(
        n65936) );
  AOI22_X1 U49612 ( .A1(n67441), .A2(n58399), .B1(n67435), .B2(OUT2[20]), .ZN(
        n65915) );
  AOI22_X1 U49613 ( .A1(n67393), .A2(n58803), .B1(n67387), .B2(n58459), .ZN(
        n65917) );
  AOI22_X1 U49614 ( .A1(n67369), .A2(n57545), .B1(n67363), .B2(n8938), .ZN(
        n65918) );
  AOI22_X1 U49615 ( .A1(n67441), .A2(n58400), .B1(n67435), .B2(OUT2[21]), .ZN(
        n65897) );
  AOI22_X1 U49616 ( .A1(n67393), .A2(n58804), .B1(n67387), .B2(n58460), .ZN(
        n65899) );
  AOI22_X1 U49617 ( .A1(n67369), .A2(n57521), .B1(n67363), .B2(n8937), .ZN(
        n65900) );
  AOI22_X1 U49618 ( .A1(n67441), .A2(n58401), .B1(n67436), .B2(OUT2[22]), .ZN(
        n65879) );
  AOI22_X1 U49619 ( .A1(n67393), .A2(n58805), .B1(n67387), .B2(n58461), .ZN(
        n65881) );
  AOI22_X1 U49620 ( .A1(n67369), .A2(n57497), .B1(n67363), .B2(n8936), .ZN(
        n65882) );
  AOI22_X1 U49621 ( .A1(n67441), .A2(n58402), .B1(n67436), .B2(OUT2[23]), .ZN(
        n65861) );
  AOI22_X1 U49622 ( .A1(n67393), .A2(n58806), .B1(n67387), .B2(n58462), .ZN(
        n65863) );
  AOI22_X1 U49623 ( .A1(n67369), .A2(n57473), .B1(n67363), .B2(n8935), .ZN(
        n65864) );
  AOI22_X1 U49624 ( .A1(n67442), .A2(n58403), .B1(n67436), .B2(OUT2[24]), .ZN(
        n65843) );
  AOI22_X1 U49625 ( .A1(n67394), .A2(n58807), .B1(n67388), .B2(n58463), .ZN(
        n65845) );
  AOI22_X1 U49626 ( .A1(n67370), .A2(n57449), .B1(n67364), .B2(n8934), .ZN(
        n65846) );
  AOI22_X1 U49627 ( .A1(n67442), .A2(n58404), .B1(n67436), .B2(OUT2[25]), .ZN(
        n65825) );
  AOI22_X1 U49628 ( .A1(n67394), .A2(n58808), .B1(n67388), .B2(n58464), .ZN(
        n65827) );
  AOI22_X1 U49629 ( .A1(n67370), .A2(n57425), .B1(n67364), .B2(n8933), .ZN(
        n65828) );
  AOI22_X1 U49630 ( .A1(n67442), .A2(n58405), .B1(n67436), .B2(OUT2[26]), .ZN(
        n65807) );
  AOI22_X1 U49631 ( .A1(n67394), .A2(n58809), .B1(n67388), .B2(n58465), .ZN(
        n65809) );
  AOI22_X1 U49632 ( .A1(n67370), .A2(n57401), .B1(n67364), .B2(n8932), .ZN(
        n65810) );
  AOI22_X1 U49633 ( .A1(n67442), .A2(n58406), .B1(n67436), .B2(OUT2[27]), .ZN(
        n65789) );
  AOI22_X1 U49634 ( .A1(n67394), .A2(n58810), .B1(n67388), .B2(n58466), .ZN(
        n65791) );
  AOI22_X1 U49635 ( .A1(n67370), .A2(n57377), .B1(n67364), .B2(n8931), .ZN(
        n65792) );
  AOI22_X1 U49636 ( .A1(n67442), .A2(n58407), .B1(n67436), .B2(OUT2[28]), .ZN(
        n65771) );
  AOI22_X1 U49637 ( .A1(n67394), .A2(n58811), .B1(n67388), .B2(n58467), .ZN(
        n65773) );
  AOI22_X1 U49638 ( .A1(n67370), .A2(n57353), .B1(n67364), .B2(n8930), .ZN(
        n65774) );
  AOI22_X1 U49639 ( .A1(n67442), .A2(n58408), .B1(n67436), .B2(OUT2[29]), .ZN(
        n65753) );
  AOI22_X1 U49640 ( .A1(n67394), .A2(n58812), .B1(n67388), .B2(n58468), .ZN(
        n65755) );
  AOI22_X1 U49641 ( .A1(n67370), .A2(n57329), .B1(n67364), .B2(n8929), .ZN(
        n65756) );
  AOI22_X1 U49642 ( .A1(n67442), .A2(n58409), .B1(n67436), .B2(OUT2[30]), .ZN(
        n65735) );
  AOI22_X1 U49643 ( .A1(n67394), .A2(n58813), .B1(n67388), .B2(n58469), .ZN(
        n65737) );
  AOI22_X1 U49644 ( .A1(n67370), .A2(n57305), .B1(n67364), .B2(n8928), .ZN(
        n65738) );
  AOI22_X1 U49645 ( .A1(n67442), .A2(n58410), .B1(n67436), .B2(OUT2[31]), .ZN(
        n65717) );
  AOI22_X1 U49646 ( .A1(n67394), .A2(n58814), .B1(n67388), .B2(n58470), .ZN(
        n65719) );
  AOI22_X1 U49647 ( .A1(n67370), .A2(n57281), .B1(n67364), .B2(n8927), .ZN(
        n65720) );
  AOI22_X1 U49648 ( .A1(n67442), .A2(n58411), .B1(n67436), .B2(OUT2[32]), .ZN(
        n65699) );
  AOI22_X1 U49649 ( .A1(n67394), .A2(n58815), .B1(n67388), .B2(n58471), .ZN(
        n65701) );
  AOI22_X1 U49650 ( .A1(n67370), .A2(n57257), .B1(n67364), .B2(n8926), .ZN(
        n65702) );
  AOI22_X1 U49651 ( .A1(n67442), .A2(n58412), .B1(n67436), .B2(OUT2[33]), .ZN(
        n65681) );
  AOI22_X1 U49652 ( .A1(n67394), .A2(n58816), .B1(n67388), .B2(n58472), .ZN(
        n65683) );
  AOI22_X1 U49653 ( .A1(n67370), .A2(n57233), .B1(n67364), .B2(n8925), .ZN(
        n65684) );
  AOI22_X1 U49654 ( .A1(n67442), .A2(n58413), .B1(n67436), .B2(OUT2[34]), .ZN(
        n65663) );
  AOI22_X1 U49655 ( .A1(n67394), .A2(n58817), .B1(n67388), .B2(n58473), .ZN(
        n65665) );
  AOI22_X1 U49656 ( .A1(n67370), .A2(n57209), .B1(n67364), .B2(n8924), .ZN(
        n65666) );
  AOI22_X1 U49657 ( .A1(n67442), .A2(n58414), .B1(n67437), .B2(OUT2[35]), .ZN(
        n65645) );
  AOI22_X1 U49658 ( .A1(n67394), .A2(n58818), .B1(n67388), .B2(n58474), .ZN(
        n65647) );
  AOI22_X1 U49659 ( .A1(n67370), .A2(n57185), .B1(n67364), .B2(n8923), .ZN(
        n65648) );
  AOI22_X1 U49660 ( .A1(n67443), .A2(n58415), .B1(n67437), .B2(OUT2[36]), .ZN(
        n65627) );
  AOI22_X1 U49661 ( .A1(n67395), .A2(n58819), .B1(n67389), .B2(n58475), .ZN(
        n65629) );
  AOI22_X1 U49662 ( .A1(n67371), .A2(n57161), .B1(n67365), .B2(n8922), .ZN(
        n65630) );
  AOI22_X1 U49663 ( .A1(n67443), .A2(n58416), .B1(n67437), .B2(OUT2[37]), .ZN(
        n65609) );
  AOI22_X1 U49664 ( .A1(n67395), .A2(n58820), .B1(n67389), .B2(n58476), .ZN(
        n65611) );
  AOI22_X1 U49665 ( .A1(n67371), .A2(n57137), .B1(n67365), .B2(n8921), .ZN(
        n65612) );
  AOI22_X1 U49666 ( .A1(n67443), .A2(n58417), .B1(n67437), .B2(OUT2[38]), .ZN(
        n65591) );
  AOI22_X1 U49667 ( .A1(n67395), .A2(n58821), .B1(n67389), .B2(n58477), .ZN(
        n65593) );
  AOI22_X1 U49668 ( .A1(n67371), .A2(n57113), .B1(n67365), .B2(n8920), .ZN(
        n65594) );
  AOI22_X1 U49669 ( .A1(n67443), .A2(n58418), .B1(n67437), .B2(OUT2[39]), .ZN(
        n65573) );
  AOI22_X1 U49670 ( .A1(n67395), .A2(n58822), .B1(n67389), .B2(n58478), .ZN(
        n65575) );
  AOI22_X1 U49671 ( .A1(n67371), .A2(n57089), .B1(n67365), .B2(n8919), .ZN(
        n65576) );
  AOI22_X1 U49672 ( .A1(n67443), .A2(n58419), .B1(n67437), .B2(OUT2[40]), .ZN(
        n65555) );
  AOI22_X1 U49673 ( .A1(n67395), .A2(n58823), .B1(n67389), .B2(n58479), .ZN(
        n65557) );
  AOI22_X1 U49674 ( .A1(n67371), .A2(n57065), .B1(n67365), .B2(n8918), .ZN(
        n65558) );
  AOI22_X1 U49675 ( .A1(n67443), .A2(n58420), .B1(n67437), .B2(OUT2[41]), .ZN(
        n65537) );
  AOI22_X1 U49676 ( .A1(n67395), .A2(n58824), .B1(n67389), .B2(n58480), .ZN(
        n65539) );
  AOI22_X1 U49677 ( .A1(n67371), .A2(n57041), .B1(n67365), .B2(n8917), .ZN(
        n65540) );
  AOI22_X1 U49678 ( .A1(n67443), .A2(n58421), .B1(n67437), .B2(OUT2[42]), .ZN(
        n65519) );
  AOI22_X1 U49679 ( .A1(n67395), .A2(n58825), .B1(n67389), .B2(n58481), .ZN(
        n65521) );
  AOI22_X1 U49680 ( .A1(n67371), .A2(n57017), .B1(n67365), .B2(n8916), .ZN(
        n65522) );
  AOI22_X1 U49681 ( .A1(n67443), .A2(n58422), .B1(n67437), .B2(OUT2[43]), .ZN(
        n65501) );
  AOI22_X1 U49682 ( .A1(n67395), .A2(n58826), .B1(n67389), .B2(n58482), .ZN(
        n65503) );
  AOI22_X1 U49683 ( .A1(n67371), .A2(n56993), .B1(n67365), .B2(n8915), .ZN(
        n65504) );
  AOI22_X1 U49684 ( .A1(n67443), .A2(n58423), .B1(n67437), .B2(OUT2[44]), .ZN(
        n65483) );
  AOI22_X1 U49685 ( .A1(n67395), .A2(n58827), .B1(n67389), .B2(n58483), .ZN(
        n65485) );
  AOI22_X1 U49686 ( .A1(n67371), .A2(n56969), .B1(n67365), .B2(n8914), .ZN(
        n65486) );
  AOI22_X1 U49687 ( .A1(n67443), .A2(n58424), .B1(n67437), .B2(OUT2[45]), .ZN(
        n65465) );
  AOI22_X1 U49688 ( .A1(n67395), .A2(n58828), .B1(n67389), .B2(n58484), .ZN(
        n65467) );
  AOI22_X1 U49689 ( .A1(n67371), .A2(n56945), .B1(n67365), .B2(n8913), .ZN(
        n65468) );
  AOI22_X1 U49690 ( .A1(n67443), .A2(n58425), .B1(n67437), .B2(OUT2[46]), .ZN(
        n65447) );
  AOI22_X1 U49691 ( .A1(n67395), .A2(n58829), .B1(n67389), .B2(n58485), .ZN(
        n65449) );
  AOI22_X1 U49692 ( .A1(n67371), .A2(n56921), .B1(n67365), .B2(n8912), .ZN(
        n65450) );
  AOI22_X1 U49693 ( .A1(n67443), .A2(n58426), .B1(n67437), .B2(OUT2[47]), .ZN(
        n65429) );
  AOI22_X1 U49694 ( .A1(n67395), .A2(n58830), .B1(n67389), .B2(n58486), .ZN(
        n65431) );
  AOI22_X1 U49695 ( .A1(n67371), .A2(n56897), .B1(n67365), .B2(n8911), .ZN(
        n65432) );
  AOI22_X1 U49696 ( .A1(n67444), .A2(n58427), .B1(n67438), .B2(OUT2[48]), .ZN(
        n65411) );
  AOI22_X1 U49697 ( .A1(n67396), .A2(n58831), .B1(n67390), .B2(n58487), .ZN(
        n65413) );
  AOI22_X1 U49698 ( .A1(n67372), .A2(n56873), .B1(n67366), .B2(n8910), .ZN(
        n65414) );
  AOI22_X1 U49699 ( .A1(n67444), .A2(n58428), .B1(n67438), .B2(OUT2[49]), .ZN(
        n65393) );
  AOI22_X1 U49700 ( .A1(n67396), .A2(n58832), .B1(n67390), .B2(n58488), .ZN(
        n65395) );
  AOI22_X1 U49701 ( .A1(n67372), .A2(n56849), .B1(n67366), .B2(n8909), .ZN(
        n65396) );
  AOI22_X1 U49702 ( .A1(n67444), .A2(n58429), .B1(n67438), .B2(OUT2[50]), .ZN(
        n65375) );
  AOI22_X1 U49703 ( .A1(n67396), .A2(n58833), .B1(n67390), .B2(n58489), .ZN(
        n65377) );
  AOI22_X1 U49704 ( .A1(n67372), .A2(n56825), .B1(n67366), .B2(n8908), .ZN(
        n65378) );
  AOI22_X1 U49705 ( .A1(n67444), .A2(n58430), .B1(n67438), .B2(OUT2[51]), .ZN(
        n65357) );
  AOI22_X1 U49706 ( .A1(n67396), .A2(n58834), .B1(n67390), .B2(n58490), .ZN(
        n65359) );
  AOI22_X1 U49707 ( .A1(n67372), .A2(n56801), .B1(n67366), .B2(n8907), .ZN(
        n65360) );
  AOI22_X1 U49708 ( .A1(n67444), .A2(n58431), .B1(n67438), .B2(OUT2[52]), .ZN(
        n65339) );
  AOI22_X1 U49709 ( .A1(n67396), .A2(n58835), .B1(n67390), .B2(n58491), .ZN(
        n65341) );
  AOI22_X1 U49710 ( .A1(n67372), .A2(n56777), .B1(n67366), .B2(n8906), .ZN(
        n65342) );
  AOI22_X1 U49711 ( .A1(n67444), .A2(n58432), .B1(n67438), .B2(OUT2[53]), .ZN(
        n65321) );
  AOI22_X1 U49712 ( .A1(n67396), .A2(n58836), .B1(n67390), .B2(n58492), .ZN(
        n65323) );
  AOI22_X1 U49713 ( .A1(n67372), .A2(n56753), .B1(n67366), .B2(n8905), .ZN(
        n65324) );
  AOI22_X1 U49714 ( .A1(n67444), .A2(n58433), .B1(n67438), .B2(OUT2[54]), .ZN(
        n65303) );
  AOI22_X1 U49715 ( .A1(n67396), .A2(n58837), .B1(n67390), .B2(n58493), .ZN(
        n65305) );
  AOI22_X1 U49716 ( .A1(n67372), .A2(n56729), .B1(n67366), .B2(n8904), .ZN(
        n65306) );
  AOI22_X1 U49717 ( .A1(n67444), .A2(n58434), .B1(n67438), .B2(OUT2[55]), .ZN(
        n65285) );
  AOI22_X1 U49718 ( .A1(n67396), .A2(n58838), .B1(n67390), .B2(n58494), .ZN(
        n65287) );
  AOI22_X1 U49719 ( .A1(n67372), .A2(n56705), .B1(n67366), .B2(n8903), .ZN(
        n65288) );
  AOI22_X1 U49720 ( .A1(n67444), .A2(n58435), .B1(n67438), .B2(OUT2[56]), .ZN(
        n65267) );
  AOI22_X1 U49721 ( .A1(n67396), .A2(n58839), .B1(n67390), .B2(n58495), .ZN(
        n65269) );
  AOI22_X1 U49722 ( .A1(n67372), .A2(n56681), .B1(n67366), .B2(n8902), .ZN(
        n65270) );
  AOI22_X1 U49723 ( .A1(n67444), .A2(n58436), .B1(n67438), .B2(OUT2[57]), .ZN(
        n65249) );
  AOI22_X1 U49724 ( .A1(n67396), .A2(n58840), .B1(n67390), .B2(n58496), .ZN(
        n65251) );
  AOI22_X1 U49725 ( .A1(n67372), .A2(n56657), .B1(n67366), .B2(n8901), .ZN(
        n65252) );
  AOI22_X1 U49726 ( .A1(n67444), .A2(n58437), .B1(n67438), .B2(OUT2[58]), .ZN(
        n65231) );
  AOI22_X1 U49727 ( .A1(n67396), .A2(n58841), .B1(n67390), .B2(n58497), .ZN(
        n65233) );
  AOI22_X1 U49728 ( .A1(n67372), .A2(n56633), .B1(n67366), .B2(n8900), .ZN(
        n65234) );
  AOI22_X1 U49729 ( .A1(n67444), .A2(n58438), .B1(n67438), .B2(OUT2[59]), .ZN(
        n65213) );
  AOI22_X1 U49730 ( .A1(n67396), .A2(n58842), .B1(n67390), .B2(n58498), .ZN(
        n65215) );
  AOI22_X1 U49731 ( .A1(n67372), .A2(n56609), .B1(n67366), .B2(n8899), .ZN(
        n65216) );
  AOI22_X1 U49732 ( .A1(n67590), .A2(n65084), .B1(n58379), .B2(n67584), .ZN(
        n65083) );
  AOI22_X1 U49733 ( .A1(n67636), .A2(n58013), .B1(n67632), .B2(OUT1[0]), .ZN(
        n65072) );
  AOI22_X1 U49734 ( .A1(n67614), .A2(n58627), .B1(n67608), .B2(n58731), .ZN(
        n65079) );
  AOI22_X1 U49735 ( .A1(n67590), .A2(n65055), .B1(n58380), .B2(n67584), .ZN(
        n65054) );
  AOI22_X1 U49736 ( .A1(n67636), .A2(n57989), .B1(n67632), .B2(OUT1[1]), .ZN(
        n65052) );
  AOI22_X1 U49737 ( .A1(n67614), .A2(n58628), .B1(n67608), .B2(n58732), .ZN(
        n65053) );
  AOI22_X1 U49738 ( .A1(n67590), .A2(n65035), .B1(n58381), .B2(n67584), .ZN(
        n65034) );
  AOI22_X1 U49739 ( .A1(n67636), .A2(n57965), .B1(n67632), .B2(OUT1[2]), .ZN(
        n65032) );
  AOI22_X1 U49740 ( .A1(n67614), .A2(n58629), .B1(n67608), .B2(n58733), .ZN(
        n65033) );
  AOI22_X1 U49741 ( .A1(n67590), .A2(n65015), .B1(n58382), .B2(n67584), .ZN(
        n65014) );
  AOI22_X1 U49742 ( .A1(n67636), .A2(n57941), .B1(n67632), .B2(OUT1[3]), .ZN(
        n65012) );
  AOI22_X1 U49743 ( .A1(n67614), .A2(n58630), .B1(n67608), .B2(n58734), .ZN(
        n65013) );
  AOI22_X1 U49744 ( .A1(n67590), .A2(n64995), .B1(n58383), .B2(n67584), .ZN(
        n64994) );
  AOI22_X1 U49745 ( .A1(n67636), .A2(n57917), .B1(n67632), .B2(OUT1[4]), .ZN(
        n64992) );
  AOI22_X1 U49746 ( .A1(n67614), .A2(n58631), .B1(n67608), .B2(n58735), .ZN(
        n64993) );
  AOI22_X1 U49747 ( .A1(n67590), .A2(n64975), .B1(n58384), .B2(n67584), .ZN(
        n64974) );
  AOI22_X1 U49748 ( .A1(n67636), .A2(n57893), .B1(n67632), .B2(OUT1[5]), .ZN(
        n64972) );
  AOI22_X1 U49749 ( .A1(n67614), .A2(n58632), .B1(n67608), .B2(n58736), .ZN(
        n64973) );
  AOI22_X1 U49750 ( .A1(n67590), .A2(n64955), .B1(n58385), .B2(n67584), .ZN(
        n64954) );
  AOI22_X1 U49751 ( .A1(n67636), .A2(n57869), .B1(n67632), .B2(OUT1[6]), .ZN(
        n64952) );
  AOI22_X1 U49752 ( .A1(n67614), .A2(n58633), .B1(n67608), .B2(n58737), .ZN(
        n64953) );
  AOI22_X1 U49753 ( .A1(n67590), .A2(n64935), .B1(n58386), .B2(n67584), .ZN(
        n64934) );
  AOI22_X1 U49754 ( .A1(n67636), .A2(n57845), .B1(n67632), .B2(OUT1[7]), .ZN(
        n64932) );
  AOI22_X1 U49755 ( .A1(n67614), .A2(n58634), .B1(n67608), .B2(n58738), .ZN(
        n64933) );
  AOI22_X1 U49756 ( .A1(n67590), .A2(n64915), .B1(n58387), .B2(n67584), .ZN(
        n64914) );
  AOI22_X1 U49757 ( .A1(n67636), .A2(n57821), .B1(n67632), .B2(OUT1[8]), .ZN(
        n64912) );
  AOI22_X1 U49758 ( .A1(n67614), .A2(n58635), .B1(n67608), .B2(n58739), .ZN(
        n64913) );
  AOI22_X1 U49759 ( .A1(n67590), .A2(n64895), .B1(n58388), .B2(n67584), .ZN(
        n64894) );
  AOI22_X1 U49760 ( .A1(n67636), .A2(n57797), .B1(n67632), .B2(OUT1[9]), .ZN(
        n64892) );
  AOI22_X1 U49761 ( .A1(n67614), .A2(n58636), .B1(n67608), .B2(n58740), .ZN(
        n64893) );
  AOI22_X1 U49762 ( .A1(n67590), .A2(n64875), .B1(n58389), .B2(n67584), .ZN(
        n64874) );
  AOI22_X1 U49763 ( .A1(n67636), .A2(n57773), .B1(n67632), .B2(OUT1[10]), .ZN(
        n64872) );
  AOI22_X1 U49764 ( .A1(n67614), .A2(n58637), .B1(n67608), .B2(n58741), .ZN(
        n64873) );
  AOI22_X1 U49765 ( .A1(n67590), .A2(n64855), .B1(n58390), .B2(n67584), .ZN(
        n64854) );
  AOI22_X1 U49766 ( .A1(n67636), .A2(n57749), .B1(n67634), .B2(OUT1[11]), .ZN(
        n64852) );
  AOI22_X1 U49767 ( .A1(n67614), .A2(n58638), .B1(n67608), .B2(n58742), .ZN(
        n64853) );
  AOI22_X1 U49768 ( .A1(n67567), .A2(n9061), .B1(n67561), .B2(n57737), .ZN(
        n64836) );
  AOI22_X1 U49769 ( .A1(n67591), .A2(n66514), .B1(n58391), .B2(n67585), .ZN(
        n64834) );
  AOI22_X1 U49770 ( .A1(n67615), .A2(n58639), .B1(n67609), .B2(n58667), .ZN(
        n64833) );
  AOI22_X1 U49771 ( .A1(n67567), .A2(n9059), .B1(n67561), .B2(n57713), .ZN(
        n64816) );
  AOI22_X1 U49772 ( .A1(n67591), .A2(n66515), .B1(n58392), .B2(n67585), .ZN(
        n64814) );
  AOI22_X1 U49773 ( .A1(n67615), .A2(n58640), .B1(n67609), .B2(n58668), .ZN(
        n64813) );
  AOI22_X1 U49774 ( .A1(n67567), .A2(n9057), .B1(n67561), .B2(n57689), .ZN(
        n64796) );
  AOI22_X1 U49775 ( .A1(n67591), .A2(n66516), .B1(n58393), .B2(n67585), .ZN(
        n64794) );
  AOI22_X1 U49776 ( .A1(n67615), .A2(n58641), .B1(n67609), .B2(n58669), .ZN(
        n64793) );
  AOI22_X1 U49777 ( .A1(n67567), .A2(n9055), .B1(n67561), .B2(n57665), .ZN(
        n64776) );
  AOI22_X1 U49778 ( .A1(n67591), .A2(n66517), .B1(n58394), .B2(n67585), .ZN(
        n64774) );
  AOI22_X1 U49779 ( .A1(n67615), .A2(n58642), .B1(n67609), .B2(n58670), .ZN(
        n64773) );
  AOI22_X1 U49780 ( .A1(n67567), .A2(n9053), .B1(n67561), .B2(n57641), .ZN(
        n64756) );
  AOI22_X1 U49781 ( .A1(n67591), .A2(n66518), .B1(n58395), .B2(n67585), .ZN(
        n64754) );
  AOI22_X1 U49782 ( .A1(n67615), .A2(n57631), .B1(n67609), .B2(n58671), .ZN(
        n64753) );
  AOI22_X1 U49783 ( .A1(n67567), .A2(n9051), .B1(n67561), .B2(n57617), .ZN(
        n64736) );
  AOI22_X1 U49784 ( .A1(n67591), .A2(n66519), .B1(n58396), .B2(n67585), .ZN(
        n64734) );
  AOI22_X1 U49785 ( .A1(n67615), .A2(n57607), .B1(n67609), .B2(n58672), .ZN(
        n64733) );
  AOI22_X1 U49786 ( .A1(n67567), .A2(n9049), .B1(n67561), .B2(n57593), .ZN(
        n64716) );
  AOI22_X1 U49787 ( .A1(n67591), .A2(n66520), .B1(n58397), .B2(n67585), .ZN(
        n64714) );
  AOI22_X1 U49788 ( .A1(n67615), .A2(n57583), .B1(n67609), .B2(n58673), .ZN(
        n64713) );
  AOI22_X1 U49789 ( .A1(n67567), .A2(n9047), .B1(n67561), .B2(n57569), .ZN(
        n64696) );
  AOI22_X1 U49790 ( .A1(n67591), .A2(n66521), .B1(n58398), .B2(n67585), .ZN(
        n64694) );
  AOI22_X1 U49791 ( .A1(n67615), .A2(n57559), .B1(n67609), .B2(n58674), .ZN(
        n64693) );
  AOI22_X1 U49792 ( .A1(n67567), .A2(n9045), .B1(n67561), .B2(n57545), .ZN(
        n64676) );
  AOI22_X1 U49793 ( .A1(n67591), .A2(n66522), .B1(n58399), .B2(n67585), .ZN(
        n64674) );
  AOI22_X1 U49794 ( .A1(n67615), .A2(n57535), .B1(n67609), .B2(n58675), .ZN(
        n64673) );
  AOI22_X1 U49795 ( .A1(n67567), .A2(n9043), .B1(n67561), .B2(n57521), .ZN(
        n64656) );
  AOI22_X1 U49796 ( .A1(n67591), .A2(n66523), .B1(n58400), .B2(n67585), .ZN(
        n64654) );
  AOI22_X1 U49797 ( .A1(n67615), .A2(n57511), .B1(n67609), .B2(n58676), .ZN(
        n64653) );
  AOI22_X1 U49798 ( .A1(n67567), .A2(n9041), .B1(n67561), .B2(n57497), .ZN(
        n64636) );
  AOI22_X1 U49799 ( .A1(n67591), .A2(n66524), .B1(n58401), .B2(n67585), .ZN(
        n64634) );
  AOI22_X1 U49800 ( .A1(n67615), .A2(n57487), .B1(n67609), .B2(n58677), .ZN(
        n64633) );
  AOI22_X1 U49801 ( .A1(n67567), .A2(n9039), .B1(n67561), .B2(n57473), .ZN(
        n64616) );
  AOI22_X1 U49802 ( .A1(n67591), .A2(n66525), .B1(n58402), .B2(n67585), .ZN(
        n64614) );
  AOI22_X1 U49803 ( .A1(n67615), .A2(n57463), .B1(n67609), .B2(n58678), .ZN(
        n64613) );
  AOI22_X1 U49804 ( .A1(n67568), .A2(n9037), .B1(n67562), .B2(n57449), .ZN(
        n64596) );
  AOI22_X1 U49805 ( .A1(n67592), .A2(n66526), .B1(n58403), .B2(n67586), .ZN(
        n64594) );
  AOI22_X1 U49806 ( .A1(n67616), .A2(n57439), .B1(n67610), .B2(n58679), .ZN(
        n64593) );
  AOI22_X1 U49807 ( .A1(n67568), .A2(n9035), .B1(n67562), .B2(n57425), .ZN(
        n64576) );
  AOI22_X1 U49808 ( .A1(n67592), .A2(n66527), .B1(n58404), .B2(n67586), .ZN(
        n64574) );
  AOI22_X1 U49809 ( .A1(n67616), .A2(n57415), .B1(n67610), .B2(n58680), .ZN(
        n64573) );
  AOI22_X1 U49810 ( .A1(n67568), .A2(n9033), .B1(n67562), .B2(n57401), .ZN(
        n64556) );
  AOI22_X1 U49811 ( .A1(n67592), .A2(n66528), .B1(n58405), .B2(n67586), .ZN(
        n64554) );
  AOI22_X1 U49812 ( .A1(n67616), .A2(n57391), .B1(n67610), .B2(n58681), .ZN(
        n64553) );
  AOI22_X1 U49813 ( .A1(n67568), .A2(n9031), .B1(n67562), .B2(n57377), .ZN(
        n64536) );
  AOI22_X1 U49814 ( .A1(n67592), .A2(n66529), .B1(n58406), .B2(n67586), .ZN(
        n64534) );
  AOI22_X1 U49815 ( .A1(n67616), .A2(n57367), .B1(n67610), .B2(n58682), .ZN(
        n64533) );
  AOI22_X1 U49816 ( .A1(n67568), .A2(n9029), .B1(n67562), .B2(n57353), .ZN(
        n64516) );
  AOI22_X1 U49817 ( .A1(n67592), .A2(n66530), .B1(n58407), .B2(n67586), .ZN(
        n64514) );
  AOI22_X1 U49818 ( .A1(n67616), .A2(n57343), .B1(n67610), .B2(n58683), .ZN(
        n64513) );
  AOI22_X1 U49819 ( .A1(n67568), .A2(n9027), .B1(n67562), .B2(n57329), .ZN(
        n64496) );
  AOI22_X1 U49820 ( .A1(n67592), .A2(n66531), .B1(n58408), .B2(n67586), .ZN(
        n64494) );
  AOI22_X1 U49821 ( .A1(n67616), .A2(n57319), .B1(n67610), .B2(n58684), .ZN(
        n64493) );
  AOI22_X1 U49822 ( .A1(n67568), .A2(n9025), .B1(n67562), .B2(n57305), .ZN(
        n64476) );
  AOI22_X1 U49823 ( .A1(n67592), .A2(n66532), .B1(n58409), .B2(n67586), .ZN(
        n64474) );
  AOI22_X1 U49824 ( .A1(n67616), .A2(n57295), .B1(n67610), .B2(n58685), .ZN(
        n64473) );
  AOI22_X1 U49825 ( .A1(n67568), .A2(n9023), .B1(n67562), .B2(n57281), .ZN(
        n64456) );
  AOI22_X1 U49826 ( .A1(n67592), .A2(n66533), .B1(n58410), .B2(n67586), .ZN(
        n64454) );
  AOI22_X1 U49827 ( .A1(n67616), .A2(n57271), .B1(n67610), .B2(n58686), .ZN(
        n64453) );
  AOI22_X1 U49828 ( .A1(n67568), .A2(n9021), .B1(n67562), .B2(n57257), .ZN(
        n64436) );
  AOI22_X1 U49829 ( .A1(n67592), .A2(n66534), .B1(n58411), .B2(n67586), .ZN(
        n64434) );
  AOI22_X1 U49830 ( .A1(n67616), .A2(n57247), .B1(n67610), .B2(n58687), .ZN(
        n64433) );
  AOI22_X1 U49831 ( .A1(n67568), .A2(n9019), .B1(n67562), .B2(n57233), .ZN(
        n64416) );
  AOI22_X1 U49832 ( .A1(n67592), .A2(n66535), .B1(n58412), .B2(n67586), .ZN(
        n64414) );
  AOI22_X1 U49833 ( .A1(n67616), .A2(n57223), .B1(n67610), .B2(n58688), .ZN(
        n64413) );
  AOI22_X1 U49834 ( .A1(n67568), .A2(n9017), .B1(n67562), .B2(n57209), .ZN(
        n64396) );
  AOI22_X1 U49835 ( .A1(n67592), .A2(n66536), .B1(n58413), .B2(n67586), .ZN(
        n64394) );
  AOI22_X1 U49836 ( .A1(n67616), .A2(n57199), .B1(n67610), .B2(n58689), .ZN(
        n64393) );
  AOI22_X1 U49837 ( .A1(n67568), .A2(n9015), .B1(n67562), .B2(n57185), .ZN(
        n64376) );
  AOI22_X1 U49838 ( .A1(n67592), .A2(n66537), .B1(n58414), .B2(n67586), .ZN(
        n64374) );
  AOI22_X1 U49839 ( .A1(n67616), .A2(n57175), .B1(n67610), .B2(n58690), .ZN(
        n64373) );
  AOI22_X1 U49840 ( .A1(n67569), .A2(n9013), .B1(n67563), .B2(n57161), .ZN(
        n64356) );
  AOI22_X1 U49841 ( .A1(n67593), .A2(n66538), .B1(n58415), .B2(n67587), .ZN(
        n64354) );
  AOI22_X1 U49842 ( .A1(n67617), .A2(n57151), .B1(n67611), .B2(n58691), .ZN(
        n64353) );
  AOI22_X1 U49843 ( .A1(n67569), .A2(n9011), .B1(n67563), .B2(n57137), .ZN(
        n64336) );
  AOI22_X1 U49844 ( .A1(n67593), .A2(n66539), .B1(n58416), .B2(n67587), .ZN(
        n64334) );
  AOI22_X1 U49845 ( .A1(n67617), .A2(n57127), .B1(n67611), .B2(n58692), .ZN(
        n64333) );
  AOI22_X1 U49846 ( .A1(n67569), .A2(n9009), .B1(n67563), .B2(n57113), .ZN(
        n64316) );
  AOI22_X1 U49847 ( .A1(n67593), .A2(n66540), .B1(n58417), .B2(n67587), .ZN(
        n64314) );
  AOI22_X1 U49848 ( .A1(n67617), .A2(n57103), .B1(n67611), .B2(n58693), .ZN(
        n64313) );
  AOI22_X1 U49849 ( .A1(n67569), .A2(n9007), .B1(n67563), .B2(n57089), .ZN(
        n64296) );
  AOI22_X1 U49850 ( .A1(n67593), .A2(n66541), .B1(n58418), .B2(n67587), .ZN(
        n64294) );
  AOI22_X1 U49851 ( .A1(n67617), .A2(n57079), .B1(n67611), .B2(n58694), .ZN(
        n64293) );
  AOI22_X1 U49852 ( .A1(n67569), .A2(n9005), .B1(n67563), .B2(n57065), .ZN(
        n64276) );
  AOI22_X1 U49853 ( .A1(n67593), .A2(n66542), .B1(n58419), .B2(n67587), .ZN(
        n64274) );
  AOI22_X1 U49854 ( .A1(n67617), .A2(n57055), .B1(n67611), .B2(n58695), .ZN(
        n64273) );
  AOI22_X1 U49855 ( .A1(n67569), .A2(n9003), .B1(n67563), .B2(n57041), .ZN(
        n64256) );
  AOI22_X1 U49856 ( .A1(n67593), .A2(n66543), .B1(n58420), .B2(n67587), .ZN(
        n64254) );
  AOI22_X1 U49857 ( .A1(n67617), .A2(n57031), .B1(n67611), .B2(n58696), .ZN(
        n64253) );
  AOI22_X1 U49858 ( .A1(n67569), .A2(n9001), .B1(n67563), .B2(n57017), .ZN(
        n64236) );
  AOI22_X1 U49859 ( .A1(n67593), .A2(n66544), .B1(n58421), .B2(n67587), .ZN(
        n64234) );
  AOI22_X1 U49860 ( .A1(n67617), .A2(n57007), .B1(n67611), .B2(n58697), .ZN(
        n64233) );
  AOI22_X1 U49861 ( .A1(n67569), .A2(n8999), .B1(n67563), .B2(n56993), .ZN(
        n64216) );
  AOI22_X1 U49862 ( .A1(n67593), .A2(n66545), .B1(n58422), .B2(n67587), .ZN(
        n64214) );
  AOI22_X1 U49863 ( .A1(n67617), .A2(n56983), .B1(n67611), .B2(n58698), .ZN(
        n64213) );
  AOI22_X1 U49864 ( .A1(n67569), .A2(n8997), .B1(n67563), .B2(n56969), .ZN(
        n64196) );
  AOI22_X1 U49865 ( .A1(n67593), .A2(n66546), .B1(n58423), .B2(n67587), .ZN(
        n64194) );
  AOI22_X1 U49866 ( .A1(n67617), .A2(n56959), .B1(n67611), .B2(n58699), .ZN(
        n64193) );
  AOI22_X1 U49867 ( .A1(n67569), .A2(n8995), .B1(n67563), .B2(n56945), .ZN(
        n64176) );
  AOI22_X1 U49868 ( .A1(n67593), .A2(n66547), .B1(n58424), .B2(n67587), .ZN(
        n64174) );
  AOI22_X1 U49869 ( .A1(n67617), .A2(n56935), .B1(n67611), .B2(n58700), .ZN(
        n64173) );
  AOI22_X1 U49870 ( .A1(n67569), .A2(n8993), .B1(n67563), .B2(n56921), .ZN(
        n64156) );
  AOI22_X1 U49871 ( .A1(n67593), .A2(n66548), .B1(n58425), .B2(n67587), .ZN(
        n64154) );
  AOI22_X1 U49872 ( .A1(n67617), .A2(n56911), .B1(n67611), .B2(n58701), .ZN(
        n64153) );
  AOI22_X1 U49873 ( .A1(n67569), .A2(n8991), .B1(n67563), .B2(n56897), .ZN(
        n64136) );
  AOI22_X1 U49874 ( .A1(n67593), .A2(n66549), .B1(n58426), .B2(n67587), .ZN(
        n64134) );
  AOI22_X1 U49875 ( .A1(n67617), .A2(n56887), .B1(n67611), .B2(n58702), .ZN(
        n64133) );
  AOI22_X1 U49876 ( .A1(n67570), .A2(n8989), .B1(n67564), .B2(n56873), .ZN(
        n64116) );
  AOI22_X1 U49877 ( .A1(n67618), .A2(n56863), .B1(n67612), .B2(n58703), .ZN(
        n64113) );
  AOI22_X1 U49878 ( .A1(n67570), .A2(n8987), .B1(n67564), .B2(n56849), .ZN(
        n64096) );
  AOI22_X1 U49879 ( .A1(n67618), .A2(n56839), .B1(n67612), .B2(n58704), .ZN(
        n64093) );
  AOI22_X1 U49880 ( .A1(n67570), .A2(n8985), .B1(n67564), .B2(n56825), .ZN(
        n64076) );
  AOI22_X1 U49881 ( .A1(n67618), .A2(n56815), .B1(n67612), .B2(n58705), .ZN(
        n64073) );
  AOI22_X1 U49882 ( .A1(n67570), .A2(n8983), .B1(n67564), .B2(n56801), .ZN(
        n64056) );
  AOI22_X1 U49883 ( .A1(n67618), .A2(n56791), .B1(n67612), .B2(n58706), .ZN(
        n64053) );
  AOI22_X1 U49884 ( .A1(n67570), .A2(n8981), .B1(n67564), .B2(n56777), .ZN(
        n64036) );
  AOI22_X1 U49885 ( .A1(n67618), .A2(n58643), .B1(n67612), .B2(n58707), .ZN(
        n64033) );
  AOI22_X1 U49886 ( .A1(n67570), .A2(n8979), .B1(n67564), .B2(n56753), .ZN(
        n64016) );
  AOI22_X1 U49887 ( .A1(n67618), .A2(n58644), .B1(n67612), .B2(n58708), .ZN(
        n64013) );
  AOI22_X1 U49888 ( .A1(n67570), .A2(n8977), .B1(n67564), .B2(n56729), .ZN(
        n63996) );
  AOI22_X1 U49889 ( .A1(n67618), .A2(n58645), .B1(n67612), .B2(n58709), .ZN(
        n63993) );
  AOI22_X1 U49890 ( .A1(n67570), .A2(n8975), .B1(n67564), .B2(n56705), .ZN(
        n63976) );
  AOI22_X1 U49891 ( .A1(n67618), .A2(n58646), .B1(n67612), .B2(n58710), .ZN(
        n63973) );
  AOI22_X1 U49892 ( .A1(n67570), .A2(n8973), .B1(n67564), .B2(n56681), .ZN(
        n63956) );
  AOI22_X1 U49893 ( .A1(n67618), .A2(n58647), .B1(n67612), .B2(n58711), .ZN(
        n63953) );
  AOI22_X1 U49894 ( .A1(n67570), .A2(n8971), .B1(n67564), .B2(n56657), .ZN(
        n63936) );
  AOI22_X1 U49895 ( .A1(n67618), .A2(n58648), .B1(n67612), .B2(n58712), .ZN(
        n63933) );
  AOI22_X1 U49896 ( .A1(n67570), .A2(n8969), .B1(n67564), .B2(n56633), .ZN(
        n63916) );
  AOI22_X1 U49897 ( .A1(n67618), .A2(n58649), .B1(n67612), .B2(n58713), .ZN(
        n63913) );
  AOI22_X1 U49898 ( .A1(n67570), .A2(n8967), .B1(n67564), .B2(n56609), .ZN(
        n63896) );
  AOI22_X1 U49899 ( .A1(n67618), .A2(n58650), .B1(n67612), .B2(n58714), .ZN(
        n63893) );
  OAI221_X1 U49900 ( .B1(n63427), .B2(n67452), .C1(n49232), .C2(n67446), .A(
        n66275), .ZN(n66274) );
  AOI22_X1 U49901 ( .A1(n67440), .A2(n58379), .B1(n67434), .B2(OUT2[0]), .ZN(
        n66275) );
  OAI221_X1 U49902 ( .B1(n63426), .B2(n67452), .C1(n49233), .C2(n67446), .A(
        n66257), .ZN(n66256) );
  AOI22_X1 U49903 ( .A1(n67440), .A2(n58380), .B1(n67434), .B2(OUT2[1]), .ZN(
        n66257) );
  OAI221_X1 U49904 ( .B1(n63425), .B2(n67452), .C1(n49234), .C2(n67446), .A(
        n66239), .ZN(n66238) );
  AOI22_X1 U49905 ( .A1(n67440), .A2(n58381), .B1(n67434), .B2(OUT2[2]), .ZN(
        n66239) );
  OAI221_X1 U49906 ( .B1(n63424), .B2(n67452), .C1(n49235), .C2(n67446), .A(
        n66221), .ZN(n66220) );
  AOI22_X1 U49907 ( .A1(n67440), .A2(n58382), .B1(n67434), .B2(OUT2[3]), .ZN(
        n66221) );
  OAI221_X1 U49908 ( .B1(n63423), .B2(n67452), .C1(n49236), .C2(n67446), .A(
        n66203), .ZN(n66202) );
  AOI22_X1 U49909 ( .A1(n67440), .A2(n58383), .B1(n67434), .B2(OUT2[4]), .ZN(
        n66203) );
  OAI221_X1 U49910 ( .B1(n63422), .B2(n67452), .C1(n49237), .C2(n67446), .A(
        n66185), .ZN(n66184) );
  AOI22_X1 U49911 ( .A1(n67440), .A2(n58384), .B1(n67434), .B2(OUT2[5]), .ZN(
        n66185) );
  OAI221_X1 U49912 ( .B1(n63421), .B2(n67452), .C1(n49238), .C2(n67446), .A(
        n66167), .ZN(n66166) );
  AOI22_X1 U49913 ( .A1(n67440), .A2(n58385), .B1(n67434), .B2(OUT2[6]), .ZN(
        n66167) );
  OAI221_X1 U49914 ( .B1(n63420), .B2(n67452), .C1(n49239), .C2(n67446), .A(
        n66149), .ZN(n66148) );
  AOI22_X1 U49915 ( .A1(n67440), .A2(n58386), .B1(n67434), .B2(OUT2[7]), .ZN(
        n66149) );
  OAI221_X1 U49916 ( .B1(n63419), .B2(n67452), .C1(n49240), .C2(n67446), .A(
        n66131), .ZN(n66130) );
  AOI22_X1 U49917 ( .A1(n67440), .A2(n58387), .B1(n67434), .B2(OUT2[8]), .ZN(
        n66131) );
  OAI221_X1 U49918 ( .B1(n63418), .B2(n67452), .C1(n49241), .C2(n67446), .A(
        n66113), .ZN(n66112) );
  AOI22_X1 U49919 ( .A1(n67440), .A2(n58388), .B1(n67435), .B2(OUT2[9]), .ZN(
        n66113) );
  OAI221_X1 U49920 ( .B1(n63417), .B2(n67452), .C1(n49242), .C2(n67446), .A(
        n66095), .ZN(n66094) );
  AOI22_X1 U49921 ( .A1(n67440), .A2(n58389), .B1(n67435), .B2(OUT2[10]), .ZN(
        n66095) );
  OAI221_X1 U49922 ( .B1(n63416), .B2(n67452), .C1(n49243), .C2(n67446), .A(
        n66077), .ZN(n66076) );
  AOI22_X1 U49923 ( .A1(n67440), .A2(n58390), .B1(n67435), .B2(OUT2[11]), .ZN(
        n66077) );
  OAI221_X1 U49924 ( .B1(n63100), .B2(n67631), .C1(n62229), .C2(n67625), .A(
        n63872), .ZN(n63869) );
  AOI22_X1 U49925 ( .A1(n67619), .A2(n58651), .B1(n67613), .B2(n58715), .ZN(
        n63872) );
  OAI221_X1 U49926 ( .B1(n63099), .B2(n67631), .C1(n62228), .C2(n67625), .A(
        n63851), .ZN(n63848) );
  AOI22_X1 U49927 ( .A1(n67619), .A2(n58652), .B1(n67613), .B2(n58716), .ZN(
        n63851) );
  OAI221_X1 U49928 ( .B1(n63098), .B2(n67631), .C1(n62227), .C2(n67625), .A(
        n63830), .ZN(n63827) );
  AOI22_X1 U49929 ( .A1(n67619), .A2(n58653), .B1(n67613), .B2(n58717), .ZN(
        n63830) );
  OAI221_X1 U49930 ( .B1(n62424), .B2(n67607), .C1(n63501), .C2(n67601), .A(
        n63787), .ZN(n63772) );
  AOI22_X1 U49931 ( .A1(n67595), .A2(n66550), .B1(n67589), .B2(n58378), .ZN(
        n63787) );
  OAI221_X1 U49932 ( .B1(n63096), .B2(n67631), .C1(n62225), .C2(n67625), .A(
        n63782), .ZN(n63773) );
  AOI22_X1 U49933 ( .A1(n67619), .A2(n58654), .B1(n67613), .B2(n58718), .ZN(
        n63782) );
  OAI22_X1 U49934 ( .A1(n54670), .A2(n67725), .B1(n68060), .B2(n67719), .ZN(
        n5759) );
  OAI22_X1 U49935 ( .A1(n54669), .A2(n67725), .B1(n68063), .B2(n67719), .ZN(
        n5760) );
  OAI22_X1 U49936 ( .A1(n54668), .A2(n67725), .B1(n68066), .B2(n67719), .ZN(
        n5761) );
  OAI22_X1 U49937 ( .A1(n54667), .A2(n67725), .B1(n68069), .B2(n67719), .ZN(
        n5762) );
  OAI22_X1 U49938 ( .A1(n54666), .A2(n67725), .B1(n68072), .B2(n67719), .ZN(
        n5763) );
  OAI22_X1 U49939 ( .A1(n54665), .A2(n67725), .B1(n68075), .B2(n67719), .ZN(
        n5764) );
  OAI22_X1 U49940 ( .A1(n54664), .A2(n67725), .B1(n68078), .B2(n67719), .ZN(
        n5765) );
  OAI22_X1 U49941 ( .A1(n54663), .A2(n67725), .B1(n68081), .B2(n67719), .ZN(
        n5766) );
  OAI22_X1 U49942 ( .A1(n54662), .A2(n67725), .B1(n68084), .B2(n67719), .ZN(
        n5767) );
  OAI22_X1 U49943 ( .A1(n54661), .A2(n67725), .B1(n68087), .B2(n67719), .ZN(
        n5768) );
  OAI22_X1 U49944 ( .A1(n54660), .A2(n67725), .B1(n68090), .B2(n67719), .ZN(
        n5769) );
  OAI22_X1 U49945 ( .A1(n54659), .A2(n67726), .B1(n68093), .B2(n67719), .ZN(
        n5770) );
  OAI22_X1 U49946 ( .A1(n54658), .A2(n67726), .B1(n68096), .B2(n67720), .ZN(
        n5771) );
  OAI22_X1 U49947 ( .A1(n54657), .A2(n67726), .B1(n68099), .B2(n67720), .ZN(
        n5772) );
  OAI22_X1 U49948 ( .A1(n54656), .A2(n67726), .B1(n68102), .B2(n67720), .ZN(
        n5773) );
  OAI22_X1 U49949 ( .A1(n54655), .A2(n67726), .B1(n68105), .B2(n67720), .ZN(
        n5774) );
  OAI22_X1 U49950 ( .A1(n54654), .A2(n67726), .B1(n68108), .B2(n67720), .ZN(
        n5775) );
  OAI22_X1 U49951 ( .A1(n54653), .A2(n67726), .B1(n68111), .B2(n67720), .ZN(
        n5776) );
  OAI22_X1 U49952 ( .A1(n54652), .A2(n67726), .B1(n68114), .B2(n67720), .ZN(
        n5777) );
  OAI22_X1 U49953 ( .A1(n54651), .A2(n67726), .B1(n68117), .B2(n67720), .ZN(
        n5778) );
  OAI22_X1 U49954 ( .A1(n54650), .A2(n67726), .B1(n68120), .B2(n67720), .ZN(
        n5779) );
  OAI22_X1 U49955 ( .A1(n54649), .A2(n67726), .B1(n68123), .B2(n67720), .ZN(
        n5780) );
  OAI22_X1 U49956 ( .A1(n54648), .A2(n67726), .B1(n68126), .B2(n67720), .ZN(
        n5781) );
  OAI22_X1 U49957 ( .A1(n54647), .A2(n67727), .B1(n68129), .B2(n67720), .ZN(
        n5782) );
  OAI22_X1 U49958 ( .A1(n54646), .A2(n67727), .B1(n68132), .B2(n67721), .ZN(
        n5783) );
  OAI22_X1 U49959 ( .A1(n54645), .A2(n67727), .B1(n68135), .B2(n67721), .ZN(
        n5784) );
  OAI22_X1 U49960 ( .A1(n54644), .A2(n67727), .B1(n68138), .B2(n67721), .ZN(
        n5785) );
  OAI22_X1 U49961 ( .A1(n54643), .A2(n67727), .B1(n68141), .B2(n67721), .ZN(
        n5786) );
  OAI22_X1 U49962 ( .A1(n54642), .A2(n67727), .B1(n68144), .B2(n67721), .ZN(
        n5787) );
  OAI22_X1 U49963 ( .A1(n54641), .A2(n67727), .B1(n68147), .B2(n67721), .ZN(
        n5788) );
  OAI22_X1 U49964 ( .A1(n54640), .A2(n67727), .B1(n68150), .B2(n67721), .ZN(
        n5789) );
  OAI22_X1 U49965 ( .A1(n54639), .A2(n67727), .B1(n68153), .B2(n67721), .ZN(
        n5790) );
  OAI22_X1 U49966 ( .A1(n54638), .A2(n67727), .B1(n68156), .B2(n67721), .ZN(
        n5791) );
  OAI22_X1 U49967 ( .A1(n54637), .A2(n67727), .B1(n68159), .B2(n67721), .ZN(
        n5792) );
  OAI22_X1 U49968 ( .A1(n54636), .A2(n67727), .B1(n68162), .B2(n67721), .ZN(
        n5793) );
  OAI22_X1 U49969 ( .A1(n54635), .A2(n67728), .B1(n68165), .B2(n67721), .ZN(
        n5794) );
  OAI22_X1 U49970 ( .A1(n54634), .A2(n67728), .B1(n68168), .B2(n67722), .ZN(
        n5795) );
  OAI22_X1 U49971 ( .A1(n54633), .A2(n67728), .B1(n68171), .B2(n67722), .ZN(
        n5796) );
  OAI22_X1 U49972 ( .A1(n54632), .A2(n67728), .B1(n68174), .B2(n67722), .ZN(
        n5797) );
  OAI22_X1 U49973 ( .A1(n54631), .A2(n67728), .B1(n68177), .B2(n67722), .ZN(
        n5798) );
  OAI22_X1 U49974 ( .A1(n54630), .A2(n67728), .B1(n68180), .B2(n67722), .ZN(
        n5799) );
  OAI22_X1 U49975 ( .A1(n54629), .A2(n67728), .B1(n68183), .B2(n67722), .ZN(
        n5800) );
  OAI22_X1 U49976 ( .A1(n54628), .A2(n67728), .B1(n68186), .B2(n67722), .ZN(
        n5801) );
  OAI22_X1 U49977 ( .A1(n54627), .A2(n67728), .B1(n68189), .B2(n67722), .ZN(
        n5802) );
  OAI22_X1 U49978 ( .A1(n54626), .A2(n67728), .B1(n68192), .B2(n67722), .ZN(
        n5803) );
  OAI22_X1 U49979 ( .A1(n54625), .A2(n67728), .B1(n68195), .B2(n67722), .ZN(
        n5804) );
  OAI22_X1 U49980 ( .A1(n54624), .A2(n67728), .B1(n68198), .B2(n67722), .ZN(
        n5805) );
  OAI22_X1 U49981 ( .A1(n54623), .A2(n67729), .B1(n68201), .B2(n67722), .ZN(
        n5806) );
  OAI22_X1 U49982 ( .A1(n54622), .A2(n67729), .B1(n68204), .B2(n67723), .ZN(
        n5807) );
  OAI22_X1 U49983 ( .A1(n54621), .A2(n67729), .B1(n68207), .B2(n67723), .ZN(
        n5808) );
  OAI22_X1 U49984 ( .A1(n54620), .A2(n67729), .B1(n68210), .B2(n67723), .ZN(
        n5809) );
  OAI22_X1 U49985 ( .A1(n54619), .A2(n67729), .B1(n68213), .B2(n67723), .ZN(
        n5810) );
  OAI22_X1 U49986 ( .A1(n54618), .A2(n67729), .B1(n68216), .B2(n67723), .ZN(
        n5811) );
  OAI22_X1 U49987 ( .A1(n54617), .A2(n67729), .B1(n68219), .B2(n67723), .ZN(
        n5812) );
  OAI22_X1 U49988 ( .A1(n54616), .A2(n67729), .B1(n68222), .B2(n67723), .ZN(
        n5813) );
  OAI22_X1 U49989 ( .A1(n54615), .A2(n67729), .B1(n68225), .B2(n67723), .ZN(
        n5814) );
  OAI22_X1 U49990 ( .A1(n54614), .A2(n67729), .B1(n68228), .B2(n67723), .ZN(
        n5815) );
  OAI22_X1 U49991 ( .A1(n54613), .A2(n67729), .B1(n68231), .B2(n67723), .ZN(
        n5816) );
  OAI22_X1 U49992 ( .A1(n54612), .A2(n67729), .B1(n68234), .B2(n67723), .ZN(
        n5817) );
  OAI22_X1 U49993 ( .A1(n54611), .A2(n67730), .B1(n68237), .B2(n67723), .ZN(
        n5818) );
  OAI22_X1 U49994 ( .A1(n67662), .A2(n65063), .B1(n68060), .B2(n67654), .ZN(
        n5376) );
  OAI22_X1 U49995 ( .A1(n67662), .A2(n65043), .B1(n68063), .B2(n67654), .ZN(
        n5378) );
  OAI22_X1 U49996 ( .A1(n67662), .A2(n65023), .B1(n68066), .B2(n67654), .ZN(
        n5380) );
  OAI22_X1 U49997 ( .A1(n67662), .A2(n65003), .B1(n68069), .B2(n67654), .ZN(
        n5382) );
  OAI22_X1 U49998 ( .A1(n67662), .A2(n64983), .B1(n68072), .B2(n67654), .ZN(
        n5384) );
  OAI22_X1 U49999 ( .A1(n67662), .A2(n64963), .B1(n68075), .B2(n67654), .ZN(
        n5386) );
  OAI22_X1 U50000 ( .A1(n67662), .A2(n64943), .B1(n68078), .B2(n67654), .ZN(
        n5388) );
  OAI22_X1 U50001 ( .A1(n67662), .A2(n64923), .B1(n68081), .B2(n67654), .ZN(
        n5390) );
  OAI22_X1 U50002 ( .A1(n67662), .A2(n64903), .B1(n68084), .B2(n67654), .ZN(
        n5392) );
  OAI22_X1 U50003 ( .A1(n67662), .A2(n64883), .B1(n68087), .B2(n67654), .ZN(
        n5394) );
  OAI22_X1 U50004 ( .A1(n67662), .A2(n64863), .B1(n68090), .B2(n67654), .ZN(
        n5396) );
  OAI22_X1 U50005 ( .A1(n67662), .A2(n64843), .B1(n68093), .B2(n67654), .ZN(
        n5398) );
  OAI22_X1 U50006 ( .A1(n67663), .A2(n64823), .B1(n68096), .B2(n67655), .ZN(
        n5400) );
  OAI22_X1 U50007 ( .A1(n67663), .A2(n64803), .B1(n68099), .B2(n67655), .ZN(
        n5402) );
  OAI22_X1 U50008 ( .A1(n67663), .A2(n64783), .B1(n68102), .B2(n67655), .ZN(
        n5404) );
  OAI22_X1 U50009 ( .A1(n67663), .A2(n64763), .B1(n68105), .B2(n67655), .ZN(
        n5406) );
  OAI22_X1 U50010 ( .A1(n67663), .A2(n64743), .B1(n68108), .B2(n67655), .ZN(
        n5408) );
  OAI22_X1 U50011 ( .A1(n67663), .A2(n64723), .B1(n68111), .B2(n67655), .ZN(
        n5410) );
  OAI22_X1 U50012 ( .A1(n67663), .A2(n64703), .B1(n68114), .B2(n67655), .ZN(
        n5412) );
  OAI22_X1 U50013 ( .A1(n67663), .A2(n64683), .B1(n68117), .B2(n67655), .ZN(
        n5414) );
  OAI22_X1 U50014 ( .A1(n67663), .A2(n64663), .B1(n68120), .B2(n67655), .ZN(
        n5416) );
  OAI22_X1 U50015 ( .A1(n67663), .A2(n64643), .B1(n68123), .B2(n67655), .ZN(
        n5418) );
  OAI22_X1 U50016 ( .A1(n67663), .A2(n64623), .B1(n68126), .B2(n67655), .ZN(
        n5420) );
  OAI22_X1 U50017 ( .A1(n67663), .A2(n64603), .B1(n68129), .B2(n67655), .ZN(
        n5422) );
  OAI22_X1 U50018 ( .A1(n67663), .A2(n64583), .B1(n68132), .B2(n67656), .ZN(
        n5424) );
  OAI22_X1 U50019 ( .A1(n67664), .A2(n64563), .B1(n68135), .B2(n67656), .ZN(
        n5426) );
  OAI22_X1 U50020 ( .A1(n67664), .A2(n64543), .B1(n68138), .B2(n67656), .ZN(
        n5428) );
  OAI22_X1 U50021 ( .A1(n67664), .A2(n64523), .B1(n68141), .B2(n67656), .ZN(
        n5430) );
  OAI22_X1 U50022 ( .A1(n67664), .A2(n64503), .B1(n68144), .B2(n67656), .ZN(
        n5432) );
  OAI22_X1 U50023 ( .A1(n67664), .A2(n64483), .B1(n68147), .B2(n67656), .ZN(
        n5434) );
  OAI22_X1 U50024 ( .A1(n67664), .A2(n64463), .B1(n68150), .B2(n67656), .ZN(
        n5436) );
  OAI22_X1 U50025 ( .A1(n67664), .A2(n64443), .B1(n68153), .B2(n67656), .ZN(
        n5438) );
  OAI22_X1 U50026 ( .A1(n67664), .A2(n64423), .B1(n68156), .B2(n67656), .ZN(
        n5440) );
  OAI22_X1 U50027 ( .A1(n67664), .A2(n64403), .B1(n68159), .B2(n67656), .ZN(
        n5442) );
  OAI22_X1 U50028 ( .A1(n67664), .A2(n64383), .B1(n68162), .B2(n67656), .ZN(
        n5444) );
  OAI22_X1 U50029 ( .A1(n67664), .A2(n64363), .B1(n68165), .B2(n67656), .ZN(
        n5446) );
  OAI22_X1 U50030 ( .A1(n67664), .A2(n64343), .B1(n68168), .B2(n67657), .ZN(
        n5448) );
  OAI22_X1 U50031 ( .A1(n67664), .A2(n64323), .B1(n68171), .B2(n67657), .ZN(
        n5450) );
  OAI22_X1 U50032 ( .A1(n67665), .A2(n64303), .B1(n68174), .B2(n67657), .ZN(
        n5452) );
  OAI22_X1 U50033 ( .A1(n67665), .A2(n64283), .B1(n68177), .B2(n67657), .ZN(
        n5454) );
  OAI22_X1 U50034 ( .A1(n67665), .A2(n64263), .B1(n68180), .B2(n67657), .ZN(
        n5456) );
  OAI22_X1 U50035 ( .A1(n67665), .A2(n64243), .B1(n68183), .B2(n67657), .ZN(
        n5458) );
  OAI22_X1 U50036 ( .A1(n67665), .A2(n64223), .B1(n68186), .B2(n67657), .ZN(
        n5460) );
  OAI22_X1 U50037 ( .A1(n67665), .A2(n64203), .B1(n68189), .B2(n67657), .ZN(
        n5462) );
  OAI22_X1 U50038 ( .A1(n67665), .A2(n64183), .B1(n68192), .B2(n67657), .ZN(
        n5464) );
  OAI22_X1 U50039 ( .A1(n67665), .A2(n64163), .B1(n68195), .B2(n67657), .ZN(
        n5466) );
  OAI22_X1 U50040 ( .A1(n67665), .A2(n64143), .B1(n68198), .B2(n67657), .ZN(
        n5468) );
  OAI22_X1 U50041 ( .A1(n67665), .A2(n64123), .B1(n68201), .B2(n67657), .ZN(
        n5470) );
  OAI22_X1 U50042 ( .A1(n67665), .A2(n64103), .B1(n68204), .B2(n67658), .ZN(
        n5472) );
  OAI22_X1 U50043 ( .A1(n67665), .A2(n64083), .B1(n68207), .B2(n67658), .ZN(
        n5474) );
  OAI22_X1 U50044 ( .A1(n67665), .A2(n64063), .B1(n68210), .B2(n67658), .ZN(
        n5476) );
  OAI22_X1 U50045 ( .A1(n67666), .A2(n64043), .B1(n68213), .B2(n67658), .ZN(
        n5478) );
  OAI22_X1 U50046 ( .A1(n67666), .A2(n64023), .B1(n68216), .B2(n67658), .ZN(
        n5480) );
  OAI22_X1 U50047 ( .A1(n67666), .A2(n64003), .B1(n68219), .B2(n67658), .ZN(
        n5482) );
  OAI22_X1 U50048 ( .A1(n67666), .A2(n63983), .B1(n68222), .B2(n67658), .ZN(
        n5484) );
  OAI22_X1 U50049 ( .A1(n67666), .A2(n63963), .B1(n68225), .B2(n67658), .ZN(
        n5486) );
  OAI22_X1 U50050 ( .A1(n67666), .A2(n63943), .B1(n68228), .B2(n67658), .ZN(
        n5488) );
  OAI22_X1 U50051 ( .A1(n67666), .A2(n63923), .B1(n68231), .B2(n67658), .ZN(
        n5490) );
  OAI22_X1 U50052 ( .A1(n67666), .A2(n63903), .B1(n68234), .B2(n67658), .ZN(
        n5492) );
  OAI22_X1 U50053 ( .A1(n67666), .A2(n63883), .B1(n68237), .B2(n67658), .ZN(
        n5494) );
  OAI22_X1 U50054 ( .A1(n67675), .A2(n63763), .B1(n68060), .B2(n67667), .ZN(
        n5503) );
  OAI22_X1 U50055 ( .A1(n67675), .A2(n63762), .B1(n68063), .B2(n67667), .ZN(
        n5504) );
  OAI22_X1 U50056 ( .A1(n67675), .A2(n63761), .B1(n68066), .B2(n67667), .ZN(
        n5505) );
  OAI22_X1 U50057 ( .A1(n67675), .A2(n63760), .B1(n68069), .B2(n67667), .ZN(
        n5506) );
  OAI22_X1 U50058 ( .A1(n67675), .A2(n63759), .B1(n68072), .B2(n67667), .ZN(
        n5507) );
  OAI22_X1 U50059 ( .A1(n67675), .A2(n63758), .B1(n68075), .B2(n67667), .ZN(
        n5508) );
  OAI22_X1 U50060 ( .A1(n67675), .A2(n63757), .B1(n68078), .B2(n67667), .ZN(
        n5509) );
  OAI22_X1 U50061 ( .A1(n67675), .A2(n63756), .B1(n68081), .B2(n67667), .ZN(
        n5510) );
  OAI22_X1 U50062 ( .A1(n67675), .A2(n63755), .B1(n68084), .B2(n67667), .ZN(
        n5511) );
  OAI22_X1 U50063 ( .A1(n67675), .A2(n63754), .B1(n68087), .B2(n67667), .ZN(
        n5512) );
  OAI22_X1 U50064 ( .A1(n67675), .A2(n63753), .B1(n68090), .B2(n67667), .ZN(
        n5513) );
  OAI22_X1 U50065 ( .A1(n67675), .A2(n63752), .B1(n68093), .B2(n67667), .ZN(
        n5514) );
  OAI22_X1 U50066 ( .A1(n67676), .A2(n63751), .B1(n68096), .B2(n67668), .ZN(
        n5515) );
  OAI22_X1 U50067 ( .A1(n67676), .A2(n63750), .B1(n68099), .B2(n67668), .ZN(
        n5516) );
  OAI22_X1 U50068 ( .A1(n67676), .A2(n63749), .B1(n68102), .B2(n67668), .ZN(
        n5517) );
  OAI22_X1 U50069 ( .A1(n67676), .A2(n63748), .B1(n68105), .B2(n67668), .ZN(
        n5518) );
  OAI22_X1 U50070 ( .A1(n67676), .A2(n63747), .B1(n68108), .B2(n67668), .ZN(
        n5519) );
  OAI22_X1 U50071 ( .A1(n67676), .A2(n63746), .B1(n68111), .B2(n67668), .ZN(
        n5520) );
  OAI22_X1 U50072 ( .A1(n67676), .A2(n63745), .B1(n68114), .B2(n67668), .ZN(
        n5521) );
  OAI22_X1 U50073 ( .A1(n67676), .A2(n63744), .B1(n68117), .B2(n67668), .ZN(
        n5522) );
  OAI22_X1 U50074 ( .A1(n67676), .A2(n63743), .B1(n68120), .B2(n67668), .ZN(
        n5523) );
  OAI22_X1 U50075 ( .A1(n67676), .A2(n63742), .B1(n68123), .B2(n67668), .ZN(
        n5524) );
  OAI22_X1 U50076 ( .A1(n67676), .A2(n63741), .B1(n68126), .B2(n67668), .ZN(
        n5525) );
  OAI22_X1 U50077 ( .A1(n67676), .A2(n63740), .B1(n68129), .B2(n67668), .ZN(
        n5526) );
  OAI22_X1 U50078 ( .A1(n67676), .A2(n63739), .B1(n68132), .B2(n67669), .ZN(
        n5527) );
  OAI22_X1 U50079 ( .A1(n67677), .A2(n63738), .B1(n68135), .B2(n67669), .ZN(
        n5528) );
  OAI22_X1 U50080 ( .A1(n67677), .A2(n63737), .B1(n68138), .B2(n67669), .ZN(
        n5529) );
  OAI22_X1 U50081 ( .A1(n67677), .A2(n63736), .B1(n68141), .B2(n67669), .ZN(
        n5530) );
  OAI22_X1 U50082 ( .A1(n67677), .A2(n63735), .B1(n68144), .B2(n67669), .ZN(
        n5531) );
  OAI22_X1 U50083 ( .A1(n67677), .A2(n63734), .B1(n68147), .B2(n67669), .ZN(
        n5532) );
  OAI22_X1 U50084 ( .A1(n67677), .A2(n63733), .B1(n68150), .B2(n67669), .ZN(
        n5533) );
  OAI22_X1 U50085 ( .A1(n67677), .A2(n63732), .B1(n68153), .B2(n67669), .ZN(
        n5534) );
  OAI22_X1 U50086 ( .A1(n67677), .A2(n63731), .B1(n68156), .B2(n67669), .ZN(
        n5535) );
  OAI22_X1 U50087 ( .A1(n67677), .A2(n63730), .B1(n68159), .B2(n67669), .ZN(
        n5536) );
  OAI22_X1 U50088 ( .A1(n67677), .A2(n63729), .B1(n68162), .B2(n67669), .ZN(
        n5537) );
  OAI22_X1 U50089 ( .A1(n67677), .A2(n63728), .B1(n68165), .B2(n67669), .ZN(
        n5538) );
  OAI22_X1 U50090 ( .A1(n67677), .A2(n63727), .B1(n68168), .B2(n67670), .ZN(
        n5539) );
  OAI22_X1 U50091 ( .A1(n67677), .A2(n63726), .B1(n68171), .B2(n67670), .ZN(
        n5540) );
  OAI22_X1 U50092 ( .A1(n67678), .A2(n63725), .B1(n68174), .B2(n67670), .ZN(
        n5541) );
  OAI22_X1 U50093 ( .A1(n67678), .A2(n63724), .B1(n68177), .B2(n67670), .ZN(
        n5542) );
  OAI22_X1 U50094 ( .A1(n67678), .A2(n63723), .B1(n68180), .B2(n67670), .ZN(
        n5543) );
  OAI22_X1 U50095 ( .A1(n67678), .A2(n63722), .B1(n68183), .B2(n67670), .ZN(
        n5544) );
  OAI22_X1 U50096 ( .A1(n67678), .A2(n63721), .B1(n68186), .B2(n67670), .ZN(
        n5545) );
  OAI22_X1 U50097 ( .A1(n67678), .A2(n63720), .B1(n68189), .B2(n67670), .ZN(
        n5546) );
  OAI22_X1 U50098 ( .A1(n67678), .A2(n63719), .B1(n68192), .B2(n67670), .ZN(
        n5547) );
  OAI22_X1 U50099 ( .A1(n67678), .A2(n63718), .B1(n68195), .B2(n67670), .ZN(
        n5548) );
  OAI22_X1 U50100 ( .A1(n67678), .A2(n63717), .B1(n68198), .B2(n67670), .ZN(
        n5549) );
  OAI22_X1 U50101 ( .A1(n67678), .A2(n63716), .B1(n68201), .B2(n67670), .ZN(
        n5550) );
  OAI22_X1 U50102 ( .A1(n67678), .A2(n63715), .B1(n68204), .B2(n67671), .ZN(
        n5551) );
  OAI22_X1 U50103 ( .A1(n67678), .A2(n63714), .B1(n68207), .B2(n67671), .ZN(
        n5552) );
  OAI22_X1 U50104 ( .A1(n67678), .A2(n63713), .B1(n68210), .B2(n67671), .ZN(
        n5553) );
  OAI22_X1 U50105 ( .A1(n67679), .A2(n63712), .B1(n68213), .B2(n67671), .ZN(
        n5554) );
  OAI22_X1 U50106 ( .A1(n67679), .A2(n63711), .B1(n68216), .B2(n67671), .ZN(
        n5555) );
  OAI22_X1 U50107 ( .A1(n67679), .A2(n63710), .B1(n68219), .B2(n67671), .ZN(
        n5556) );
  OAI22_X1 U50108 ( .A1(n67679), .A2(n63709), .B1(n68222), .B2(n67671), .ZN(
        n5557) );
  OAI22_X1 U50109 ( .A1(n67679), .A2(n63708), .B1(n68225), .B2(n67671), .ZN(
        n5558) );
  OAI22_X1 U50110 ( .A1(n67679), .A2(n63707), .B1(n68228), .B2(n67671), .ZN(
        n5559) );
  OAI22_X1 U50111 ( .A1(n67679), .A2(n63706), .B1(n68231), .B2(n67671), .ZN(
        n5560) );
  OAI22_X1 U50112 ( .A1(n67679), .A2(n63705), .B1(n68234), .B2(n67671), .ZN(
        n5561) );
  OAI22_X1 U50113 ( .A1(n67679), .A2(n63704), .B1(n68237), .B2(n67671), .ZN(
        n5562) );
  OAI22_X1 U50114 ( .A1(n54246), .A2(n67929), .B1(n68058), .B2(n67923), .ZN(
        n6783) );
  OAI22_X1 U50115 ( .A1(n54245), .A2(n67929), .B1(n68061), .B2(n67923), .ZN(
        n6784) );
  OAI22_X1 U50116 ( .A1(n54244), .A2(n67929), .B1(n68064), .B2(n67923), .ZN(
        n6785) );
  OAI22_X1 U50117 ( .A1(n54243), .A2(n67929), .B1(n68067), .B2(n67923), .ZN(
        n6786) );
  OAI22_X1 U50118 ( .A1(n54242), .A2(n67929), .B1(n68070), .B2(n67923), .ZN(
        n6787) );
  OAI22_X1 U50119 ( .A1(n54241), .A2(n67929), .B1(n68073), .B2(n67923), .ZN(
        n6788) );
  OAI22_X1 U50120 ( .A1(n54240), .A2(n67929), .B1(n68076), .B2(n67923), .ZN(
        n6789) );
  OAI22_X1 U50121 ( .A1(n54239), .A2(n67929), .B1(n68079), .B2(n67923), .ZN(
        n6790) );
  OAI22_X1 U50122 ( .A1(n54238), .A2(n67929), .B1(n68082), .B2(n67923), .ZN(
        n6791) );
  OAI22_X1 U50123 ( .A1(n54237), .A2(n67929), .B1(n68085), .B2(n67923), .ZN(
        n6792) );
  OAI22_X1 U50124 ( .A1(n54236), .A2(n67929), .B1(n68088), .B2(n67923), .ZN(
        n6793) );
  OAI22_X1 U50125 ( .A1(n54235), .A2(n67930), .B1(n68091), .B2(n67923), .ZN(
        n6794) );
  OAI22_X1 U50126 ( .A1(n54234), .A2(n67930), .B1(n68094), .B2(n67924), .ZN(
        n6795) );
  OAI22_X1 U50127 ( .A1(n54233), .A2(n67930), .B1(n68097), .B2(n67924), .ZN(
        n6796) );
  OAI22_X1 U50128 ( .A1(n54232), .A2(n67930), .B1(n68100), .B2(n67924), .ZN(
        n6797) );
  OAI22_X1 U50129 ( .A1(n54231), .A2(n67930), .B1(n68103), .B2(n67924), .ZN(
        n6798) );
  OAI22_X1 U50130 ( .A1(n54230), .A2(n67930), .B1(n68106), .B2(n67924), .ZN(
        n6799) );
  OAI22_X1 U50131 ( .A1(n54229), .A2(n67930), .B1(n68109), .B2(n67924), .ZN(
        n6800) );
  OAI22_X1 U50132 ( .A1(n54228), .A2(n67930), .B1(n68112), .B2(n67924), .ZN(
        n6801) );
  OAI22_X1 U50133 ( .A1(n54227), .A2(n67930), .B1(n68115), .B2(n67924), .ZN(
        n6802) );
  OAI22_X1 U50134 ( .A1(n54226), .A2(n67930), .B1(n68118), .B2(n67924), .ZN(
        n6803) );
  OAI22_X1 U50135 ( .A1(n54225), .A2(n67930), .B1(n68121), .B2(n67924), .ZN(
        n6804) );
  OAI22_X1 U50136 ( .A1(n54224), .A2(n67930), .B1(n68124), .B2(n67924), .ZN(
        n6805) );
  OAI22_X1 U50137 ( .A1(n54223), .A2(n67931), .B1(n68127), .B2(n67924), .ZN(
        n6806) );
  OAI22_X1 U50138 ( .A1(n54222), .A2(n67931), .B1(n68130), .B2(n67925), .ZN(
        n6807) );
  OAI22_X1 U50139 ( .A1(n54221), .A2(n67931), .B1(n68133), .B2(n67925), .ZN(
        n6808) );
  OAI22_X1 U50140 ( .A1(n54220), .A2(n67931), .B1(n68136), .B2(n67925), .ZN(
        n6809) );
  OAI22_X1 U50141 ( .A1(n54219), .A2(n67931), .B1(n68139), .B2(n67925), .ZN(
        n6810) );
  OAI22_X1 U50142 ( .A1(n54218), .A2(n67931), .B1(n68142), .B2(n67925), .ZN(
        n6811) );
  OAI22_X1 U50143 ( .A1(n54217), .A2(n67931), .B1(n68145), .B2(n67925), .ZN(
        n6812) );
  OAI22_X1 U50144 ( .A1(n54216), .A2(n67931), .B1(n68148), .B2(n67925), .ZN(
        n6813) );
  OAI22_X1 U50145 ( .A1(n54215), .A2(n67931), .B1(n68151), .B2(n67925), .ZN(
        n6814) );
  OAI22_X1 U50146 ( .A1(n54214), .A2(n67931), .B1(n68154), .B2(n67925), .ZN(
        n6815) );
  OAI22_X1 U50147 ( .A1(n54213), .A2(n67931), .B1(n68157), .B2(n67925), .ZN(
        n6816) );
  OAI22_X1 U50148 ( .A1(n54212), .A2(n67931), .B1(n68160), .B2(n67925), .ZN(
        n6817) );
  OAI22_X1 U50149 ( .A1(n54211), .A2(n67932), .B1(n68163), .B2(n67925), .ZN(
        n6818) );
  OAI22_X1 U50150 ( .A1(n54210), .A2(n67932), .B1(n68166), .B2(n67926), .ZN(
        n6819) );
  OAI22_X1 U50151 ( .A1(n54209), .A2(n67932), .B1(n68169), .B2(n67926), .ZN(
        n6820) );
  OAI22_X1 U50152 ( .A1(n54208), .A2(n67932), .B1(n68172), .B2(n67926), .ZN(
        n6821) );
  OAI22_X1 U50153 ( .A1(n54207), .A2(n67932), .B1(n68175), .B2(n67926), .ZN(
        n6822) );
  OAI22_X1 U50154 ( .A1(n54206), .A2(n67932), .B1(n68178), .B2(n67926), .ZN(
        n6823) );
  OAI22_X1 U50155 ( .A1(n54205), .A2(n67932), .B1(n68181), .B2(n67926), .ZN(
        n6824) );
  OAI22_X1 U50156 ( .A1(n54204), .A2(n67932), .B1(n68184), .B2(n67926), .ZN(
        n6825) );
  OAI22_X1 U50157 ( .A1(n54203), .A2(n67932), .B1(n68187), .B2(n67926), .ZN(
        n6826) );
  OAI22_X1 U50158 ( .A1(n54202), .A2(n67932), .B1(n68190), .B2(n67926), .ZN(
        n6827) );
  OAI22_X1 U50159 ( .A1(n54201), .A2(n67932), .B1(n68193), .B2(n67926), .ZN(
        n6828) );
  OAI22_X1 U50160 ( .A1(n54200), .A2(n67932), .B1(n68196), .B2(n67926), .ZN(
        n6829) );
  OAI22_X1 U50161 ( .A1(n54199), .A2(n67933), .B1(n68199), .B2(n67926), .ZN(
        n6830) );
  OAI22_X1 U50162 ( .A1(n54198), .A2(n67933), .B1(n68202), .B2(n67927), .ZN(
        n6831) );
  OAI22_X1 U50163 ( .A1(n54197), .A2(n67933), .B1(n68205), .B2(n67927), .ZN(
        n6832) );
  OAI22_X1 U50164 ( .A1(n54196), .A2(n67933), .B1(n68208), .B2(n67927), .ZN(
        n6833) );
  OAI22_X1 U50165 ( .A1(n54195), .A2(n67933), .B1(n68211), .B2(n67927), .ZN(
        n6834) );
  OAI22_X1 U50166 ( .A1(n54194), .A2(n67933), .B1(n68214), .B2(n67927), .ZN(
        n6835) );
  OAI22_X1 U50167 ( .A1(n54193), .A2(n67933), .B1(n68217), .B2(n67927), .ZN(
        n6836) );
  OAI22_X1 U50168 ( .A1(n54192), .A2(n67933), .B1(n68220), .B2(n67927), .ZN(
        n6837) );
  OAI22_X1 U50169 ( .A1(n54191), .A2(n67933), .B1(n68223), .B2(n67927), .ZN(
        n6838) );
  OAI22_X1 U50170 ( .A1(n54190), .A2(n67933), .B1(n68226), .B2(n67927), .ZN(
        n6839) );
  OAI22_X1 U50171 ( .A1(n54189), .A2(n67933), .B1(n68229), .B2(n67927), .ZN(
        n6840) );
  OAI22_X1 U50172 ( .A1(n54188), .A2(n67933), .B1(n68232), .B2(n67927), .ZN(
        n6841) );
  OAI22_X1 U50173 ( .A1(n54187), .A2(n67934), .B1(n68235), .B2(n67927), .ZN(
        n6842) );
  OAI22_X1 U50174 ( .A1(n49232), .A2(n67904), .B1(n68059), .B2(n67898), .ZN(
        n6655) );
  OAI22_X1 U50175 ( .A1(n49233), .A2(n67904), .B1(n68062), .B2(n67898), .ZN(
        n6656) );
  OAI22_X1 U50176 ( .A1(n49234), .A2(n67904), .B1(n68065), .B2(n67898), .ZN(
        n6657) );
  OAI22_X1 U50177 ( .A1(n49235), .A2(n67904), .B1(n68068), .B2(n67898), .ZN(
        n6658) );
  OAI22_X1 U50178 ( .A1(n49236), .A2(n67904), .B1(n68071), .B2(n67898), .ZN(
        n6659) );
  OAI22_X1 U50179 ( .A1(n49237), .A2(n67904), .B1(n68074), .B2(n67898), .ZN(
        n6660) );
  OAI22_X1 U50180 ( .A1(n49238), .A2(n67904), .B1(n68077), .B2(n67898), .ZN(
        n6661) );
  OAI22_X1 U50181 ( .A1(n49239), .A2(n67904), .B1(n68080), .B2(n67898), .ZN(
        n6662) );
  OAI22_X1 U50182 ( .A1(n49240), .A2(n67904), .B1(n68083), .B2(n67898), .ZN(
        n6663) );
  OAI22_X1 U50183 ( .A1(n49241), .A2(n67904), .B1(n68086), .B2(n67898), .ZN(
        n6664) );
  OAI22_X1 U50184 ( .A1(n49242), .A2(n67904), .B1(n68089), .B2(n67898), .ZN(
        n6665) );
  OAI22_X1 U50185 ( .A1(n49243), .A2(n67905), .B1(n68092), .B2(n67898), .ZN(
        n6666) );
  OAI22_X1 U50186 ( .A1(n49244), .A2(n67905), .B1(n68095), .B2(n67899), .ZN(
        n6667) );
  OAI22_X1 U50187 ( .A1(n49245), .A2(n67905), .B1(n68098), .B2(n67899), .ZN(
        n6668) );
  OAI22_X1 U50188 ( .A1(n49246), .A2(n67905), .B1(n68101), .B2(n67899), .ZN(
        n6669) );
  OAI22_X1 U50189 ( .A1(n49247), .A2(n67905), .B1(n68104), .B2(n67899), .ZN(
        n6670) );
  OAI22_X1 U50190 ( .A1(n49248), .A2(n67905), .B1(n68107), .B2(n67899), .ZN(
        n6671) );
  OAI22_X1 U50191 ( .A1(n49249), .A2(n67905), .B1(n68110), .B2(n67899), .ZN(
        n6672) );
  OAI22_X1 U50192 ( .A1(n49250), .A2(n67905), .B1(n68113), .B2(n67899), .ZN(
        n6673) );
  OAI22_X1 U50193 ( .A1(n49251), .A2(n67905), .B1(n68116), .B2(n67899), .ZN(
        n6674) );
  OAI22_X1 U50194 ( .A1(n49252), .A2(n67905), .B1(n68119), .B2(n67899), .ZN(
        n6675) );
  OAI22_X1 U50195 ( .A1(n49253), .A2(n67905), .B1(n68122), .B2(n67899), .ZN(
        n6676) );
  OAI22_X1 U50196 ( .A1(n49254), .A2(n67905), .B1(n68125), .B2(n67899), .ZN(
        n6677) );
  OAI22_X1 U50197 ( .A1(n49255), .A2(n67906), .B1(n68128), .B2(n67899), .ZN(
        n6678) );
  OAI22_X1 U50198 ( .A1(n49256), .A2(n67906), .B1(n68131), .B2(n67900), .ZN(
        n6679) );
  OAI22_X1 U50199 ( .A1(n49257), .A2(n67906), .B1(n68134), .B2(n67900), .ZN(
        n6680) );
  OAI22_X1 U50200 ( .A1(n49258), .A2(n67906), .B1(n68137), .B2(n67900), .ZN(
        n6681) );
  OAI22_X1 U50201 ( .A1(n49259), .A2(n67906), .B1(n68140), .B2(n67900), .ZN(
        n6682) );
  OAI22_X1 U50202 ( .A1(n49260), .A2(n67906), .B1(n68143), .B2(n67900), .ZN(
        n6683) );
  OAI22_X1 U50203 ( .A1(n49261), .A2(n67906), .B1(n68146), .B2(n67900), .ZN(
        n6684) );
  OAI22_X1 U50204 ( .A1(n49262), .A2(n67906), .B1(n68149), .B2(n67900), .ZN(
        n6685) );
  OAI22_X1 U50205 ( .A1(n49263), .A2(n67906), .B1(n68152), .B2(n67900), .ZN(
        n6686) );
  OAI22_X1 U50206 ( .A1(n49264), .A2(n67906), .B1(n68155), .B2(n67900), .ZN(
        n6687) );
  OAI22_X1 U50207 ( .A1(n49265), .A2(n67906), .B1(n68158), .B2(n67900), .ZN(
        n6688) );
  OAI22_X1 U50208 ( .A1(n49266), .A2(n67906), .B1(n68161), .B2(n67900), .ZN(
        n6689) );
  OAI22_X1 U50209 ( .A1(n49267), .A2(n67907), .B1(n68164), .B2(n67900), .ZN(
        n6690) );
  OAI22_X1 U50210 ( .A1(n49268), .A2(n67907), .B1(n68167), .B2(n67901), .ZN(
        n6691) );
  OAI22_X1 U50211 ( .A1(n49269), .A2(n67907), .B1(n68170), .B2(n67901), .ZN(
        n6692) );
  OAI22_X1 U50212 ( .A1(n49270), .A2(n67907), .B1(n68173), .B2(n67901), .ZN(
        n6693) );
  OAI22_X1 U50213 ( .A1(n49271), .A2(n67907), .B1(n68176), .B2(n67901), .ZN(
        n6694) );
  OAI22_X1 U50214 ( .A1(n49272), .A2(n67907), .B1(n68179), .B2(n67901), .ZN(
        n6695) );
  OAI22_X1 U50215 ( .A1(n49273), .A2(n67907), .B1(n68182), .B2(n67901), .ZN(
        n6696) );
  OAI22_X1 U50216 ( .A1(n49274), .A2(n67907), .B1(n68185), .B2(n67901), .ZN(
        n6697) );
  OAI22_X1 U50217 ( .A1(n49275), .A2(n67907), .B1(n68188), .B2(n67901), .ZN(
        n6698) );
  OAI22_X1 U50218 ( .A1(n49276), .A2(n67907), .B1(n68191), .B2(n67901), .ZN(
        n6699) );
  OAI22_X1 U50219 ( .A1(n49277), .A2(n67907), .B1(n68194), .B2(n67901), .ZN(
        n6700) );
  OAI22_X1 U50220 ( .A1(n49278), .A2(n67907), .B1(n68197), .B2(n67901), .ZN(
        n6701) );
  OAI22_X1 U50221 ( .A1(n49279), .A2(n67908), .B1(n68200), .B2(n67901), .ZN(
        n6702) );
  OAI22_X1 U50222 ( .A1(n49280), .A2(n67908), .B1(n68203), .B2(n67902), .ZN(
        n6703) );
  OAI22_X1 U50223 ( .A1(n49281), .A2(n67908), .B1(n68206), .B2(n67902), .ZN(
        n6704) );
  OAI22_X1 U50224 ( .A1(n49282), .A2(n67908), .B1(n68209), .B2(n67902), .ZN(
        n6705) );
  OAI22_X1 U50225 ( .A1(n49283), .A2(n67908), .B1(n68212), .B2(n67902), .ZN(
        n6706) );
  OAI22_X1 U50226 ( .A1(n49284), .A2(n67908), .B1(n68215), .B2(n67902), .ZN(
        n6707) );
  OAI22_X1 U50227 ( .A1(n49285), .A2(n67908), .B1(n68218), .B2(n67902), .ZN(
        n6708) );
  OAI22_X1 U50228 ( .A1(n49286), .A2(n67908), .B1(n68221), .B2(n67902), .ZN(
        n6709) );
  OAI22_X1 U50229 ( .A1(n49287), .A2(n67908), .B1(n68224), .B2(n67902), .ZN(
        n6710) );
  OAI22_X1 U50230 ( .A1(n49288), .A2(n67908), .B1(n68227), .B2(n67902), .ZN(
        n6711) );
  OAI22_X1 U50231 ( .A1(n49289), .A2(n67908), .B1(n68230), .B2(n67902), .ZN(
        n6712) );
  OAI22_X1 U50232 ( .A1(n49290), .A2(n67908), .B1(n68233), .B2(n67902), .ZN(
        n6713) );
  OAI22_X1 U50233 ( .A1(n49291), .A2(n67909), .B1(n68236), .B2(n67902), .ZN(
        n6714) );
  OAI22_X1 U50234 ( .A1(n68258), .A2(n62085), .B1(n68250), .B2(n68058), .ZN(
        n7423) );
  OAI22_X1 U50235 ( .A1(n68258), .A2(n62083), .B1(n68250), .B2(n68061), .ZN(
        n7424) );
  OAI22_X1 U50236 ( .A1(n68258), .A2(n62081), .B1(n68250), .B2(n68064), .ZN(
        n7425) );
  OAI22_X1 U50237 ( .A1(n68258), .A2(n62079), .B1(n68250), .B2(n68067), .ZN(
        n7426) );
  OAI22_X1 U50238 ( .A1(n68258), .A2(n62077), .B1(n68250), .B2(n68070), .ZN(
        n7427) );
  OAI22_X1 U50239 ( .A1(n68258), .A2(n62075), .B1(n68250), .B2(n68073), .ZN(
        n7428) );
  OAI22_X1 U50240 ( .A1(n68258), .A2(n62073), .B1(n68250), .B2(n68076), .ZN(
        n7429) );
  OAI22_X1 U50241 ( .A1(n68258), .A2(n62071), .B1(n68250), .B2(n68079), .ZN(
        n7430) );
  OAI22_X1 U50242 ( .A1(n68258), .A2(n62069), .B1(n68250), .B2(n68082), .ZN(
        n7431) );
  OAI22_X1 U50243 ( .A1(n68258), .A2(n62067), .B1(n68250), .B2(n68085), .ZN(
        n7432) );
  OAI22_X1 U50244 ( .A1(n68258), .A2(n62065), .B1(n68250), .B2(n68088), .ZN(
        n7433) );
  OAI22_X1 U50245 ( .A1(n68258), .A2(n62063), .B1(n68250), .B2(n68091), .ZN(
        n7434) );
  OAI22_X1 U50246 ( .A1(n49420), .A2(n67827), .B1(n68059), .B2(n67821), .ZN(
        n6271) );
  OAI22_X1 U50247 ( .A1(n49421), .A2(n67827), .B1(n68062), .B2(n67821), .ZN(
        n6272) );
  OAI22_X1 U50248 ( .A1(n49422), .A2(n67827), .B1(n68065), .B2(n67821), .ZN(
        n6273) );
  OAI22_X1 U50249 ( .A1(n49423), .A2(n67827), .B1(n68068), .B2(n67821), .ZN(
        n6274) );
  OAI22_X1 U50250 ( .A1(n49424), .A2(n67827), .B1(n68071), .B2(n67821), .ZN(
        n6275) );
  OAI22_X1 U50251 ( .A1(n49425), .A2(n67827), .B1(n68074), .B2(n67821), .ZN(
        n6276) );
  OAI22_X1 U50252 ( .A1(n49426), .A2(n67827), .B1(n68077), .B2(n67821), .ZN(
        n6277) );
  OAI22_X1 U50253 ( .A1(n49427), .A2(n67827), .B1(n68080), .B2(n67821), .ZN(
        n6278) );
  OAI22_X1 U50254 ( .A1(n49428), .A2(n67827), .B1(n68083), .B2(n67821), .ZN(
        n6279) );
  OAI22_X1 U50255 ( .A1(n49429), .A2(n67827), .B1(n68086), .B2(n67821), .ZN(
        n6280) );
  OAI22_X1 U50256 ( .A1(n49430), .A2(n67827), .B1(n68089), .B2(n67821), .ZN(
        n6281) );
  OAI22_X1 U50257 ( .A1(n49431), .A2(n67828), .B1(n68092), .B2(n67821), .ZN(
        n6282) );
  OAI22_X1 U50258 ( .A1(n49432), .A2(n67828), .B1(n68095), .B2(n67822), .ZN(
        n6283) );
  OAI22_X1 U50259 ( .A1(n49433), .A2(n67828), .B1(n68098), .B2(n67822), .ZN(
        n6284) );
  OAI22_X1 U50260 ( .A1(n49434), .A2(n67828), .B1(n68101), .B2(n67822), .ZN(
        n6285) );
  OAI22_X1 U50261 ( .A1(n49435), .A2(n67828), .B1(n68104), .B2(n67822), .ZN(
        n6286) );
  OAI22_X1 U50262 ( .A1(n49436), .A2(n67828), .B1(n68107), .B2(n67822), .ZN(
        n6287) );
  OAI22_X1 U50263 ( .A1(n49437), .A2(n67828), .B1(n68110), .B2(n67822), .ZN(
        n6288) );
  OAI22_X1 U50264 ( .A1(n49438), .A2(n67828), .B1(n68113), .B2(n67822), .ZN(
        n6289) );
  OAI22_X1 U50265 ( .A1(n49439), .A2(n67828), .B1(n68116), .B2(n67822), .ZN(
        n6290) );
  OAI22_X1 U50266 ( .A1(n49440), .A2(n67828), .B1(n68119), .B2(n67822), .ZN(
        n6291) );
  OAI22_X1 U50267 ( .A1(n49441), .A2(n67828), .B1(n68122), .B2(n67822), .ZN(
        n6292) );
  OAI22_X1 U50268 ( .A1(n49442), .A2(n67828), .B1(n68125), .B2(n67822), .ZN(
        n6293) );
  OAI22_X1 U50269 ( .A1(n49443), .A2(n67829), .B1(n68128), .B2(n67822), .ZN(
        n6294) );
  OAI22_X1 U50270 ( .A1(n49444), .A2(n67829), .B1(n68131), .B2(n67823), .ZN(
        n6295) );
  OAI22_X1 U50271 ( .A1(n49445), .A2(n67829), .B1(n68134), .B2(n67823), .ZN(
        n6296) );
  OAI22_X1 U50272 ( .A1(n49446), .A2(n67829), .B1(n68137), .B2(n67823), .ZN(
        n6297) );
  OAI22_X1 U50273 ( .A1(n49447), .A2(n67829), .B1(n68140), .B2(n67823), .ZN(
        n6298) );
  OAI22_X1 U50274 ( .A1(n49448), .A2(n67829), .B1(n68143), .B2(n67823), .ZN(
        n6299) );
  OAI22_X1 U50275 ( .A1(n49449), .A2(n67829), .B1(n68146), .B2(n67823), .ZN(
        n6300) );
  OAI22_X1 U50276 ( .A1(n49450), .A2(n67829), .B1(n68149), .B2(n67823), .ZN(
        n6301) );
  OAI22_X1 U50277 ( .A1(n49451), .A2(n67829), .B1(n68152), .B2(n67823), .ZN(
        n6302) );
  OAI22_X1 U50278 ( .A1(n49452), .A2(n67829), .B1(n68155), .B2(n67823), .ZN(
        n6303) );
  OAI22_X1 U50279 ( .A1(n49453), .A2(n67829), .B1(n68158), .B2(n67823), .ZN(
        n6304) );
  OAI22_X1 U50280 ( .A1(n49454), .A2(n67829), .B1(n68161), .B2(n67823), .ZN(
        n6305) );
  OAI22_X1 U50281 ( .A1(n49455), .A2(n67830), .B1(n68164), .B2(n67823), .ZN(
        n6306) );
  OAI22_X1 U50282 ( .A1(n49456), .A2(n67830), .B1(n68167), .B2(n67824), .ZN(
        n6307) );
  OAI22_X1 U50283 ( .A1(n49457), .A2(n67830), .B1(n68170), .B2(n67824), .ZN(
        n6308) );
  OAI22_X1 U50284 ( .A1(n49458), .A2(n67830), .B1(n68173), .B2(n67824), .ZN(
        n6309) );
  OAI22_X1 U50285 ( .A1(n49459), .A2(n67830), .B1(n68176), .B2(n67824), .ZN(
        n6310) );
  OAI22_X1 U50286 ( .A1(n49460), .A2(n67830), .B1(n68179), .B2(n67824), .ZN(
        n6311) );
  OAI22_X1 U50287 ( .A1(n49461), .A2(n67830), .B1(n68182), .B2(n67824), .ZN(
        n6312) );
  OAI22_X1 U50288 ( .A1(n49462), .A2(n67830), .B1(n68185), .B2(n67824), .ZN(
        n6313) );
  OAI22_X1 U50289 ( .A1(n49463), .A2(n67830), .B1(n68188), .B2(n67824), .ZN(
        n6314) );
  OAI22_X1 U50290 ( .A1(n49464), .A2(n67830), .B1(n68191), .B2(n67824), .ZN(
        n6315) );
  OAI22_X1 U50291 ( .A1(n49465), .A2(n67830), .B1(n68194), .B2(n67824), .ZN(
        n6316) );
  OAI22_X1 U50292 ( .A1(n49466), .A2(n67830), .B1(n68197), .B2(n67824), .ZN(
        n6317) );
  OAI22_X1 U50293 ( .A1(n49467), .A2(n67831), .B1(n68200), .B2(n67824), .ZN(
        n6318) );
  OAI22_X1 U50294 ( .A1(n49468), .A2(n67831), .B1(n68203), .B2(n67825), .ZN(
        n6319) );
  OAI22_X1 U50295 ( .A1(n49469), .A2(n67831), .B1(n68206), .B2(n67825), .ZN(
        n6320) );
  OAI22_X1 U50296 ( .A1(n49470), .A2(n67831), .B1(n68209), .B2(n67825), .ZN(
        n6321) );
  OAI22_X1 U50297 ( .A1(n49471), .A2(n67831), .B1(n68212), .B2(n67825), .ZN(
        n6322) );
  OAI22_X1 U50298 ( .A1(n49472), .A2(n67831), .B1(n68215), .B2(n67825), .ZN(
        n6323) );
  OAI22_X1 U50299 ( .A1(n49473), .A2(n67831), .B1(n68218), .B2(n67825), .ZN(
        n6324) );
  OAI22_X1 U50300 ( .A1(n49474), .A2(n67831), .B1(n68221), .B2(n67825), .ZN(
        n6325) );
  OAI22_X1 U50301 ( .A1(n49475), .A2(n67831), .B1(n68224), .B2(n67825), .ZN(
        n6326) );
  OAI22_X1 U50302 ( .A1(n49476), .A2(n67831), .B1(n68227), .B2(n67825), .ZN(
        n6327) );
  OAI22_X1 U50303 ( .A1(n49477), .A2(n67831), .B1(n68230), .B2(n67825), .ZN(
        n6328) );
  OAI22_X1 U50304 ( .A1(n49478), .A2(n67831), .B1(n68233), .B2(n67825), .ZN(
        n6329) );
  OAI22_X1 U50305 ( .A1(n49479), .A2(n67832), .B1(n68236), .B2(n67825), .ZN(
        n6330) );
  OAI22_X1 U50306 ( .A1(n67778), .A2(n63294), .B1(n68059), .B2(n67770), .ZN(
        n6015) );
  OAI22_X1 U50307 ( .A1(n67778), .A2(n63293), .B1(n68062), .B2(n67770), .ZN(
        n6016) );
  OAI22_X1 U50308 ( .A1(n67778), .A2(n63292), .B1(n68065), .B2(n67770), .ZN(
        n6017) );
  OAI22_X1 U50309 ( .A1(n67778), .A2(n63291), .B1(n68068), .B2(n67770), .ZN(
        n6018) );
  OAI22_X1 U50310 ( .A1(n67778), .A2(n63290), .B1(n68071), .B2(n67770), .ZN(
        n6019) );
  OAI22_X1 U50311 ( .A1(n67778), .A2(n63289), .B1(n68074), .B2(n67770), .ZN(
        n6020) );
  OAI22_X1 U50312 ( .A1(n67778), .A2(n63288), .B1(n68077), .B2(n67770), .ZN(
        n6021) );
  OAI22_X1 U50313 ( .A1(n67778), .A2(n63287), .B1(n68080), .B2(n67770), .ZN(
        n6022) );
  OAI22_X1 U50314 ( .A1(n67778), .A2(n63286), .B1(n68083), .B2(n67770), .ZN(
        n6023) );
  OAI22_X1 U50315 ( .A1(n67778), .A2(n63285), .B1(n68086), .B2(n67770), .ZN(
        n6024) );
  OAI22_X1 U50316 ( .A1(n67778), .A2(n63284), .B1(n68089), .B2(n67770), .ZN(
        n6025) );
  OAI22_X1 U50317 ( .A1(n67778), .A2(n63283), .B1(n68092), .B2(n67770), .ZN(
        n6026) );
  OAI22_X1 U50318 ( .A1(n67779), .A2(n63282), .B1(n68095), .B2(n67771), .ZN(
        n6027) );
  OAI22_X1 U50319 ( .A1(n67779), .A2(n63281), .B1(n68098), .B2(n67771), .ZN(
        n6028) );
  OAI22_X1 U50320 ( .A1(n67779), .A2(n63280), .B1(n68101), .B2(n67771), .ZN(
        n6029) );
  OAI22_X1 U50321 ( .A1(n67779), .A2(n63279), .B1(n68104), .B2(n67771), .ZN(
        n6030) );
  OAI22_X1 U50322 ( .A1(n67779), .A2(n63278), .B1(n68107), .B2(n67771), .ZN(
        n6031) );
  OAI22_X1 U50323 ( .A1(n67779), .A2(n63277), .B1(n68110), .B2(n67771), .ZN(
        n6032) );
  OAI22_X1 U50324 ( .A1(n67779), .A2(n63276), .B1(n68113), .B2(n67771), .ZN(
        n6033) );
  OAI22_X1 U50325 ( .A1(n67779), .A2(n63275), .B1(n68116), .B2(n67771), .ZN(
        n6034) );
  OAI22_X1 U50326 ( .A1(n67779), .A2(n63274), .B1(n68119), .B2(n67771), .ZN(
        n6035) );
  OAI22_X1 U50327 ( .A1(n67779), .A2(n63273), .B1(n68122), .B2(n67771), .ZN(
        n6036) );
  OAI22_X1 U50328 ( .A1(n67779), .A2(n63272), .B1(n68125), .B2(n67771), .ZN(
        n6037) );
  OAI22_X1 U50329 ( .A1(n67779), .A2(n63271), .B1(n68128), .B2(n67771), .ZN(
        n6038) );
  OAI22_X1 U50330 ( .A1(n67779), .A2(n63270), .B1(n68131), .B2(n67772), .ZN(
        n6039) );
  OAI22_X1 U50331 ( .A1(n67780), .A2(n63269), .B1(n68134), .B2(n67772), .ZN(
        n6040) );
  OAI22_X1 U50332 ( .A1(n67780), .A2(n63268), .B1(n68137), .B2(n67772), .ZN(
        n6041) );
  OAI22_X1 U50333 ( .A1(n67780), .A2(n63267), .B1(n68140), .B2(n67772), .ZN(
        n6042) );
  OAI22_X1 U50334 ( .A1(n67780), .A2(n63266), .B1(n68143), .B2(n67772), .ZN(
        n6043) );
  OAI22_X1 U50335 ( .A1(n67780), .A2(n63265), .B1(n68146), .B2(n67772), .ZN(
        n6044) );
  OAI22_X1 U50336 ( .A1(n67780), .A2(n63264), .B1(n68149), .B2(n67772), .ZN(
        n6045) );
  OAI22_X1 U50337 ( .A1(n67780), .A2(n63263), .B1(n68152), .B2(n67772), .ZN(
        n6046) );
  OAI22_X1 U50338 ( .A1(n67780), .A2(n63262), .B1(n68155), .B2(n67772), .ZN(
        n6047) );
  OAI22_X1 U50339 ( .A1(n67780), .A2(n63261), .B1(n68158), .B2(n67772), .ZN(
        n6048) );
  OAI22_X1 U50340 ( .A1(n67780), .A2(n63260), .B1(n68161), .B2(n67772), .ZN(
        n6049) );
  OAI22_X1 U50341 ( .A1(n67780), .A2(n63259), .B1(n68164), .B2(n67772), .ZN(
        n6050) );
  OAI22_X1 U50342 ( .A1(n67780), .A2(n63258), .B1(n68167), .B2(n67773), .ZN(
        n6051) );
  OAI22_X1 U50343 ( .A1(n67780), .A2(n63257), .B1(n68170), .B2(n67773), .ZN(
        n6052) );
  OAI22_X1 U50344 ( .A1(n67781), .A2(n63256), .B1(n68173), .B2(n67773), .ZN(
        n6053) );
  OAI22_X1 U50345 ( .A1(n67781), .A2(n63255), .B1(n68176), .B2(n67773), .ZN(
        n6054) );
  OAI22_X1 U50346 ( .A1(n67781), .A2(n63254), .B1(n68179), .B2(n67773), .ZN(
        n6055) );
  OAI22_X1 U50347 ( .A1(n67781), .A2(n63253), .B1(n68182), .B2(n67773), .ZN(
        n6056) );
  OAI22_X1 U50348 ( .A1(n67781), .A2(n63252), .B1(n68185), .B2(n67773), .ZN(
        n6057) );
  OAI22_X1 U50349 ( .A1(n67781), .A2(n63251), .B1(n68188), .B2(n67773), .ZN(
        n6058) );
  OAI22_X1 U50350 ( .A1(n67781), .A2(n63250), .B1(n68191), .B2(n67773), .ZN(
        n6059) );
  OAI22_X1 U50351 ( .A1(n67781), .A2(n63249), .B1(n68194), .B2(n67773), .ZN(
        n6060) );
  OAI22_X1 U50352 ( .A1(n67781), .A2(n63248), .B1(n68197), .B2(n67773), .ZN(
        n6061) );
  OAI22_X1 U50353 ( .A1(n67781), .A2(n63247), .B1(n68200), .B2(n67773), .ZN(
        n6062) );
  OAI22_X1 U50354 ( .A1(n67781), .A2(n63246), .B1(n68203), .B2(n67774), .ZN(
        n6063) );
  OAI22_X1 U50355 ( .A1(n67781), .A2(n63245), .B1(n68206), .B2(n67774), .ZN(
        n6064) );
  OAI22_X1 U50356 ( .A1(n67781), .A2(n63244), .B1(n68209), .B2(n67774), .ZN(
        n6065) );
  OAI22_X1 U50357 ( .A1(n67782), .A2(n63243), .B1(n68212), .B2(n67774), .ZN(
        n6066) );
  OAI22_X1 U50358 ( .A1(n67782), .A2(n63242), .B1(n68215), .B2(n67774), .ZN(
        n6067) );
  OAI22_X1 U50359 ( .A1(n67782), .A2(n63241), .B1(n68218), .B2(n67774), .ZN(
        n6068) );
  OAI22_X1 U50360 ( .A1(n67782), .A2(n63240), .B1(n68221), .B2(n67774), .ZN(
        n6069) );
  OAI22_X1 U50361 ( .A1(n67782), .A2(n63239), .B1(n68224), .B2(n67774), .ZN(
        n6070) );
  OAI22_X1 U50362 ( .A1(n67782), .A2(n63238), .B1(n68227), .B2(n67774), .ZN(
        n6071) );
  OAI22_X1 U50363 ( .A1(n67782), .A2(n63237), .B1(n68230), .B2(n67774), .ZN(
        n6072) );
  OAI22_X1 U50364 ( .A1(n67782), .A2(n63236), .B1(n68233), .B2(n67774), .ZN(
        n6073) );
  OAI22_X1 U50365 ( .A1(n67782), .A2(n63235), .B1(n68236), .B2(n67774), .ZN(
        n6074) );
  OAI22_X1 U50366 ( .A1(n7489), .A2(n67789), .B1(n68059), .B2(n67783), .ZN(
        n6079) );
  OAI22_X1 U50367 ( .A1(n7505), .A2(n67789), .B1(n68062), .B2(n67783), .ZN(
        n6080) );
  OAI22_X1 U50368 ( .A1(n7521), .A2(n67789), .B1(n68065), .B2(n67783), .ZN(
        n6081) );
  OAI22_X1 U50369 ( .A1(n7537), .A2(n67789), .B1(n68068), .B2(n67783), .ZN(
        n6082) );
  OAI22_X1 U50370 ( .A1(n7553), .A2(n67789), .B1(n68071), .B2(n67783), .ZN(
        n6083) );
  OAI22_X1 U50371 ( .A1(n7569), .A2(n67789), .B1(n68074), .B2(n67783), .ZN(
        n6084) );
  OAI22_X1 U50372 ( .A1(n7585), .A2(n67789), .B1(n68077), .B2(n67783), .ZN(
        n6085) );
  OAI22_X1 U50373 ( .A1(n7601), .A2(n67789), .B1(n68080), .B2(n67783), .ZN(
        n6086) );
  OAI22_X1 U50374 ( .A1(n7617), .A2(n67789), .B1(n68083), .B2(n67783), .ZN(
        n6087) );
  OAI22_X1 U50375 ( .A1(n7633), .A2(n67789), .B1(n68086), .B2(n67783), .ZN(
        n6088) );
  OAI22_X1 U50376 ( .A1(n7649), .A2(n67789), .B1(n68089), .B2(n67783), .ZN(
        n6089) );
  OAI22_X1 U50377 ( .A1(n7665), .A2(n67790), .B1(n68092), .B2(n67783), .ZN(
        n6090) );
  OAI22_X1 U50378 ( .A1(n7681), .A2(n67790), .B1(n68095), .B2(n67784), .ZN(
        n6091) );
  OAI22_X1 U50379 ( .A1(n7697), .A2(n67790), .B1(n68098), .B2(n67784), .ZN(
        n6092) );
  OAI22_X1 U50380 ( .A1(n7713), .A2(n67790), .B1(n68101), .B2(n67784), .ZN(
        n6093) );
  OAI22_X1 U50381 ( .A1(n7729), .A2(n67790), .B1(n68104), .B2(n67784), .ZN(
        n6094) );
  OAI22_X1 U50382 ( .A1(n7745), .A2(n67790), .B1(n68107), .B2(n67784), .ZN(
        n6095) );
  OAI22_X1 U50383 ( .A1(n7761), .A2(n67790), .B1(n68110), .B2(n67784), .ZN(
        n6096) );
  OAI22_X1 U50384 ( .A1(n7777), .A2(n67790), .B1(n68113), .B2(n67784), .ZN(
        n6097) );
  OAI22_X1 U50385 ( .A1(n7793), .A2(n67790), .B1(n68116), .B2(n67784), .ZN(
        n6098) );
  OAI22_X1 U50386 ( .A1(n7809), .A2(n67790), .B1(n68119), .B2(n67784), .ZN(
        n6099) );
  OAI22_X1 U50387 ( .A1(n7825), .A2(n67790), .B1(n68122), .B2(n67784), .ZN(
        n6100) );
  OAI22_X1 U50388 ( .A1(n7841), .A2(n67790), .B1(n68125), .B2(n67784), .ZN(
        n6101) );
  OAI22_X1 U50389 ( .A1(n7857), .A2(n67791), .B1(n68128), .B2(n67784), .ZN(
        n6102) );
  OAI22_X1 U50390 ( .A1(n7873), .A2(n67791), .B1(n68131), .B2(n67785), .ZN(
        n6103) );
  OAI22_X1 U50391 ( .A1(n7889), .A2(n67791), .B1(n68134), .B2(n67785), .ZN(
        n6104) );
  OAI22_X1 U50392 ( .A1(n7905), .A2(n67791), .B1(n68137), .B2(n67785), .ZN(
        n6105) );
  OAI22_X1 U50393 ( .A1(n7921), .A2(n67791), .B1(n68140), .B2(n67785), .ZN(
        n6106) );
  OAI22_X1 U50394 ( .A1(n7937), .A2(n67791), .B1(n68143), .B2(n67785), .ZN(
        n6107) );
  OAI22_X1 U50395 ( .A1(n7953), .A2(n67791), .B1(n68146), .B2(n67785), .ZN(
        n6108) );
  OAI22_X1 U50396 ( .A1(n7969), .A2(n67791), .B1(n68149), .B2(n67785), .ZN(
        n6109) );
  OAI22_X1 U50397 ( .A1(n7985), .A2(n67791), .B1(n68152), .B2(n67785), .ZN(
        n6110) );
  OAI22_X1 U50398 ( .A1(n8001), .A2(n67791), .B1(n68155), .B2(n67785), .ZN(
        n6111) );
  OAI22_X1 U50399 ( .A1(n8017), .A2(n67791), .B1(n68158), .B2(n67785), .ZN(
        n6112) );
  OAI22_X1 U50400 ( .A1(n8033), .A2(n67791), .B1(n68161), .B2(n67785), .ZN(
        n6113) );
  OAI22_X1 U50401 ( .A1(n8049), .A2(n67792), .B1(n68164), .B2(n67785), .ZN(
        n6114) );
  OAI22_X1 U50402 ( .A1(n8065), .A2(n67792), .B1(n68167), .B2(n67786), .ZN(
        n6115) );
  OAI22_X1 U50403 ( .A1(n8081), .A2(n67792), .B1(n68170), .B2(n67786), .ZN(
        n6116) );
  OAI22_X1 U50404 ( .A1(n8097), .A2(n67792), .B1(n68173), .B2(n67786), .ZN(
        n6117) );
  OAI22_X1 U50405 ( .A1(n8113), .A2(n67792), .B1(n68176), .B2(n67786), .ZN(
        n6118) );
  OAI22_X1 U50406 ( .A1(n8129), .A2(n67792), .B1(n68179), .B2(n67786), .ZN(
        n6119) );
  OAI22_X1 U50407 ( .A1(n8145), .A2(n67792), .B1(n68182), .B2(n67786), .ZN(
        n6120) );
  OAI22_X1 U50408 ( .A1(n8161), .A2(n67792), .B1(n68185), .B2(n67786), .ZN(
        n6121) );
  OAI22_X1 U50409 ( .A1(n8177), .A2(n67792), .B1(n68188), .B2(n67786), .ZN(
        n6122) );
  OAI22_X1 U50410 ( .A1(n8193), .A2(n67792), .B1(n68191), .B2(n67786), .ZN(
        n6123) );
  OAI22_X1 U50411 ( .A1(n8209), .A2(n67792), .B1(n68194), .B2(n67786), .ZN(
        n6124) );
  OAI22_X1 U50412 ( .A1(n8225), .A2(n67792), .B1(n68197), .B2(n67786), .ZN(
        n6125) );
  OAI22_X1 U50413 ( .A1(n8241), .A2(n67793), .B1(n68200), .B2(n67786), .ZN(
        n6126) );
  OAI22_X1 U50414 ( .A1(n8257), .A2(n67793), .B1(n68203), .B2(n67787), .ZN(
        n6127) );
  OAI22_X1 U50415 ( .A1(n8273), .A2(n67793), .B1(n68206), .B2(n67787), .ZN(
        n6128) );
  OAI22_X1 U50416 ( .A1(n8289), .A2(n67793), .B1(n68209), .B2(n67787), .ZN(
        n6129) );
  OAI22_X1 U50417 ( .A1(n8305), .A2(n67793), .B1(n68212), .B2(n67787), .ZN(
        n6130) );
  OAI22_X1 U50418 ( .A1(n8321), .A2(n67793), .B1(n68215), .B2(n67787), .ZN(
        n6131) );
  OAI22_X1 U50419 ( .A1(n8337), .A2(n67793), .B1(n68218), .B2(n67787), .ZN(
        n6132) );
  OAI22_X1 U50420 ( .A1(n8353), .A2(n67793), .B1(n68221), .B2(n67787), .ZN(
        n6133) );
  OAI22_X1 U50421 ( .A1(n8369), .A2(n67793), .B1(n68224), .B2(n67787), .ZN(
        n6134) );
  OAI22_X1 U50422 ( .A1(n8385), .A2(n67793), .B1(n68227), .B2(n67787), .ZN(
        n6135) );
  OAI22_X1 U50423 ( .A1(n8401), .A2(n67793), .B1(n68230), .B2(n67787), .ZN(
        n6136) );
  OAI22_X1 U50424 ( .A1(n8417), .A2(n67793), .B1(n68233), .B2(n67787), .ZN(
        n6137) );
  OAI22_X1 U50425 ( .A1(n8433), .A2(n67794), .B1(n68236), .B2(n67787), .ZN(
        n6138) );
  OAI22_X1 U50426 ( .A1(n67893), .A2(n62825), .B1(n68059), .B2(n67885), .ZN(
        n6591) );
  OAI22_X1 U50427 ( .A1(n67897), .A2(n62824), .B1(n68062), .B2(n67885), .ZN(
        n6592) );
  OAI22_X1 U50428 ( .A1(n67897), .A2(n62823), .B1(n68065), .B2(n67885), .ZN(
        n6593) );
  OAI22_X1 U50429 ( .A1(n67897), .A2(n62822), .B1(n68068), .B2(n67885), .ZN(
        n6594) );
  OAI22_X1 U50430 ( .A1(n67897), .A2(n62821), .B1(n68071), .B2(n67885), .ZN(
        n6595) );
  OAI22_X1 U50431 ( .A1(n67897), .A2(n62820), .B1(n68074), .B2(n67885), .ZN(
        n6596) );
  OAI22_X1 U50432 ( .A1(n67897), .A2(n62819), .B1(n68077), .B2(n67885), .ZN(
        n6597) );
  OAI22_X1 U50433 ( .A1(n67897), .A2(n62818), .B1(n68080), .B2(n67885), .ZN(
        n6598) );
  OAI22_X1 U50434 ( .A1(n67897), .A2(n62817), .B1(n68083), .B2(n67885), .ZN(
        n6599) );
  OAI22_X1 U50435 ( .A1(n67897), .A2(n62816), .B1(n68086), .B2(n67885), .ZN(
        n6600) );
  OAI22_X1 U50436 ( .A1(n67897), .A2(n62815), .B1(n68089), .B2(n67885), .ZN(
        n6601) );
  OAI22_X1 U50437 ( .A1(n67897), .A2(n62814), .B1(n68092), .B2(n67885), .ZN(
        n6602) );
  OAI22_X1 U50438 ( .A1(n67897), .A2(n62813), .B1(n68095), .B2(n67886), .ZN(
        n6603) );
  OAI22_X1 U50439 ( .A1(n67897), .A2(n62812), .B1(n68098), .B2(n67886), .ZN(
        n6604) );
  OAI22_X1 U50440 ( .A1(n67896), .A2(n62811), .B1(n68101), .B2(n67886), .ZN(
        n6605) );
  OAI22_X1 U50441 ( .A1(n67896), .A2(n62810), .B1(n68104), .B2(n67886), .ZN(
        n6606) );
  OAI22_X1 U50442 ( .A1(n67896), .A2(n62809), .B1(n68107), .B2(n67886), .ZN(
        n6607) );
  OAI22_X1 U50443 ( .A1(n67896), .A2(n62808), .B1(n68110), .B2(n67886), .ZN(
        n6608) );
  OAI22_X1 U50444 ( .A1(n67896), .A2(n62807), .B1(n68113), .B2(n67886), .ZN(
        n6609) );
  OAI22_X1 U50445 ( .A1(n67896), .A2(n62806), .B1(n68116), .B2(n67886), .ZN(
        n6610) );
  OAI22_X1 U50446 ( .A1(n67896), .A2(n62805), .B1(n68119), .B2(n67886), .ZN(
        n6611) );
  OAI22_X1 U50447 ( .A1(n67896), .A2(n62804), .B1(n68122), .B2(n67886), .ZN(
        n6612) );
  OAI22_X1 U50448 ( .A1(n67896), .A2(n62803), .B1(n68125), .B2(n67886), .ZN(
        n6613) );
  OAI22_X1 U50449 ( .A1(n67896), .A2(n62802), .B1(n68128), .B2(n67886), .ZN(
        n6614) );
  OAI22_X1 U50450 ( .A1(n67896), .A2(n62801), .B1(n68131), .B2(n67887), .ZN(
        n6615) );
  OAI22_X1 U50451 ( .A1(n67896), .A2(n62800), .B1(n68134), .B2(n67887), .ZN(
        n6616) );
  OAI22_X1 U50452 ( .A1(n67896), .A2(n62799), .B1(n68137), .B2(n67887), .ZN(
        n6617) );
  OAI22_X1 U50453 ( .A1(n67895), .A2(n62798), .B1(n68140), .B2(n67887), .ZN(
        n6618) );
  OAI22_X1 U50454 ( .A1(n67895), .A2(n62797), .B1(n68143), .B2(n67887), .ZN(
        n6619) );
  OAI22_X1 U50455 ( .A1(n67895), .A2(n62796), .B1(n68146), .B2(n67887), .ZN(
        n6620) );
  OAI22_X1 U50456 ( .A1(n67895), .A2(n62795), .B1(n68149), .B2(n67887), .ZN(
        n6621) );
  OAI22_X1 U50457 ( .A1(n67895), .A2(n62794), .B1(n68152), .B2(n67887), .ZN(
        n6622) );
  OAI22_X1 U50458 ( .A1(n67895), .A2(n62793), .B1(n68155), .B2(n67887), .ZN(
        n6623) );
  OAI22_X1 U50459 ( .A1(n67895), .A2(n62792), .B1(n68158), .B2(n67887), .ZN(
        n6624) );
  OAI22_X1 U50460 ( .A1(n67895), .A2(n62791), .B1(n68161), .B2(n67887), .ZN(
        n6625) );
  OAI22_X1 U50461 ( .A1(n67895), .A2(n62790), .B1(n68164), .B2(n67887), .ZN(
        n6626) );
  OAI22_X1 U50462 ( .A1(n67895), .A2(n62789), .B1(n68167), .B2(n67888), .ZN(
        n6627) );
  OAI22_X1 U50463 ( .A1(n67895), .A2(n62788), .B1(n68170), .B2(n67888), .ZN(
        n6628) );
  OAI22_X1 U50464 ( .A1(n67895), .A2(n62787), .B1(n68173), .B2(n67888), .ZN(
        n6629) );
  OAI22_X1 U50465 ( .A1(n67894), .A2(n62786), .B1(n68176), .B2(n67888), .ZN(
        n6630) );
  OAI22_X1 U50466 ( .A1(n67894), .A2(n62785), .B1(n68179), .B2(n67888), .ZN(
        n6631) );
  OAI22_X1 U50467 ( .A1(n67894), .A2(n62784), .B1(n68182), .B2(n67888), .ZN(
        n6632) );
  OAI22_X1 U50468 ( .A1(n67894), .A2(n62783), .B1(n68185), .B2(n67888), .ZN(
        n6633) );
  OAI22_X1 U50469 ( .A1(n67894), .A2(n62782), .B1(n68188), .B2(n67888), .ZN(
        n6634) );
  OAI22_X1 U50470 ( .A1(n67894), .A2(n62781), .B1(n68191), .B2(n67888), .ZN(
        n6635) );
  OAI22_X1 U50471 ( .A1(n67894), .A2(n62780), .B1(n68194), .B2(n67888), .ZN(
        n6636) );
  OAI22_X1 U50472 ( .A1(n67894), .A2(n62779), .B1(n68197), .B2(n67888), .ZN(
        n6637) );
  OAI22_X1 U50473 ( .A1(n67895), .A2(n62778), .B1(n68200), .B2(n67888), .ZN(
        n6638) );
  OAI22_X1 U50474 ( .A1(n67894), .A2(n62777), .B1(n68203), .B2(n67889), .ZN(
        n6639) );
  OAI22_X1 U50475 ( .A1(n67894), .A2(n62776), .B1(n68206), .B2(n67889), .ZN(
        n6640) );
  OAI22_X1 U50476 ( .A1(n67894), .A2(n62775), .B1(n68209), .B2(n67889), .ZN(
        n6641) );
  OAI22_X1 U50477 ( .A1(n67894), .A2(n62774), .B1(n68212), .B2(n67889), .ZN(
        n6642) );
  OAI22_X1 U50478 ( .A1(n67894), .A2(n62773), .B1(n68215), .B2(n67889), .ZN(
        n6643) );
  OAI22_X1 U50479 ( .A1(n67893), .A2(n62772), .B1(n68218), .B2(n67889), .ZN(
        n6644) );
  OAI22_X1 U50480 ( .A1(n67893), .A2(n62771), .B1(n68221), .B2(n67889), .ZN(
        n6645) );
  OAI22_X1 U50481 ( .A1(n67893), .A2(n62770), .B1(n68224), .B2(n67889), .ZN(
        n6646) );
  OAI22_X1 U50482 ( .A1(n67893), .A2(n62769), .B1(n68227), .B2(n67889), .ZN(
        n6647) );
  OAI22_X1 U50483 ( .A1(n67893), .A2(n62768), .B1(n68230), .B2(n67889), .ZN(
        n6648) );
  OAI22_X1 U50484 ( .A1(n67893), .A2(n62767), .B1(n68233), .B2(n67889), .ZN(
        n6649) );
  OAI22_X1 U50485 ( .A1(n67893), .A2(n62766), .B1(n68236), .B2(n67889), .ZN(
        n6650) );
  INV_X1 U50486 ( .A(ADD_RD2[3]), .ZN(n66292) );
  INV_X1 U50487 ( .A(ADD_RD1[3]), .ZN(n65093) );
  INV_X1 U50488 ( .A(ADD_RD2[4]), .ZN(n66291) );
  INV_X1 U50489 ( .A(ADD_RD1[4]), .ZN(n65095) );
  INV_X1 U50490 ( .A(ADD_RD2[0]), .ZN(n66297) );
  INV_X1 U50491 ( .A(ADD_RD1[0]), .ZN(n65094) );
  NAND4_X1 U50492 ( .A1(n65151), .A2(n65152), .A3(n65153), .A4(n65154), .ZN(
        n5373) );
  NOR4_X1 U50493 ( .A1(n65155), .A2(n65156), .A3(n65157), .A4(n65158), .ZN(
        n65154) );
  AOI221_X1 U50494 ( .B1(n67283), .B2(n56531), .C1(n67277), .C2(n58049), .A(
        n65168), .ZN(n65151) );
  NOR4_X1 U50495 ( .A1(n65163), .A2(n65164), .A3(n65165), .A4(n65166), .ZN(
        n65153) );
  NAND4_X1 U50496 ( .A1(n65100), .A2(n65101), .A3(n65102), .A4(n65103), .ZN(
        n5374) );
  NOR4_X1 U50497 ( .A1(n65104), .A2(n65105), .A3(n65106), .A4(n65107), .ZN(
        n65103) );
  AOI221_X1 U50498 ( .B1(n67283), .B2(n56490), .C1(n67277), .C2(n58050), .A(
        n65148), .ZN(n65100) );
  NOR4_X1 U50499 ( .A1(n65128), .A2(n65129), .A3(n65130), .A4(n65131), .ZN(
        n65102) );
  NAND4_X1 U50500 ( .A1(n66267), .A2(n66268), .A3(n66269), .A4(n66270), .ZN(
        n5311) );
  AOI221_X1 U50501 ( .B1(n67278), .B2(n58028), .C1(n67272), .C2(n58051), .A(
        n66300), .ZN(n66267) );
  NOR4_X1 U50502 ( .A1(n66293), .A2(n66294), .A3(n66295), .A4(n66296), .ZN(
        n66269) );
  AOI221_X1 U50503 ( .B1(n67302), .B2(n58731), .C1(n67296), .C2(n58283), .A(
        n66298), .ZN(n66268) );
  NAND4_X1 U50504 ( .A1(n66249), .A2(n66250), .A3(n66251), .A4(n66252), .ZN(
        n5312) );
  AOI221_X1 U50505 ( .B1(n67278), .B2(n57995), .C1(n67272), .C2(n58052), .A(
        n66266), .ZN(n66249) );
  NOR4_X1 U50506 ( .A1(n66261), .A2(n66262), .A3(n66263), .A4(n66264), .ZN(
        n66251) );
  AOI221_X1 U50507 ( .B1(n67302), .B2(n58732), .C1(n67296), .C2(n58284), .A(
        n66265), .ZN(n66250) );
  NAND4_X1 U50508 ( .A1(n66231), .A2(n66232), .A3(n66233), .A4(n66234), .ZN(
        n5313) );
  AOI221_X1 U50509 ( .B1(n67278), .B2(n57971), .C1(n67272), .C2(n58053), .A(
        n66248), .ZN(n66231) );
  NOR4_X1 U50510 ( .A1(n66243), .A2(n66244), .A3(n66245), .A4(n66246), .ZN(
        n66233) );
  AOI221_X1 U50511 ( .B1(n67302), .B2(n58733), .C1(n67296), .C2(n58285), .A(
        n66247), .ZN(n66232) );
  NAND4_X1 U50512 ( .A1(n66213), .A2(n66214), .A3(n66215), .A4(n66216), .ZN(
        n5314) );
  AOI221_X1 U50513 ( .B1(n67278), .B2(n57947), .C1(n67272), .C2(n58054), .A(
        n66230), .ZN(n66213) );
  NOR4_X1 U50514 ( .A1(n66225), .A2(n66226), .A3(n66227), .A4(n66228), .ZN(
        n66215) );
  AOI221_X1 U50515 ( .B1(n67302), .B2(n58734), .C1(n67296), .C2(n58286), .A(
        n66229), .ZN(n66214) );
  NAND4_X1 U50516 ( .A1(n66195), .A2(n66196), .A3(n66197), .A4(n66198), .ZN(
        n5315) );
  AOI221_X1 U50517 ( .B1(n67278), .B2(n57923), .C1(n67272), .C2(n58055), .A(
        n66212), .ZN(n66195) );
  NOR4_X1 U50518 ( .A1(n66207), .A2(n66208), .A3(n66209), .A4(n66210), .ZN(
        n66197) );
  AOI221_X1 U50519 ( .B1(n67302), .B2(n58735), .C1(n67296), .C2(n58287), .A(
        n66211), .ZN(n66196) );
  NAND4_X1 U50520 ( .A1(n66177), .A2(n66178), .A3(n66179), .A4(n66180), .ZN(
        n5316) );
  AOI221_X1 U50521 ( .B1(n67278), .B2(n57899), .C1(n67272), .C2(n58056), .A(
        n66194), .ZN(n66177) );
  NOR4_X1 U50522 ( .A1(n66189), .A2(n66190), .A3(n66191), .A4(n66192), .ZN(
        n66179) );
  AOI221_X1 U50523 ( .B1(n67302), .B2(n58736), .C1(n67296), .C2(n58288), .A(
        n66193), .ZN(n66178) );
  NAND4_X1 U50524 ( .A1(n66159), .A2(n66160), .A3(n66161), .A4(n66162), .ZN(
        n5317) );
  AOI221_X1 U50525 ( .B1(n67278), .B2(n57875), .C1(n67272), .C2(n58057), .A(
        n66176), .ZN(n66159) );
  NOR4_X1 U50526 ( .A1(n66171), .A2(n66172), .A3(n66173), .A4(n66174), .ZN(
        n66161) );
  AOI221_X1 U50527 ( .B1(n67302), .B2(n58737), .C1(n67296), .C2(n58289), .A(
        n66175), .ZN(n66160) );
  NAND4_X1 U50528 ( .A1(n66141), .A2(n66142), .A3(n66143), .A4(n66144), .ZN(
        n5318) );
  AOI221_X1 U50529 ( .B1(n67278), .B2(n57851), .C1(n67272), .C2(n58058), .A(
        n66158), .ZN(n66141) );
  NOR4_X1 U50530 ( .A1(n66153), .A2(n66154), .A3(n66155), .A4(n66156), .ZN(
        n66143) );
  AOI221_X1 U50531 ( .B1(n67302), .B2(n58738), .C1(n67296), .C2(n58290), .A(
        n66157), .ZN(n66142) );
  NAND4_X1 U50532 ( .A1(n66123), .A2(n66124), .A3(n66125), .A4(n66126), .ZN(
        n5319) );
  AOI221_X1 U50533 ( .B1(n67278), .B2(n57827), .C1(n67272), .C2(n58059), .A(
        n66140), .ZN(n66123) );
  NOR4_X1 U50534 ( .A1(n66135), .A2(n66136), .A3(n66137), .A4(n66138), .ZN(
        n66125) );
  AOI221_X1 U50535 ( .B1(n67302), .B2(n58739), .C1(n67296), .C2(n58291), .A(
        n66139), .ZN(n66124) );
  NAND4_X1 U50536 ( .A1(n66105), .A2(n66106), .A3(n66107), .A4(n66108), .ZN(
        n5320) );
  AOI221_X1 U50537 ( .B1(n67278), .B2(n57803), .C1(n67272), .C2(n58060), .A(
        n66122), .ZN(n66105) );
  NOR4_X1 U50538 ( .A1(n66117), .A2(n66118), .A3(n66119), .A4(n66120), .ZN(
        n66107) );
  AOI221_X1 U50539 ( .B1(n67302), .B2(n58740), .C1(n67296), .C2(n58292), .A(
        n66121), .ZN(n66106) );
  NAND4_X1 U50540 ( .A1(n66087), .A2(n66088), .A3(n66089), .A4(n66090), .ZN(
        n5321) );
  AOI221_X1 U50541 ( .B1(n67278), .B2(n57779), .C1(n67272), .C2(n58061), .A(
        n66104), .ZN(n66087) );
  NOR4_X1 U50542 ( .A1(n66099), .A2(n66100), .A3(n66101), .A4(n66102), .ZN(
        n66089) );
  AOI221_X1 U50543 ( .B1(n67302), .B2(n58741), .C1(n67296), .C2(n58293), .A(
        n66103), .ZN(n66088) );
  NAND4_X1 U50544 ( .A1(n66069), .A2(n66070), .A3(n66071), .A4(n66072), .ZN(
        n5322) );
  AOI221_X1 U50545 ( .B1(n67278), .B2(n57755), .C1(n67272), .C2(n58062), .A(
        n66086), .ZN(n66069) );
  NOR4_X1 U50546 ( .A1(n66081), .A2(n66082), .A3(n66083), .A4(n66084), .ZN(
        n66071) );
  AOI221_X1 U50547 ( .B1(n67302), .B2(n58742), .C1(n67296), .C2(n58294), .A(
        n66085), .ZN(n66070) );
  NAND4_X1 U50548 ( .A1(n66051), .A2(n66052), .A3(n66053), .A4(n66054), .ZN(
        n5323) );
  AOI221_X1 U50549 ( .B1(n67279), .B2(n57731), .C1(n67273), .C2(n58063), .A(
        n66068), .ZN(n66051) );
  NOR4_X1 U50550 ( .A1(n66063), .A2(n66064), .A3(n66065), .A4(n66066), .ZN(
        n66053) );
  AOI221_X1 U50551 ( .B1(n67303), .B2(n58667), .C1(n67297), .C2(n58235), .A(
        n66067), .ZN(n66052) );
  NAND4_X1 U50552 ( .A1(n66033), .A2(n66034), .A3(n66035), .A4(n66036), .ZN(
        n5324) );
  AOI221_X1 U50553 ( .B1(n67279), .B2(n57707), .C1(n67273), .C2(n58064), .A(
        n66050), .ZN(n66033) );
  NOR4_X1 U50554 ( .A1(n66045), .A2(n66046), .A3(n66047), .A4(n66048), .ZN(
        n66035) );
  AOI221_X1 U50555 ( .B1(n67303), .B2(n58668), .C1(n67297), .C2(n58236), .A(
        n66049), .ZN(n66034) );
  NAND4_X1 U50556 ( .A1(n66015), .A2(n66016), .A3(n66017), .A4(n66018), .ZN(
        n5325) );
  AOI221_X1 U50557 ( .B1(n67279), .B2(n57683), .C1(n67273), .C2(n58065), .A(
        n66032), .ZN(n66015) );
  NOR4_X1 U50558 ( .A1(n66027), .A2(n66028), .A3(n66029), .A4(n66030), .ZN(
        n66017) );
  AOI221_X1 U50559 ( .B1(n67303), .B2(n58669), .C1(n67297), .C2(n58237), .A(
        n66031), .ZN(n66016) );
  NAND4_X1 U50560 ( .A1(n65997), .A2(n65998), .A3(n65999), .A4(n66000), .ZN(
        n5326) );
  AOI221_X1 U50561 ( .B1(n67279), .B2(n57659), .C1(n67273), .C2(n58066), .A(
        n66014), .ZN(n65997) );
  NOR4_X1 U50562 ( .A1(n66009), .A2(n66010), .A3(n66011), .A4(n66012), .ZN(
        n65999) );
  AOI221_X1 U50563 ( .B1(n67303), .B2(n58670), .C1(n67297), .C2(n58238), .A(
        n66013), .ZN(n65998) );
  NAND4_X1 U50564 ( .A1(n65979), .A2(n65980), .A3(n65981), .A4(n65982), .ZN(
        n5327) );
  AOI221_X1 U50565 ( .B1(n67279), .B2(n57635), .C1(n67273), .C2(n58067), .A(
        n65996), .ZN(n65979) );
  NOR4_X1 U50566 ( .A1(n65991), .A2(n65992), .A3(n65993), .A4(n65994), .ZN(
        n65981) );
  AOI221_X1 U50567 ( .B1(n67303), .B2(n58671), .C1(n67297), .C2(n58239), .A(
        n65995), .ZN(n65980) );
  NAND4_X1 U50568 ( .A1(n65961), .A2(n65962), .A3(n65963), .A4(n65964), .ZN(
        n5328) );
  AOI221_X1 U50569 ( .B1(n67279), .B2(n57611), .C1(n67273), .C2(n58068), .A(
        n65978), .ZN(n65961) );
  NOR4_X1 U50570 ( .A1(n65973), .A2(n65974), .A3(n65975), .A4(n65976), .ZN(
        n65963) );
  AOI221_X1 U50571 ( .B1(n67303), .B2(n58672), .C1(n67297), .C2(n58240), .A(
        n65977), .ZN(n65962) );
  NAND4_X1 U50572 ( .A1(n65943), .A2(n65944), .A3(n65945), .A4(n65946), .ZN(
        n5329) );
  AOI221_X1 U50573 ( .B1(n67279), .B2(n57587), .C1(n67273), .C2(n58069), .A(
        n65960), .ZN(n65943) );
  NOR4_X1 U50574 ( .A1(n65955), .A2(n65956), .A3(n65957), .A4(n65958), .ZN(
        n65945) );
  AOI221_X1 U50575 ( .B1(n67303), .B2(n58673), .C1(n67297), .C2(n58241), .A(
        n65959), .ZN(n65944) );
  NAND4_X1 U50576 ( .A1(n65925), .A2(n65926), .A3(n65927), .A4(n65928), .ZN(
        n5330) );
  AOI221_X1 U50577 ( .B1(n67279), .B2(n57563), .C1(n67273), .C2(n58070), .A(
        n65942), .ZN(n65925) );
  NOR4_X1 U50578 ( .A1(n65937), .A2(n65938), .A3(n65939), .A4(n65940), .ZN(
        n65927) );
  AOI221_X1 U50579 ( .B1(n67303), .B2(n58674), .C1(n67297), .C2(n58242), .A(
        n65941), .ZN(n65926) );
  NAND4_X1 U50580 ( .A1(n65907), .A2(n65908), .A3(n65909), .A4(n65910), .ZN(
        n5331) );
  AOI221_X1 U50581 ( .B1(n67279), .B2(n57539), .C1(n67273), .C2(n58071), .A(
        n65924), .ZN(n65907) );
  NOR4_X1 U50582 ( .A1(n65919), .A2(n65920), .A3(n65921), .A4(n65922), .ZN(
        n65909) );
  AOI221_X1 U50583 ( .B1(n67303), .B2(n58675), .C1(n67297), .C2(n58243), .A(
        n65923), .ZN(n65908) );
  NAND4_X1 U50584 ( .A1(n65889), .A2(n65890), .A3(n65891), .A4(n65892), .ZN(
        n5332) );
  AOI221_X1 U50585 ( .B1(n67279), .B2(n57515), .C1(n67273), .C2(n58072), .A(
        n65906), .ZN(n65889) );
  NOR4_X1 U50586 ( .A1(n65901), .A2(n65902), .A3(n65903), .A4(n65904), .ZN(
        n65891) );
  AOI221_X1 U50587 ( .B1(n67303), .B2(n58676), .C1(n67297), .C2(n58244), .A(
        n65905), .ZN(n65890) );
  NAND4_X1 U50588 ( .A1(n65871), .A2(n65872), .A3(n65873), .A4(n65874), .ZN(
        n5333) );
  AOI221_X1 U50589 ( .B1(n67279), .B2(n57491), .C1(n67273), .C2(n58073), .A(
        n65888), .ZN(n65871) );
  NOR4_X1 U50590 ( .A1(n65883), .A2(n65884), .A3(n65885), .A4(n65886), .ZN(
        n65873) );
  AOI221_X1 U50591 ( .B1(n67303), .B2(n58677), .C1(n67297), .C2(n58245), .A(
        n65887), .ZN(n65872) );
  NAND4_X1 U50592 ( .A1(n65853), .A2(n65854), .A3(n65855), .A4(n65856), .ZN(
        n5334) );
  AOI221_X1 U50593 ( .B1(n67279), .B2(n57467), .C1(n67273), .C2(n58074), .A(
        n65870), .ZN(n65853) );
  NOR4_X1 U50594 ( .A1(n65865), .A2(n65866), .A3(n65867), .A4(n65868), .ZN(
        n65855) );
  AOI221_X1 U50595 ( .B1(n67303), .B2(n58678), .C1(n67297), .C2(n58246), .A(
        n65869), .ZN(n65854) );
  NAND4_X1 U50596 ( .A1(n65835), .A2(n65836), .A3(n65837), .A4(n65838), .ZN(
        n5335) );
  AOI221_X1 U50597 ( .B1(n67280), .B2(n57443), .C1(n67274), .C2(n58075), .A(
        n65852), .ZN(n65835) );
  NOR4_X1 U50598 ( .A1(n65847), .A2(n65848), .A3(n65849), .A4(n65850), .ZN(
        n65837) );
  AOI221_X1 U50599 ( .B1(n67304), .B2(n58679), .C1(n67298), .C2(n58247), .A(
        n65851), .ZN(n65836) );
  NAND4_X1 U50600 ( .A1(n65817), .A2(n65818), .A3(n65819), .A4(n65820), .ZN(
        n5336) );
  AOI221_X1 U50601 ( .B1(n67280), .B2(n57419), .C1(n67274), .C2(n58076), .A(
        n65834), .ZN(n65817) );
  NOR4_X1 U50602 ( .A1(n65829), .A2(n65830), .A3(n65831), .A4(n65832), .ZN(
        n65819) );
  AOI221_X1 U50603 ( .B1(n67304), .B2(n58680), .C1(n67298), .C2(n58248), .A(
        n65833), .ZN(n65818) );
  NAND4_X1 U50604 ( .A1(n65799), .A2(n65800), .A3(n65801), .A4(n65802), .ZN(
        n5337) );
  AOI221_X1 U50605 ( .B1(n67280), .B2(n57395), .C1(n67274), .C2(n58077), .A(
        n65816), .ZN(n65799) );
  NOR4_X1 U50606 ( .A1(n65811), .A2(n65812), .A3(n65813), .A4(n65814), .ZN(
        n65801) );
  AOI221_X1 U50607 ( .B1(n67304), .B2(n58681), .C1(n67298), .C2(n58249), .A(
        n65815), .ZN(n65800) );
  NAND4_X1 U50608 ( .A1(n65781), .A2(n65782), .A3(n65783), .A4(n65784), .ZN(
        n5338) );
  AOI221_X1 U50609 ( .B1(n67280), .B2(n57371), .C1(n67274), .C2(n58078), .A(
        n65798), .ZN(n65781) );
  NOR4_X1 U50610 ( .A1(n65793), .A2(n65794), .A3(n65795), .A4(n65796), .ZN(
        n65783) );
  AOI221_X1 U50611 ( .B1(n67304), .B2(n58682), .C1(n67298), .C2(n58250), .A(
        n65797), .ZN(n65782) );
  NAND4_X1 U50612 ( .A1(n65763), .A2(n65764), .A3(n65765), .A4(n65766), .ZN(
        n5339) );
  AOI221_X1 U50613 ( .B1(n67280), .B2(n57347), .C1(n67274), .C2(n58079), .A(
        n65780), .ZN(n65763) );
  NOR4_X1 U50614 ( .A1(n65775), .A2(n65776), .A3(n65777), .A4(n65778), .ZN(
        n65765) );
  AOI221_X1 U50615 ( .B1(n67304), .B2(n58683), .C1(n67298), .C2(n58251), .A(
        n65779), .ZN(n65764) );
  NAND4_X1 U50616 ( .A1(n65745), .A2(n65746), .A3(n65747), .A4(n65748), .ZN(
        n5340) );
  AOI221_X1 U50617 ( .B1(n67280), .B2(n57323), .C1(n67274), .C2(n58080), .A(
        n65762), .ZN(n65745) );
  NOR4_X1 U50618 ( .A1(n65757), .A2(n65758), .A3(n65759), .A4(n65760), .ZN(
        n65747) );
  AOI221_X1 U50619 ( .B1(n67304), .B2(n58684), .C1(n67298), .C2(n58252), .A(
        n65761), .ZN(n65746) );
  NAND4_X1 U50620 ( .A1(n65727), .A2(n65728), .A3(n65729), .A4(n65730), .ZN(
        n5341) );
  AOI221_X1 U50621 ( .B1(n67280), .B2(n57299), .C1(n67274), .C2(n58081), .A(
        n65744), .ZN(n65727) );
  NOR4_X1 U50622 ( .A1(n65739), .A2(n65740), .A3(n65741), .A4(n65742), .ZN(
        n65729) );
  AOI221_X1 U50623 ( .B1(n67304), .B2(n58685), .C1(n67298), .C2(n58253), .A(
        n65743), .ZN(n65728) );
  NAND4_X1 U50624 ( .A1(n65709), .A2(n65710), .A3(n65711), .A4(n65712), .ZN(
        n5342) );
  AOI221_X1 U50625 ( .B1(n67280), .B2(n57275), .C1(n67274), .C2(n58082), .A(
        n65726), .ZN(n65709) );
  NOR4_X1 U50626 ( .A1(n65721), .A2(n65722), .A3(n65723), .A4(n65724), .ZN(
        n65711) );
  AOI221_X1 U50627 ( .B1(n67304), .B2(n58686), .C1(n67298), .C2(n58254), .A(
        n65725), .ZN(n65710) );
  NAND4_X1 U50628 ( .A1(n65691), .A2(n65692), .A3(n65693), .A4(n65694), .ZN(
        n5343) );
  AOI221_X1 U50629 ( .B1(n67280), .B2(n57251), .C1(n67274), .C2(n58083), .A(
        n65708), .ZN(n65691) );
  NOR4_X1 U50630 ( .A1(n65703), .A2(n65704), .A3(n65705), .A4(n65706), .ZN(
        n65693) );
  AOI221_X1 U50631 ( .B1(n67304), .B2(n58687), .C1(n67298), .C2(n58255), .A(
        n65707), .ZN(n65692) );
  NAND4_X1 U50632 ( .A1(n65673), .A2(n65674), .A3(n65675), .A4(n65676), .ZN(
        n5344) );
  AOI221_X1 U50633 ( .B1(n67280), .B2(n57227), .C1(n67274), .C2(n58084), .A(
        n65690), .ZN(n65673) );
  NOR4_X1 U50634 ( .A1(n65685), .A2(n65686), .A3(n65687), .A4(n65688), .ZN(
        n65675) );
  AOI221_X1 U50635 ( .B1(n67304), .B2(n58688), .C1(n67298), .C2(n58256), .A(
        n65689), .ZN(n65674) );
  NAND4_X1 U50636 ( .A1(n65655), .A2(n65656), .A3(n65657), .A4(n65658), .ZN(
        n5345) );
  AOI221_X1 U50637 ( .B1(n67280), .B2(n57203), .C1(n67274), .C2(n58085), .A(
        n65672), .ZN(n65655) );
  NOR4_X1 U50638 ( .A1(n65667), .A2(n65668), .A3(n65669), .A4(n65670), .ZN(
        n65657) );
  AOI221_X1 U50639 ( .B1(n67304), .B2(n58689), .C1(n67298), .C2(n58257), .A(
        n65671), .ZN(n65656) );
  NAND4_X1 U50640 ( .A1(n65637), .A2(n65638), .A3(n65639), .A4(n65640), .ZN(
        n5346) );
  AOI221_X1 U50641 ( .B1(n67280), .B2(n57179), .C1(n67274), .C2(n58086), .A(
        n65654), .ZN(n65637) );
  NOR4_X1 U50642 ( .A1(n65649), .A2(n65650), .A3(n65651), .A4(n65652), .ZN(
        n65639) );
  AOI221_X1 U50643 ( .B1(n67304), .B2(n58690), .C1(n67298), .C2(n58258), .A(
        n65653), .ZN(n65638) );
  NAND4_X1 U50644 ( .A1(n65619), .A2(n65620), .A3(n65621), .A4(n65622), .ZN(
        n5347) );
  AOI221_X1 U50645 ( .B1(n67281), .B2(n57155), .C1(n67275), .C2(n58087), .A(
        n65636), .ZN(n65619) );
  NOR4_X1 U50646 ( .A1(n65631), .A2(n65632), .A3(n65633), .A4(n65634), .ZN(
        n65621) );
  AOI221_X1 U50647 ( .B1(n67305), .B2(n58691), .C1(n67299), .C2(n58259), .A(
        n65635), .ZN(n65620) );
  NAND4_X1 U50648 ( .A1(n65601), .A2(n65602), .A3(n65603), .A4(n65604), .ZN(
        n5348) );
  AOI221_X1 U50649 ( .B1(n67281), .B2(n57131), .C1(n67275), .C2(n58088), .A(
        n65618), .ZN(n65601) );
  NOR4_X1 U50650 ( .A1(n65613), .A2(n65614), .A3(n65615), .A4(n65616), .ZN(
        n65603) );
  AOI221_X1 U50651 ( .B1(n67305), .B2(n58692), .C1(n67299), .C2(n58260), .A(
        n65617), .ZN(n65602) );
  NAND4_X1 U50652 ( .A1(n65583), .A2(n65584), .A3(n65585), .A4(n65586), .ZN(
        n5349) );
  AOI221_X1 U50653 ( .B1(n67281), .B2(n57107), .C1(n67275), .C2(n58089), .A(
        n65600), .ZN(n65583) );
  NOR4_X1 U50654 ( .A1(n65595), .A2(n65596), .A3(n65597), .A4(n65598), .ZN(
        n65585) );
  AOI221_X1 U50655 ( .B1(n67305), .B2(n58693), .C1(n67299), .C2(n58261), .A(
        n65599), .ZN(n65584) );
  NAND4_X1 U50656 ( .A1(n65565), .A2(n65566), .A3(n65567), .A4(n65568), .ZN(
        n5350) );
  AOI221_X1 U50657 ( .B1(n67281), .B2(n57083), .C1(n67275), .C2(n58090), .A(
        n65582), .ZN(n65565) );
  NOR4_X1 U50658 ( .A1(n65577), .A2(n65578), .A3(n65579), .A4(n65580), .ZN(
        n65567) );
  AOI221_X1 U50659 ( .B1(n67305), .B2(n58694), .C1(n67299), .C2(n58262), .A(
        n65581), .ZN(n65566) );
  NAND4_X1 U50660 ( .A1(n65547), .A2(n65548), .A3(n65549), .A4(n65550), .ZN(
        n5351) );
  AOI221_X1 U50661 ( .B1(n67281), .B2(n57059), .C1(n67275), .C2(n58091), .A(
        n65564), .ZN(n65547) );
  NOR4_X1 U50662 ( .A1(n65559), .A2(n65560), .A3(n65561), .A4(n65562), .ZN(
        n65549) );
  AOI221_X1 U50663 ( .B1(n67305), .B2(n58695), .C1(n67299), .C2(n58263), .A(
        n65563), .ZN(n65548) );
  NAND4_X1 U50664 ( .A1(n65529), .A2(n65530), .A3(n65531), .A4(n65532), .ZN(
        n5352) );
  AOI221_X1 U50665 ( .B1(n67281), .B2(n57035), .C1(n67275), .C2(n58092), .A(
        n65546), .ZN(n65529) );
  NOR4_X1 U50666 ( .A1(n65541), .A2(n65542), .A3(n65543), .A4(n65544), .ZN(
        n65531) );
  AOI221_X1 U50667 ( .B1(n67305), .B2(n58696), .C1(n67299), .C2(n58264), .A(
        n65545), .ZN(n65530) );
  NAND4_X1 U50668 ( .A1(n65511), .A2(n65512), .A3(n65513), .A4(n65514), .ZN(
        n5353) );
  AOI221_X1 U50669 ( .B1(n67281), .B2(n57011), .C1(n67275), .C2(n58093), .A(
        n65528), .ZN(n65511) );
  NOR4_X1 U50670 ( .A1(n65523), .A2(n65524), .A3(n65525), .A4(n65526), .ZN(
        n65513) );
  AOI221_X1 U50671 ( .B1(n67305), .B2(n58697), .C1(n67299), .C2(n58265), .A(
        n65527), .ZN(n65512) );
  NAND4_X1 U50672 ( .A1(n65493), .A2(n65494), .A3(n65495), .A4(n65496), .ZN(
        n5354) );
  AOI221_X1 U50673 ( .B1(n67281), .B2(n56987), .C1(n67275), .C2(n58094), .A(
        n65510), .ZN(n65493) );
  NOR4_X1 U50674 ( .A1(n65505), .A2(n65506), .A3(n65507), .A4(n65508), .ZN(
        n65495) );
  AOI221_X1 U50675 ( .B1(n67305), .B2(n58698), .C1(n67299), .C2(n58266), .A(
        n65509), .ZN(n65494) );
  NAND4_X1 U50676 ( .A1(n65475), .A2(n65476), .A3(n65477), .A4(n65478), .ZN(
        n5355) );
  AOI221_X1 U50677 ( .B1(n67281), .B2(n56963), .C1(n67275), .C2(n58095), .A(
        n65492), .ZN(n65475) );
  NOR4_X1 U50678 ( .A1(n65487), .A2(n65488), .A3(n65489), .A4(n65490), .ZN(
        n65477) );
  AOI221_X1 U50679 ( .B1(n67305), .B2(n58699), .C1(n67299), .C2(n58267), .A(
        n65491), .ZN(n65476) );
  NAND4_X1 U50680 ( .A1(n65457), .A2(n65458), .A3(n65459), .A4(n65460), .ZN(
        n5356) );
  AOI221_X1 U50681 ( .B1(n67281), .B2(n56939), .C1(n67275), .C2(n58096), .A(
        n65474), .ZN(n65457) );
  NOR4_X1 U50682 ( .A1(n65469), .A2(n65470), .A3(n65471), .A4(n65472), .ZN(
        n65459) );
  AOI221_X1 U50683 ( .B1(n67305), .B2(n58700), .C1(n67299), .C2(n58268), .A(
        n65473), .ZN(n65458) );
  NAND4_X1 U50684 ( .A1(n65439), .A2(n65440), .A3(n65441), .A4(n65442), .ZN(
        n5357) );
  AOI221_X1 U50685 ( .B1(n67281), .B2(n56915), .C1(n67275), .C2(n58097), .A(
        n65456), .ZN(n65439) );
  NOR4_X1 U50686 ( .A1(n65451), .A2(n65452), .A3(n65453), .A4(n65454), .ZN(
        n65441) );
  AOI221_X1 U50687 ( .B1(n67305), .B2(n58701), .C1(n67299), .C2(n58269), .A(
        n65455), .ZN(n65440) );
  NAND4_X1 U50688 ( .A1(n65421), .A2(n65422), .A3(n65423), .A4(n65424), .ZN(
        n5358) );
  AOI221_X1 U50689 ( .B1(n67281), .B2(n56891), .C1(n67275), .C2(n58098), .A(
        n65438), .ZN(n65421) );
  NOR4_X1 U50690 ( .A1(n65433), .A2(n65434), .A3(n65435), .A4(n65436), .ZN(
        n65423) );
  AOI221_X1 U50691 ( .B1(n67305), .B2(n58702), .C1(n67299), .C2(n58270), .A(
        n65437), .ZN(n65422) );
  NAND4_X1 U50692 ( .A1(n65403), .A2(n65404), .A3(n65405), .A4(n65406), .ZN(
        n5359) );
  AOI221_X1 U50693 ( .B1(n67282), .B2(n56867), .C1(n67276), .C2(n58099), .A(
        n65420), .ZN(n65403) );
  NOR4_X1 U50694 ( .A1(n65415), .A2(n65416), .A3(n65417), .A4(n65418), .ZN(
        n65405) );
  AOI221_X1 U50695 ( .B1(n67306), .B2(n58703), .C1(n67300), .C2(n58271), .A(
        n65419), .ZN(n65404) );
  NAND4_X1 U50696 ( .A1(n65385), .A2(n65386), .A3(n65387), .A4(n65388), .ZN(
        n5360) );
  AOI221_X1 U50697 ( .B1(n67282), .B2(n56843), .C1(n67276), .C2(n58100), .A(
        n65402), .ZN(n65385) );
  NOR4_X1 U50698 ( .A1(n65397), .A2(n65398), .A3(n65399), .A4(n65400), .ZN(
        n65387) );
  AOI221_X1 U50699 ( .B1(n67306), .B2(n58704), .C1(n67300), .C2(n58272), .A(
        n65401), .ZN(n65386) );
  NAND4_X1 U50700 ( .A1(n65367), .A2(n65368), .A3(n65369), .A4(n65370), .ZN(
        n5361) );
  AOI221_X1 U50701 ( .B1(n67282), .B2(n56819), .C1(n67276), .C2(n58101), .A(
        n65384), .ZN(n65367) );
  NOR4_X1 U50702 ( .A1(n65379), .A2(n65380), .A3(n65381), .A4(n65382), .ZN(
        n65369) );
  AOI221_X1 U50703 ( .B1(n67306), .B2(n58705), .C1(n67300), .C2(n58273), .A(
        n65383), .ZN(n65368) );
  NAND4_X1 U50704 ( .A1(n65349), .A2(n65350), .A3(n65351), .A4(n65352), .ZN(
        n5362) );
  AOI221_X1 U50705 ( .B1(n67282), .B2(n56795), .C1(n67276), .C2(n58102), .A(
        n65366), .ZN(n65349) );
  NOR4_X1 U50706 ( .A1(n65361), .A2(n65362), .A3(n65363), .A4(n65364), .ZN(
        n65351) );
  AOI221_X1 U50707 ( .B1(n67306), .B2(n58706), .C1(n67300), .C2(n58274), .A(
        n65365), .ZN(n65350) );
  NAND4_X1 U50708 ( .A1(n65331), .A2(n65332), .A3(n65333), .A4(n65334), .ZN(
        n5363) );
  AOI221_X1 U50709 ( .B1(n67282), .B2(n56771), .C1(n67276), .C2(n58103), .A(
        n65348), .ZN(n65331) );
  NOR4_X1 U50710 ( .A1(n65343), .A2(n65344), .A3(n65345), .A4(n65346), .ZN(
        n65333) );
  AOI221_X1 U50711 ( .B1(n67306), .B2(n58707), .C1(n67300), .C2(n58275), .A(
        n65347), .ZN(n65332) );
  NAND4_X1 U50712 ( .A1(n65313), .A2(n65314), .A3(n65315), .A4(n65316), .ZN(
        n5364) );
  AOI221_X1 U50713 ( .B1(n67282), .B2(n56747), .C1(n67276), .C2(n58104), .A(
        n65330), .ZN(n65313) );
  NOR4_X1 U50714 ( .A1(n65325), .A2(n65326), .A3(n65327), .A4(n65328), .ZN(
        n65315) );
  AOI221_X1 U50715 ( .B1(n67306), .B2(n58708), .C1(n67300), .C2(n58276), .A(
        n65329), .ZN(n65314) );
  NAND4_X1 U50716 ( .A1(n65295), .A2(n65296), .A3(n65297), .A4(n65298), .ZN(
        n5365) );
  AOI221_X1 U50717 ( .B1(n67282), .B2(n56723), .C1(n67276), .C2(n58105), .A(
        n65312), .ZN(n65295) );
  NOR4_X1 U50718 ( .A1(n65307), .A2(n65308), .A3(n65309), .A4(n65310), .ZN(
        n65297) );
  AOI221_X1 U50719 ( .B1(n67306), .B2(n58709), .C1(n67300), .C2(n58277), .A(
        n65311), .ZN(n65296) );
  NAND4_X1 U50720 ( .A1(n65277), .A2(n65278), .A3(n65279), .A4(n65280), .ZN(
        n5366) );
  AOI221_X1 U50721 ( .B1(n67282), .B2(n56699), .C1(n67276), .C2(n58106), .A(
        n65294), .ZN(n65277) );
  NOR4_X1 U50722 ( .A1(n65289), .A2(n65290), .A3(n65291), .A4(n65292), .ZN(
        n65279) );
  AOI221_X1 U50723 ( .B1(n67306), .B2(n58710), .C1(n67300), .C2(n58278), .A(
        n65293), .ZN(n65278) );
  NAND4_X1 U50724 ( .A1(n65259), .A2(n65260), .A3(n65261), .A4(n65262), .ZN(
        n5367) );
  AOI221_X1 U50725 ( .B1(n67282), .B2(n56675), .C1(n67276), .C2(n58107), .A(
        n65276), .ZN(n65259) );
  NOR4_X1 U50726 ( .A1(n65271), .A2(n65272), .A3(n65273), .A4(n65274), .ZN(
        n65261) );
  AOI221_X1 U50727 ( .B1(n67306), .B2(n58711), .C1(n67300), .C2(n58279), .A(
        n65275), .ZN(n65260) );
  NAND4_X1 U50728 ( .A1(n65241), .A2(n65242), .A3(n65243), .A4(n65244), .ZN(
        n5368) );
  AOI221_X1 U50729 ( .B1(n67282), .B2(n56651), .C1(n67276), .C2(n58108), .A(
        n65258), .ZN(n65241) );
  NOR4_X1 U50730 ( .A1(n65253), .A2(n65254), .A3(n65255), .A4(n65256), .ZN(
        n65243) );
  AOI221_X1 U50731 ( .B1(n67306), .B2(n58712), .C1(n67300), .C2(n58280), .A(
        n65257), .ZN(n65242) );
  NAND4_X1 U50732 ( .A1(n65223), .A2(n65224), .A3(n65225), .A4(n65226), .ZN(
        n5369) );
  AOI221_X1 U50733 ( .B1(n67282), .B2(n56627), .C1(n67276), .C2(n58109), .A(
        n65240), .ZN(n65223) );
  NOR4_X1 U50734 ( .A1(n65235), .A2(n65236), .A3(n65237), .A4(n65238), .ZN(
        n65225) );
  AOI221_X1 U50735 ( .B1(n67306), .B2(n58713), .C1(n67300), .C2(n58281), .A(
        n65239), .ZN(n65224) );
  NAND4_X1 U50736 ( .A1(n65205), .A2(n65206), .A3(n65207), .A4(n65208), .ZN(
        n5370) );
  AOI221_X1 U50737 ( .B1(n67282), .B2(n56603), .C1(n67276), .C2(n58110), .A(
        n65222), .ZN(n65205) );
  NOR4_X1 U50738 ( .A1(n65217), .A2(n65218), .A3(n65219), .A4(n65220), .ZN(
        n65207) );
  AOI221_X1 U50739 ( .B1(n67306), .B2(n58714), .C1(n67300), .C2(n58282), .A(
        n65221), .ZN(n65206) );
  NAND4_X1 U50740 ( .A1(n65187), .A2(n65188), .A3(n65189), .A4(n65190), .ZN(
        n5371) );
  NOR4_X1 U50741 ( .A1(n65191), .A2(n65192), .A3(n65193), .A4(n65194), .ZN(
        n65190) );
  AOI221_X1 U50742 ( .B1(n67283), .B2(n56579), .C1(n67277), .C2(n58047), .A(
        n65204), .ZN(n65187) );
  NOR4_X1 U50743 ( .A1(n65199), .A2(n65200), .A3(n65201), .A4(n65202), .ZN(
        n65189) );
  NAND4_X1 U50744 ( .A1(n65169), .A2(n65170), .A3(n65171), .A4(n65172), .ZN(
        n5372) );
  NOR4_X1 U50745 ( .A1(n65173), .A2(n65174), .A3(n65175), .A4(n65176), .ZN(
        n65172) );
  AOI221_X1 U50746 ( .B1(n67283), .B2(n56555), .C1(n67277), .C2(n58048), .A(
        n65186), .ZN(n65169) );
  NOR4_X1 U50747 ( .A1(n65181), .A2(n65182), .A3(n65183), .A4(n65184), .ZN(
        n65171) );
  NAND4_X1 U50748 ( .A1(n65064), .A2(n65065), .A3(n65066), .A4(n65067), .ZN(
        n5375) );
  AOI221_X1 U50749 ( .B1(n67476), .B2(n58028), .C1(n67470), .C2(n59029), .A(
        n65098), .ZN(n65064) );
  AOI221_X1 U50750 ( .B1(n67500), .B2(n66313), .C1(n67494), .C2(n58112), .A(
        n65096), .ZN(n65065) );
  NOR4_X1 U50751 ( .A1(n65089), .A2(n65090), .A3(n65091), .A4(n65092), .ZN(
        n65066) );
  NAND4_X1 U50752 ( .A1(n65044), .A2(n65045), .A3(n65046), .A4(n65047), .ZN(
        n5377) );
  AOI221_X1 U50753 ( .B1(n67476), .B2(n57995), .C1(n67470), .C2(n59030), .A(
        n65062), .ZN(n65044) );
  AOI221_X1 U50754 ( .B1(n67500), .B2(n66314), .C1(n67494), .C2(n58114), .A(
        n65061), .ZN(n65045) );
  NOR4_X1 U50755 ( .A1(n65057), .A2(n65058), .A3(n65059), .A4(n65060), .ZN(
        n65046) );
  NAND4_X1 U50756 ( .A1(n65024), .A2(n65025), .A3(n65026), .A4(n65027), .ZN(
        n5379) );
  AOI221_X1 U50757 ( .B1(n67476), .B2(n57971), .C1(n67470), .C2(n59031), .A(
        n65042), .ZN(n65024) );
  AOI221_X1 U50758 ( .B1(n67500), .B2(n66315), .C1(n67494), .C2(n58116), .A(
        n65041), .ZN(n65025) );
  NOR4_X1 U50759 ( .A1(n65037), .A2(n65038), .A3(n65039), .A4(n65040), .ZN(
        n65026) );
  NAND4_X1 U50760 ( .A1(n65004), .A2(n65005), .A3(n65006), .A4(n65007), .ZN(
        n5381) );
  AOI221_X1 U50761 ( .B1(n67476), .B2(n57947), .C1(n67470), .C2(n59032), .A(
        n65022), .ZN(n65004) );
  AOI221_X1 U50762 ( .B1(n67500), .B2(n66316), .C1(n67494), .C2(n58118), .A(
        n65021), .ZN(n65005) );
  NOR4_X1 U50763 ( .A1(n65017), .A2(n65018), .A3(n65019), .A4(n65020), .ZN(
        n65006) );
  NAND4_X1 U50764 ( .A1(n64984), .A2(n64985), .A3(n64986), .A4(n64987), .ZN(
        n5383) );
  AOI221_X1 U50765 ( .B1(n67476), .B2(n57923), .C1(n67470), .C2(n59033), .A(
        n65002), .ZN(n64984) );
  AOI221_X1 U50766 ( .B1(n67500), .B2(n66317), .C1(n67494), .C2(n58120), .A(
        n65001), .ZN(n64985) );
  NOR4_X1 U50767 ( .A1(n64997), .A2(n64998), .A3(n64999), .A4(n65000), .ZN(
        n64986) );
  NAND4_X1 U50768 ( .A1(n64964), .A2(n64965), .A3(n64966), .A4(n64967), .ZN(
        n5385) );
  AOI221_X1 U50769 ( .B1(n67476), .B2(n57899), .C1(n67470), .C2(n59034), .A(
        n64982), .ZN(n64964) );
  AOI221_X1 U50770 ( .B1(n67500), .B2(n66318), .C1(n67494), .C2(n58122), .A(
        n64981), .ZN(n64965) );
  NOR4_X1 U50771 ( .A1(n64977), .A2(n64978), .A3(n64979), .A4(n64980), .ZN(
        n64966) );
  NAND4_X1 U50772 ( .A1(n64944), .A2(n64945), .A3(n64946), .A4(n64947), .ZN(
        n5387) );
  AOI221_X1 U50773 ( .B1(n67476), .B2(n57875), .C1(n67470), .C2(n59035), .A(
        n64962), .ZN(n64944) );
  AOI221_X1 U50774 ( .B1(n67500), .B2(n66319), .C1(n67494), .C2(n58124), .A(
        n64961), .ZN(n64945) );
  NOR4_X1 U50775 ( .A1(n64957), .A2(n64958), .A3(n64959), .A4(n64960), .ZN(
        n64946) );
  NAND4_X1 U50776 ( .A1(n64924), .A2(n64925), .A3(n64926), .A4(n64927), .ZN(
        n5389) );
  AOI221_X1 U50777 ( .B1(n67476), .B2(n57851), .C1(n67470), .C2(n59036), .A(
        n64942), .ZN(n64924) );
  AOI221_X1 U50778 ( .B1(n67500), .B2(n66320), .C1(n67494), .C2(n58126), .A(
        n64941), .ZN(n64925) );
  NOR4_X1 U50779 ( .A1(n64937), .A2(n64938), .A3(n64939), .A4(n64940), .ZN(
        n64926) );
  NAND4_X1 U50780 ( .A1(n64904), .A2(n64905), .A3(n64906), .A4(n64907), .ZN(
        n5391) );
  AOI221_X1 U50781 ( .B1(n67476), .B2(n57827), .C1(n67470), .C2(n59037), .A(
        n64922), .ZN(n64904) );
  AOI221_X1 U50782 ( .B1(n67500), .B2(n66321), .C1(n67494), .C2(n58128), .A(
        n64921), .ZN(n64905) );
  NOR4_X1 U50783 ( .A1(n64917), .A2(n64918), .A3(n64919), .A4(n64920), .ZN(
        n64906) );
  NAND4_X1 U50784 ( .A1(n64884), .A2(n64885), .A3(n64886), .A4(n64887), .ZN(
        n5393) );
  AOI221_X1 U50785 ( .B1(n67476), .B2(n57803), .C1(n67470), .C2(n59038), .A(
        n64902), .ZN(n64884) );
  AOI221_X1 U50786 ( .B1(n67500), .B2(n66322), .C1(n67494), .C2(n58130), .A(
        n64901), .ZN(n64885) );
  NOR4_X1 U50787 ( .A1(n64897), .A2(n64898), .A3(n64899), .A4(n64900), .ZN(
        n64886) );
  NAND4_X1 U50788 ( .A1(n64864), .A2(n64865), .A3(n64866), .A4(n64867), .ZN(
        n5395) );
  AOI221_X1 U50789 ( .B1(n67476), .B2(n57779), .C1(n67470), .C2(n59039), .A(
        n64882), .ZN(n64864) );
  AOI221_X1 U50790 ( .B1(n67500), .B2(n66323), .C1(n67494), .C2(n58132), .A(
        n64881), .ZN(n64865) );
  NOR4_X1 U50791 ( .A1(n64877), .A2(n64878), .A3(n64879), .A4(n64880), .ZN(
        n64866) );
  NAND4_X1 U50792 ( .A1(n64844), .A2(n64845), .A3(n64846), .A4(n64847), .ZN(
        n5397) );
  AOI221_X1 U50793 ( .B1(n67476), .B2(n57755), .C1(n67470), .C2(n59040), .A(
        n64862), .ZN(n64844) );
  AOI221_X1 U50794 ( .B1(n67500), .B2(n66324), .C1(n67494), .C2(n58134), .A(
        n64861), .ZN(n64845) );
  NOR4_X1 U50795 ( .A1(n64857), .A2(n64858), .A3(n64859), .A4(n64860), .ZN(
        n64846) );
  NAND4_X1 U50796 ( .A1(n64824), .A2(n64825), .A3(n64826), .A4(n64827), .ZN(
        n5399) );
  AOI221_X1 U50797 ( .B1(n67477), .B2(n57731), .C1(n67471), .C2(n59041), .A(
        n64842), .ZN(n64824) );
  AOI221_X1 U50798 ( .B1(n67501), .B2(n66325), .C1(n67495), .C2(n58135), .A(
        n64841), .ZN(n64825) );
  NOR4_X1 U50799 ( .A1(n64837), .A2(n64838), .A3(n64839), .A4(n64840), .ZN(
        n64826) );
  NAND4_X1 U50800 ( .A1(n64804), .A2(n64805), .A3(n64806), .A4(n64807), .ZN(
        n5401) );
  AOI221_X1 U50801 ( .B1(n67477), .B2(n57707), .C1(n67471), .C2(n59042), .A(
        n64822), .ZN(n64804) );
  AOI221_X1 U50802 ( .B1(n67501), .B2(n66326), .C1(n67495), .C2(n58137), .A(
        n64821), .ZN(n64805) );
  NOR4_X1 U50803 ( .A1(n64817), .A2(n64818), .A3(n64819), .A4(n64820), .ZN(
        n64806) );
  NAND4_X1 U50804 ( .A1(n64784), .A2(n64785), .A3(n64786), .A4(n64787), .ZN(
        n5403) );
  AOI221_X1 U50805 ( .B1(n67477), .B2(n57683), .C1(n67471), .C2(n59043), .A(
        n64802), .ZN(n64784) );
  AOI221_X1 U50806 ( .B1(n67501), .B2(n66327), .C1(n67495), .C2(n58139), .A(
        n64801), .ZN(n64785) );
  NOR4_X1 U50807 ( .A1(n64797), .A2(n64798), .A3(n64799), .A4(n64800), .ZN(
        n64786) );
  NAND4_X1 U50808 ( .A1(n64764), .A2(n64765), .A3(n64766), .A4(n64767), .ZN(
        n5405) );
  AOI221_X1 U50809 ( .B1(n67477), .B2(n57659), .C1(n67471), .C2(n59044), .A(
        n64782), .ZN(n64764) );
  AOI221_X1 U50810 ( .B1(n67501), .B2(n66328), .C1(n67495), .C2(n58141), .A(
        n64781), .ZN(n64765) );
  NOR4_X1 U50811 ( .A1(n64777), .A2(n64778), .A3(n64779), .A4(n64780), .ZN(
        n64766) );
  NAND4_X1 U50812 ( .A1(n64744), .A2(n64745), .A3(n64746), .A4(n64747), .ZN(
        n5407) );
  AOI221_X1 U50813 ( .B1(n67477), .B2(n57635), .C1(n67471), .C2(n59045), .A(
        n64762), .ZN(n64744) );
  AOI221_X1 U50814 ( .B1(n67501), .B2(n66329), .C1(n67495), .C2(n58143), .A(
        n64761), .ZN(n64745) );
  NOR4_X1 U50815 ( .A1(n64757), .A2(n64758), .A3(n64759), .A4(n64760), .ZN(
        n64746) );
  NAND4_X1 U50816 ( .A1(n64724), .A2(n64725), .A3(n64726), .A4(n64727), .ZN(
        n5409) );
  AOI221_X1 U50817 ( .B1(n67477), .B2(n57611), .C1(n67471), .C2(n59046), .A(
        n64742), .ZN(n64724) );
  AOI221_X1 U50818 ( .B1(n67501), .B2(n66330), .C1(n67495), .C2(n58145), .A(
        n64741), .ZN(n64725) );
  NOR4_X1 U50819 ( .A1(n64737), .A2(n64738), .A3(n64739), .A4(n64740), .ZN(
        n64726) );
  NAND4_X1 U50820 ( .A1(n64704), .A2(n64705), .A3(n64706), .A4(n64707), .ZN(
        n5411) );
  AOI221_X1 U50821 ( .B1(n67477), .B2(n57587), .C1(n67471), .C2(n59047), .A(
        n64722), .ZN(n64704) );
  AOI221_X1 U50822 ( .B1(n67501), .B2(n66331), .C1(n67495), .C2(n58147), .A(
        n64721), .ZN(n64705) );
  NOR4_X1 U50823 ( .A1(n64717), .A2(n64718), .A3(n64719), .A4(n64720), .ZN(
        n64706) );
  NAND4_X1 U50824 ( .A1(n64684), .A2(n64685), .A3(n64686), .A4(n64687), .ZN(
        n5413) );
  AOI221_X1 U50825 ( .B1(n67477), .B2(n57563), .C1(n67471), .C2(n59048), .A(
        n64702), .ZN(n64684) );
  AOI221_X1 U50826 ( .B1(n67501), .B2(n66332), .C1(n67495), .C2(n58149), .A(
        n64701), .ZN(n64685) );
  NOR4_X1 U50827 ( .A1(n64697), .A2(n64698), .A3(n64699), .A4(n64700), .ZN(
        n64686) );
  NAND4_X1 U50828 ( .A1(n64664), .A2(n64665), .A3(n64666), .A4(n64667), .ZN(
        n5415) );
  AOI221_X1 U50829 ( .B1(n67477), .B2(n57539), .C1(n67471), .C2(n59049), .A(
        n64682), .ZN(n64664) );
  AOI221_X1 U50830 ( .B1(n67501), .B2(n66333), .C1(n67495), .C2(n58151), .A(
        n64681), .ZN(n64665) );
  NOR4_X1 U50831 ( .A1(n64677), .A2(n64678), .A3(n64679), .A4(n64680), .ZN(
        n64666) );
  NAND4_X1 U50832 ( .A1(n64644), .A2(n64645), .A3(n64646), .A4(n64647), .ZN(
        n5417) );
  AOI221_X1 U50833 ( .B1(n67477), .B2(n57515), .C1(n67471), .C2(n59050), .A(
        n64662), .ZN(n64644) );
  AOI221_X1 U50834 ( .B1(n67501), .B2(n66334), .C1(n67495), .C2(n58153), .A(
        n64661), .ZN(n64645) );
  NOR4_X1 U50835 ( .A1(n64657), .A2(n64658), .A3(n64659), .A4(n64660), .ZN(
        n64646) );
  NAND4_X1 U50836 ( .A1(n64624), .A2(n64625), .A3(n64626), .A4(n64627), .ZN(
        n5419) );
  AOI221_X1 U50837 ( .B1(n67477), .B2(n57491), .C1(n67471), .C2(n59051), .A(
        n64642), .ZN(n64624) );
  AOI221_X1 U50838 ( .B1(n67501), .B2(n66335), .C1(n67495), .C2(n58155), .A(
        n64641), .ZN(n64625) );
  NOR4_X1 U50839 ( .A1(n64637), .A2(n64638), .A3(n64639), .A4(n64640), .ZN(
        n64626) );
  NAND4_X1 U50840 ( .A1(n64604), .A2(n64605), .A3(n64606), .A4(n64607), .ZN(
        n5421) );
  AOI221_X1 U50841 ( .B1(n67477), .B2(n57467), .C1(n67471), .C2(n59052), .A(
        n64622), .ZN(n64604) );
  AOI221_X1 U50842 ( .B1(n67501), .B2(n66336), .C1(n67495), .C2(n58157), .A(
        n64621), .ZN(n64605) );
  NOR4_X1 U50843 ( .A1(n64617), .A2(n64618), .A3(n64619), .A4(n64620), .ZN(
        n64606) );
  NAND4_X1 U50844 ( .A1(n64584), .A2(n64585), .A3(n64586), .A4(n64587), .ZN(
        n5423) );
  AOI221_X1 U50845 ( .B1(n67478), .B2(n57443), .C1(n67472), .C2(n59053), .A(
        n64602), .ZN(n64584) );
  AOI221_X1 U50846 ( .B1(n67502), .B2(n66337), .C1(n67496), .C2(n58159), .A(
        n64601), .ZN(n64585) );
  NOR4_X1 U50847 ( .A1(n64597), .A2(n64598), .A3(n64599), .A4(n64600), .ZN(
        n64586) );
  NAND4_X1 U50848 ( .A1(n64564), .A2(n64565), .A3(n64566), .A4(n64567), .ZN(
        n5425) );
  AOI221_X1 U50849 ( .B1(n67478), .B2(n57419), .C1(n67472), .C2(n59054), .A(
        n64582), .ZN(n64564) );
  AOI221_X1 U50850 ( .B1(n67502), .B2(n66338), .C1(n67496), .C2(n58161), .A(
        n64581), .ZN(n64565) );
  NOR4_X1 U50851 ( .A1(n64577), .A2(n64578), .A3(n64579), .A4(n64580), .ZN(
        n64566) );
  NAND4_X1 U50852 ( .A1(n64544), .A2(n64545), .A3(n64546), .A4(n64547), .ZN(
        n5427) );
  AOI221_X1 U50853 ( .B1(n67478), .B2(n57395), .C1(n67472), .C2(n59055), .A(
        n64562), .ZN(n64544) );
  AOI221_X1 U50854 ( .B1(n67502), .B2(n66339), .C1(n67496), .C2(n58163), .A(
        n64561), .ZN(n64545) );
  NOR4_X1 U50855 ( .A1(n64557), .A2(n64558), .A3(n64559), .A4(n64560), .ZN(
        n64546) );
  NAND4_X1 U50856 ( .A1(n64524), .A2(n64525), .A3(n64526), .A4(n64527), .ZN(
        n5429) );
  AOI221_X1 U50857 ( .B1(n67478), .B2(n57371), .C1(n67472), .C2(n59056), .A(
        n64542), .ZN(n64524) );
  AOI221_X1 U50858 ( .B1(n67502), .B2(n66340), .C1(n67496), .C2(n58165), .A(
        n64541), .ZN(n64525) );
  NOR4_X1 U50859 ( .A1(n64537), .A2(n64538), .A3(n64539), .A4(n64540), .ZN(
        n64526) );
  NAND4_X1 U50860 ( .A1(n64504), .A2(n64505), .A3(n64506), .A4(n64507), .ZN(
        n5431) );
  AOI221_X1 U50861 ( .B1(n67478), .B2(n57347), .C1(n67472), .C2(n59057), .A(
        n64522), .ZN(n64504) );
  AOI221_X1 U50862 ( .B1(n67502), .B2(n66341), .C1(n67496), .C2(n58167), .A(
        n64521), .ZN(n64505) );
  NOR4_X1 U50863 ( .A1(n64517), .A2(n64518), .A3(n64519), .A4(n64520), .ZN(
        n64506) );
  NAND4_X1 U50864 ( .A1(n64484), .A2(n64485), .A3(n64486), .A4(n64487), .ZN(
        n5433) );
  AOI221_X1 U50865 ( .B1(n67478), .B2(n57323), .C1(n67472), .C2(n59058), .A(
        n64502), .ZN(n64484) );
  AOI221_X1 U50866 ( .B1(n67502), .B2(n66342), .C1(n67496), .C2(n58169), .A(
        n64501), .ZN(n64485) );
  NOR4_X1 U50867 ( .A1(n64497), .A2(n64498), .A3(n64499), .A4(n64500), .ZN(
        n64486) );
  NAND4_X1 U50868 ( .A1(n64464), .A2(n64465), .A3(n64466), .A4(n64467), .ZN(
        n5435) );
  AOI221_X1 U50869 ( .B1(n67478), .B2(n57299), .C1(n67472), .C2(n59059), .A(
        n64482), .ZN(n64464) );
  AOI221_X1 U50870 ( .B1(n67502), .B2(n66343), .C1(n67496), .C2(n58171), .A(
        n64481), .ZN(n64465) );
  NOR4_X1 U50871 ( .A1(n64477), .A2(n64478), .A3(n64479), .A4(n64480), .ZN(
        n64466) );
  NAND4_X1 U50872 ( .A1(n64444), .A2(n64445), .A3(n64446), .A4(n64447), .ZN(
        n5437) );
  AOI221_X1 U50873 ( .B1(n67478), .B2(n57275), .C1(n67472), .C2(n59060), .A(
        n64462), .ZN(n64444) );
  AOI221_X1 U50874 ( .B1(n67502), .B2(n66344), .C1(n67496), .C2(n58173), .A(
        n64461), .ZN(n64445) );
  NOR4_X1 U50875 ( .A1(n64457), .A2(n64458), .A3(n64459), .A4(n64460), .ZN(
        n64446) );
  NAND4_X1 U50876 ( .A1(n64424), .A2(n64425), .A3(n64426), .A4(n64427), .ZN(
        n5439) );
  AOI221_X1 U50877 ( .B1(n67478), .B2(n57251), .C1(n67472), .C2(n59061), .A(
        n64442), .ZN(n64424) );
  AOI221_X1 U50878 ( .B1(n67502), .B2(n66345), .C1(n67496), .C2(n58175), .A(
        n64441), .ZN(n64425) );
  NOR4_X1 U50879 ( .A1(n64437), .A2(n64438), .A3(n64439), .A4(n64440), .ZN(
        n64426) );
  NAND4_X1 U50880 ( .A1(n64404), .A2(n64405), .A3(n64406), .A4(n64407), .ZN(
        n5441) );
  AOI221_X1 U50881 ( .B1(n67478), .B2(n57227), .C1(n67472), .C2(n59062), .A(
        n64422), .ZN(n64404) );
  AOI221_X1 U50882 ( .B1(n67502), .B2(n66346), .C1(n67496), .C2(n58177), .A(
        n64421), .ZN(n64405) );
  NOR4_X1 U50883 ( .A1(n64417), .A2(n64418), .A3(n64419), .A4(n64420), .ZN(
        n64406) );
  NAND4_X1 U50884 ( .A1(n64384), .A2(n64385), .A3(n64386), .A4(n64387), .ZN(
        n5443) );
  AOI221_X1 U50885 ( .B1(n67478), .B2(n57203), .C1(n67472), .C2(n59063), .A(
        n64402), .ZN(n64384) );
  AOI221_X1 U50886 ( .B1(n67502), .B2(n66347), .C1(n67496), .C2(n58179), .A(
        n64401), .ZN(n64385) );
  NOR4_X1 U50887 ( .A1(n64397), .A2(n64398), .A3(n64399), .A4(n64400), .ZN(
        n64386) );
  NAND4_X1 U50888 ( .A1(n64364), .A2(n64365), .A3(n64366), .A4(n64367), .ZN(
        n5445) );
  AOI221_X1 U50889 ( .B1(n67478), .B2(n57179), .C1(n67472), .C2(n59064), .A(
        n64382), .ZN(n64364) );
  AOI221_X1 U50890 ( .B1(n67502), .B2(n66348), .C1(n67496), .C2(n58181), .A(
        n64381), .ZN(n64365) );
  NOR4_X1 U50891 ( .A1(n64377), .A2(n64378), .A3(n64379), .A4(n64380), .ZN(
        n64366) );
  NAND4_X1 U50892 ( .A1(n64344), .A2(n64345), .A3(n64346), .A4(n64347), .ZN(
        n5447) );
  AOI221_X1 U50893 ( .B1(n67479), .B2(n57155), .C1(n67473), .C2(n59065), .A(
        n64362), .ZN(n64344) );
  AOI221_X1 U50894 ( .B1(n67503), .B2(n66349), .C1(n67497), .C2(n58183), .A(
        n64361), .ZN(n64345) );
  NOR4_X1 U50895 ( .A1(n64357), .A2(n64358), .A3(n64359), .A4(n64360), .ZN(
        n64346) );
  NAND4_X1 U50896 ( .A1(n64324), .A2(n64325), .A3(n64326), .A4(n64327), .ZN(
        n5449) );
  AOI221_X1 U50897 ( .B1(n67479), .B2(n57131), .C1(n67473), .C2(n59066), .A(
        n64342), .ZN(n64324) );
  AOI221_X1 U50898 ( .B1(n67503), .B2(n66350), .C1(n67497), .C2(n58185), .A(
        n64341), .ZN(n64325) );
  NOR4_X1 U50899 ( .A1(n64337), .A2(n64338), .A3(n64339), .A4(n64340), .ZN(
        n64326) );
  NAND4_X1 U50900 ( .A1(n64304), .A2(n64305), .A3(n64306), .A4(n64307), .ZN(
        n5451) );
  AOI221_X1 U50901 ( .B1(n67479), .B2(n57107), .C1(n67473), .C2(n59067), .A(
        n64322), .ZN(n64304) );
  AOI221_X1 U50902 ( .B1(n67503), .B2(n66351), .C1(n67497), .C2(n58187), .A(
        n64321), .ZN(n64305) );
  NOR4_X1 U50903 ( .A1(n64317), .A2(n64318), .A3(n64319), .A4(n64320), .ZN(
        n64306) );
  NAND4_X1 U50904 ( .A1(n64284), .A2(n64285), .A3(n64286), .A4(n64287), .ZN(
        n5453) );
  AOI221_X1 U50905 ( .B1(n67479), .B2(n57083), .C1(n67473), .C2(n59068), .A(
        n64302), .ZN(n64284) );
  AOI221_X1 U50906 ( .B1(n67503), .B2(n66352), .C1(n67497), .C2(n58189), .A(
        n64301), .ZN(n64285) );
  NOR4_X1 U50907 ( .A1(n64297), .A2(n64298), .A3(n64299), .A4(n64300), .ZN(
        n64286) );
  NAND4_X1 U50908 ( .A1(n64264), .A2(n64265), .A3(n64266), .A4(n64267), .ZN(
        n5455) );
  AOI221_X1 U50909 ( .B1(n67479), .B2(n57059), .C1(n67473), .C2(n59069), .A(
        n64282), .ZN(n64264) );
  AOI221_X1 U50910 ( .B1(n67503), .B2(n66353), .C1(n67497), .C2(n58191), .A(
        n64281), .ZN(n64265) );
  NOR4_X1 U50911 ( .A1(n64277), .A2(n64278), .A3(n64279), .A4(n64280), .ZN(
        n64266) );
  NAND4_X1 U50912 ( .A1(n64244), .A2(n64245), .A3(n64246), .A4(n64247), .ZN(
        n5457) );
  AOI221_X1 U50913 ( .B1(n67479), .B2(n57035), .C1(n67473), .C2(n59070), .A(
        n64262), .ZN(n64244) );
  AOI221_X1 U50914 ( .B1(n67503), .B2(n66354), .C1(n67497), .C2(n58193), .A(
        n64261), .ZN(n64245) );
  NOR4_X1 U50915 ( .A1(n64257), .A2(n64258), .A3(n64259), .A4(n64260), .ZN(
        n64246) );
  NAND4_X1 U50916 ( .A1(n64224), .A2(n64225), .A3(n64226), .A4(n64227), .ZN(
        n5459) );
  AOI221_X1 U50917 ( .B1(n67479), .B2(n57011), .C1(n67473), .C2(n59071), .A(
        n64242), .ZN(n64224) );
  AOI221_X1 U50918 ( .B1(n67503), .B2(n66355), .C1(n67497), .C2(n58195), .A(
        n64241), .ZN(n64225) );
  NOR4_X1 U50919 ( .A1(n64237), .A2(n64238), .A3(n64239), .A4(n64240), .ZN(
        n64226) );
  NAND4_X1 U50920 ( .A1(n64204), .A2(n64205), .A3(n64206), .A4(n64207), .ZN(
        n5461) );
  AOI221_X1 U50921 ( .B1(n67479), .B2(n56987), .C1(n67473), .C2(n59072), .A(
        n64222), .ZN(n64204) );
  AOI221_X1 U50922 ( .B1(n67503), .B2(n66356), .C1(n67497), .C2(n58197), .A(
        n64221), .ZN(n64205) );
  NOR4_X1 U50923 ( .A1(n64217), .A2(n64218), .A3(n64219), .A4(n64220), .ZN(
        n64206) );
  NAND4_X1 U50924 ( .A1(n64184), .A2(n64185), .A3(n64186), .A4(n64187), .ZN(
        n5463) );
  AOI221_X1 U50925 ( .B1(n67479), .B2(n56963), .C1(n67473), .C2(n59073), .A(
        n64202), .ZN(n64184) );
  AOI221_X1 U50926 ( .B1(n67503), .B2(n66357), .C1(n67497), .C2(n58199), .A(
        n64201), .ZN(n64185) );
  NOR4_X1 U50927 ( .A1(n64197), .A2(n64198), .A3(n64199), .A4(n64200), .ZN(
        n64186) );
  NAND4_X1 U50928 ( .A1(n64164), .A2(n64165), .A3(n64166), .A4(n64167), .ZN(
        n5465) );
  AOI221_X1 U50929 ( .B1(n67479), .B2(n56939), .C1(n67473), .C2(n59074), .A(
        n64182), .ZN(n64164) );
  AOI221_X1 U50930 ( .B1(n67503), .B2(n66358), .C1(n67497), .C2(n58201), .A(
        n64181), .ZN(n64165) );
  NOR4_X1 U50931 ( .A1(n64177), .A2(n64178), .A3(n64179), .A4(n64180), .ZN(
        n64166) );
  NAND4_X1 U50932 ( .A1(n64144), .A2(n64145), .A3(n64146), .A4(n64147), .ZN(
        n5467) );
  AOI221_X1 U50933 ( .B1(n67479), .B2(n56915), .C1(n67473), .C2(n59075), .A(
        n64162), .ZN(n64144) );
  AOI221_X1 U50934 ( .B1(n67503), .B2(n66359), .C1(n67497), .C2(n58203), .A(
        n64161), .ZN(n64145) );
  NOR4_X1 U50935 ( .A1(n64157), .A2(n64158), .A3(n64159), .A4(n64160), .ZN(
        n64146) );
  NAND4_X1 U50936 ( .A1(n64124), .A2(n64125), .A3(n64126), .A4(n64127), .ZN(
        n5469) );
  AOI221_X1 U50937 ( .B1(n67479), .B2(n56891), .C1(n67473), .C2(n59076), .A(
        n64142), .ZN(n64124) );
  AOI221_X1 U50938 ( .B1(n67503), .B2(n66360), .C1(n67497), .C2(n58205), .A(
        n64141), .ZN(n64125) );
  NOR4_X1 U50939 ( .A1(n64137), .A2(n64138), .A3(n64139), .A4(n64140), .ZN(
        n64126) );
  NAND4_X1 U50940 ( .A1(n64104), .A2(n64105), .A3(n64106), .A4(n64107), .ZN(
        n5471) );
  AOI221_X1 U50941 ( .B1(n67480), .B2(n56867), .C1(n67474), .C2(n59077), .A(
        n64122), .ZN(n64104) );
  AOI221_X1 U50942 ( .B1(n67504), .B2(n66361), .C1(n67498), .C2(n58207), .A(
        n64121), .ZN(n64105) );
  NOR4_X1 U50943 ( .A1(n64117), .A2(n64118), .A3(n64119), .A4(n64120), .ZN(
        n64106) );
  NAND4_X1 U50944 ( .A1(n64084), .A2(n64085), .A3(n64086), .A4(n64087), .ZN(
        n5473) );
  AOI221_X1 U50945 ( .B1(n67480), .B2(n56843), .C1(n67474), .C2(n59078), .A(
        n64102), .ZN(n64084) );
  AOI221_X1 U50946 ( .B1(n67504), .B2(n66362), .C1(n67498), .C2(n58209), .A(
        n64101), .ZN(n64085) );
  NOR4_X1 U50947 ( .A1(n64097), .A2(n64098), .A3(n64099), .A4(n64100), .ZN(
        n64086) );
  NAND4_X1 U50948 ( .A1(n64064), .A2(n64065), .A3(n64066), .A4(n64067), .ZN(
        n5475) );
  AOI221_X1 U50949 ( .B1(n67480), .B2(n56819), .C1(n67474), .C2(n59079), .A(
        n64082), .ZN(n64064) );
  AOI221_X1 U50950 ( .B1(n67504), .B2(n66363), .C1(n67498), .C2(n58211), .A(
        n64081), .ZN(n64065) );
  NOR4_X1 U50951 ( .A1(n64077), .A2(n64078), .A3(n64079), .A4(n64080), .ZN(
        n64066) );
  NAND4_X1 U50952 ( .A1(n64044), .A2(n64045), .A3(n64046), .A4(n64047), .ZN(
        n5477) );
  AOI221_X1 U50953 ( .B1(n67480), .B2(n56795), .C1(n67474), .C2(n59080), .A(
        n64062), .ZN(n64044) );
  AOI221_X1 U50954 ( .B1(n67504), .B2(n66364), .C1(n67498), .C2(n58213), .A(
        n64061), .ZN(n64045) );
  NOR4_X1 U50955 ( .A1(n64057), .A2(n64058), .A3(n64059), .A4(n64060), .ZN(
        n64046) );
  NAND4_X1 U50956 ( .A1(n64024), .A2(n64025), .A3(n64026), .A4(n64027), .ZN(
        n5479) );
  AOI221_X1 U50957 ( .B1(n67480), .B2(n56771), .C1(n67474), .C2(n59081), .A(
        n64042), .ZN(n64024) );
  AOI221_X1 U50958 ( .B1(n67504), .B2(n66365), .C1(n67498), .C2(n58215), .A(
        n64041), .ZN(n64025) );
  NOR4_X1 U50959 ( .A1(n64037), .A2(n64038), .A3(n64039), .A4(n64040), .ZN(
        n64026) );
  NAND4_X1 U50960 ( .A1(n64004), .A2(n64005), .A3(n64006), .A4(n64007), .ZN(
        n5481) );
  AOI221_X1 U50961 ( .B1(n67480), .B2(n56747), .C1(n67474), .C2(n59082), .A(
        n64022), .ZN(n64004) );
  AOI221_X1 U50962 ( .B1(n67504), .B2(n66366), .C1(n67498), .C2(n58217), .A(
        n64021), .ZN(n64005) );
  NOR4_X1 U50963 ( .A1(n64017), .A2(n64018), .A3(n64019), .A4(n64020), .ZN(
        n64006) );
  NAND4_X1 U50964 ( .A1(n63984), .A2(n63985), .A3(n63986), .A4(n63987), .ZN(
        n5483) );
  AOI221_X1 U50965 ( .B1(n67480), .B2(n56723), .C1(n67474), .C2(n59083), .A(
        n64002), .ZN(n63984) );
  AOI221_X1 U50966 ( .B1(n67504), .B2(n66367), .C1(n67498), .C2(n58219), .A(
        n64001), .ZN(n63985) );
  NOR4_X1 U50967 ( .A1(n63997), .A2(n63998), .A3(n63999), .A4(n64000), .ZN(
        n63986) );
  NAND4_X1 U50968 ( .A1(n63964), .A2(n63965), .A3(n63966), .A4(n63967), .ZN(
        n5485) );
  AOI221_X1 U50969 ( .B1(n67480), .B2(n56699), .C1(n67474), .C2(n59084), .A(
        n63982), .ZN(n63964) );
  AOI221_X1 U50970 ( .B1(n67504), .B2(n66368), .C1(n67498), .C2(n58221), .A(
        n63981), .ZN(n63965) );
  NOR4_X1 U50971 ( .A1(n63977), .A2(n63978), .A3(n63979), .A4(n63980), .ZN(
        n63966) );
  NAND4_X1 U50972 ( .A1(n63944), .A2(n63945), .A3(n63946), .A4(n63947), .ZN(
        n5487) );
  AOI221_X1 U50973 ( .B1(n67480), .B2(n56675), .C1(n67474), .C2(n59085), .A(
        n63962), .ZN(n63944) );
  AOI221_X1 U50974 ( .B1(n67504), .B2(n66369), .C1(n67498), .C2(n58223), .A(
        n63961), .ZN(n63945) );
  NOR4_X1 U50975 ( .A1(n63957), .A2(n63958), .A3(n63959), .A4(n63960), .ZN(
        n63946) );
  NAND4_X1 U50976 ( .A1(n63924), .A2(n63925), .A3(n63926), .A4(n63927), .ZN(
        n5489) );
  AOI221_X1 U50977 ( .B1(n67480), .B2(n56651), .C1(n67474), .C2(n59086), .A(
        n63942), .ZN(n63924) );
  AOI221_X1 U50978 ( .B1(n67504), .B2(n66370), .C1(n67498), .C2(n58225), .A(
        n63941), .ZN(n63925) );
  NOR4_X1 U50979 ( .A1(n63937), .A2(n63938), .A3(n63939), .A4(n63940), .ZN(
        n63926) );
  NAND4_X1 U50980 ( .A1(n63904), .A2(n63905), .A3(n63906), .A4(n63907), .ZN(
        n5491) );
  AOI221_X1 U50981 ( .B1(n67480), .B2(n56627), .C1(n67474), .C2(n59087), .A(
        n63922), .ZN(n63904) );
  AOI221_X1 U50982 ( .B1(n67504), .B2(n66371), .C1(n67498), .C2(n58227), .A(
        n63921), .ZN(n63905) );
  NOR4_X1 U50983 ( .A1(n63917), .A2(n63918), .A3(n63919), .A4(n63920), .ZN(
        n63906) );
  NAND4_X1 U50984 ( .A1(n63884), .A2(n63885), .A3(n63886), .A4(n63887), .ZN(
        n5493) );
  AOI221_X1 U50985 ( .B1(n67480), .B2(n56603), .C1(n67474), .C2(n59088), .A(
        n63902), .ZN(n63884) );
  AOI221_X1 U50986 ( .B1(n67504), .B2(n66372), .C1(n67498), .C2(n58229), .A(
        n63901), .ZN(n63885) );
  NOR4_X1 U50987 ( .A1(n63897), .A2(n63898), .A3(n63899), .A4(n63900), .ZN(
        n63886) );
  NAND4_X1 U50988 ( .A1(n63863), .A2(n63864), .A3(n63865), .A4(n63866), .ZN(
        n5495) );
  AOI221_X1 U50989 ( .B1(n67481), .B2(n56579), .C1(n67475), .C2(n59089), .A(
        n63882), .ZN(n63863) );
  AOI221_X1 U50990 ( .B1(n67505), .B2(n66305), .C1(n67499), .C2(n58231), .A(
        n63881), .ZN(n63864) );
  NOR4_X1 U50991 ( .A1(n63867), .A2(n63868), .A3(n63869), .A4(n63870), .ZN(
        n63866) );
  NAND4_X1 U50992 ( .A1(n63842), .A2(n63843), .A3(n63844), .A4(n63845), .ZN(
        n5497) );
  AOI221_X1 U50993 ( .B1(n67481), .B2(n56555), .C1(n67475), .C2(n59090), .A(
        n63861), .ZN(n63842) );
  AOI221_X1 U50994 ( .B1(n67505), .B2(n66306), .C1(n67499), .C2(n58232), .A(
        n63860), .ZN(n63843) );
  NOR4_X1 U50995 ( .A1(n63846), .A2(n63847), .A3(n63848), .A4(n63849), .ZN(
        n63845) );
  NAND4_X1 U50996 ( .A1(n63821), .A2(n63822), .A3(n63823), .A4(n63824), .ZN(
        n5499) );
  AOI221_X1 U50997 ( .B1(n67481), .B2(n56531), .C1(n67475), .C2(n59091), .A(
        n63840), .ZN(n63821) );
  AOI221_X1 U50998 ( .B1(n67505), .B2(n66307), .C1(n67499), .C2(n58233), .A(
        n63839), .ZN(n63822) );
  NOR4_X1 U50999 ( .A1(n63825), .A2(n63826), .A3(n63827), .A4(n63828), .ZN(
        n63824) );
  NAND4_X1 U51000 ( .A1(n63767), .A2(n63768), .A3(n63769), .A4(n63770), .ZN(
        n5501) );
  AOI221_X1 U51001 ( .B1(n67481), .B2(n56490), .C1(n67475), .C2(n59092), .A(
        n63817), .ZN(n63767) );
  AOI221_X1 U51002 ( .B1(n67505), .B2(n66308), .C1(n67499), .C2(n58234), .A(
        n63812), .ZN(n63768) );
  NOR4_X1 U51003 ( .A1(n63771), .A2(n63772), .A3(n63773), .A4(n63774), .ZN(
        n63770) );
  AND3_X1 U51004 ( .A1(WR), .A2(ENABLE), .A3(ADD_WR[4]), .ZN(n63295) );
  INV_X1 U51005 ( .A(RESET), .ZN(n62087) );
  INV_X1 U51006 ( .A(DATAIN[60]), .ZN(n61966) );
  INV_X1 U51007 ( .A(DATAIN[61]), .ZN(n61964) );
  INV_X1 U51008 ( .A(DATAIN[62]), .ZN(n61962) );
  INV_X1 U51009 ( .A(DATAIN[63]), .ZN(n61960) );
  INV_X1 U51010 ( .A(DATAIN[0]), .ZN(n62086) );
  INV_X1 U51011 ( .A(DATAIN[1]), .ZN(n62084) );
  INV_X1 U51012 ( .A(DATAIN[2]), .ZN(n62082) );
  INV_X1 U51013 ( .A(DATAIN[3]), .ZN(n62080) );
  INV_X1 U51014 ( .A(DATAIN[4]), .ZN(n62078) );
  INV_X1 U51015 ( .A(DATAIN[5]), .ZN(n62076) );
  INV_X1 U51016 ( .A(DATAIN[6]), .ZN(n62074) );
  INV_X1 U51017 ( .A(DATAIN[7]), .ZN(n62072) );
  INV_X1 U51018 ( .A(DATAIN[8]), .ZN(n62070) );
  INV_X1 U51019 ( .A(DATAIN[9]), .ZN(n62068) );
  INV_X1 U51020 ( .A(DATAIN[10]), .ZN(n62066) );
  INV_X1 U51021 ( .A(DATAIN[11]), .ZN(n62064) );
  INV_X1 U51022 ( .A(DATAIN[12]), .ZN(n62062) );
  INV_X1 U51023 ( .A(DATAIN[13]), .ZN(n62060) );
  INV_X1 U51024 ( .A(DATAIN[14]), .ZN(n62058) );
  INV_X1 U51025 ( .A(DATAIN[15]), .ZN(n62056) );
  INV_X1 U51026 ( .A(DATAIN[16]), .ZN(n62054) );
  INV_X1 U51027 ( .A(DATAIN[17]), .ZN(n62052) );
  INV_X1 U51028 ( .A(DATAIN[18]), .ZN(n62050) );
  INV_X1 U51029 ( .A(DATAIN[19]), .ZN(n62048) );
  INV_X1 U51030 ( .A(DATAIN[20]), .ZN(n62046) );
  INV_X1 U51031 ( .A(DATAIN[21]), .ZN(n62044) );
  INV_X1 U51032 ( .A(DATAIN[22]), .ZN(n62042) );
  INV_X1 U51033 ( .A(DATAIN[23]), .ZN(n62040) );
  INV_X1 U51034 ( .A(DATAIN[24]), .ZN(n62038) );
  INV_X1 U51035 ( .A(DATAIN[25]), .ZN(n62036) );
  INV_X1 U51036 ( .A(DATAIN[26]), .ZN(n62034) );
  INV_X1 U51037 ( .A(DATAIN[27]), .ZN(n62032) );
  INV_X1 U51038 ( .A(DATAIN[28]), .ZN(n62030) );
  INV_X1 U51039 ( .A(DATAIN[29]), .ZN(n62028) );
  INV_X1 U51040 ( .A(DATAIN[30]), .ZN(n62026) );
  INV_X1 U51041 ( .A(DATAIN[31]), .ZN(n62024) );
  INV_X1 U51042 ( .A(DATAIN[32]), .ZN(n62022) );
  INV_X1 U51043 ( .A(DATAIN[33]), .ZN(n62020) );
  INV_X1 U51044 ( .A(DATAIN[34]), .ZN(n62018) );
  INV_X1 U51045 ( .A(DATAIN[35]), .ZN(n62016) );
  INV_X1 U51046 ( .A(DATAIN[36]), .ZN(n62014) );
  INV_X1 U51047 ( .A(DATAIN[37]), .ZN(n62012) );
  INV_X1 U51048 ( .A(DATAIN[38]), .ZN(n62010) );
  INV_X1 U51049 ( .A(DATAIN[39]), .ZN(n62008) );
  INV_X1 U51050 ( .A(DATAIN[40]), .ZN(n62006) );
  INV_X1 U51051 ( .A(DATAIN[41]), .ZN(n62004) );
  INV_X1 U51052 ( .A(DATAIN[42]), .ZN(n62002) );
  INV_X1 U51053 ( .A(DATAIN[43]), .ZN(n62000) );
  INV_X1 U51054 ( .A(DATAIN[44]), .ZN(n61998) );
  INV_X1 U51055 ( .A(DATAIN[45]), .ZN(n61996) );
  INV_X1 U51056 ( .A(DATAIN[46]), .ZN(n61994) );
  INV_X1 U51057 ( .A(DATAIN[47]), .ZN(n61992) );
  INV_X1 U51058 ( .A(DATAIN[48]), .ZN(n61990) );
  INV_X1 U51059 ( .A(DATAIN[49]), .ZN(n61988) );
  INV_X1 U51060 ( .A(DATAIN[50]), .ZN(n61986) );
  INV_X1 U51061 ( .A(DATAIN[51]), .ZN(n61984) );
  INV_X1 U51062 ( .A(DATAIN[52]), .ZN(n61982) );
  INV_X1 U51063 ( .A(DATAIN[53]), .ZN(n61980) );
  INV_X1 U51064 ( .A(DATAIN[54]), .ZN(n61978) );
  INV_X1 U51065 ( .A(DATAIN[55]), .ZN(n61976) );
  INV_X1 U51066 ( .A(DATAIN[56]), .ZN(n61974) );
  INV_X1 U51067 ( .A(DATAIN[57]), .ZN(n61972) );
  INV_X1 U51068 ( .A(DATAIN[58]), .ZN(n61970) );
  INV_X1 U51069 ( .A(DATAIN[59]), .ZN(n61968) );
  INV_X1 U51070 ( .A(ADD_WR[3]), .ZN(n62491) );
  INV_X1 U51071 ( .A(ADD_WR[0]), .ZN(n62490) );
  INV_X1 U51072 ( .A(ADD_WR[1]), .ZN(n63497) );
  INV_X1 U51073 ( .A(ADD_RD2[2]), .ZN(n66299) );
  INV_X1 U51074 ( .A(ADD_RD2[1]), .ZN(n66301) );
  INV_X1 U51075 ( .A(ADD_WR[2]), .ZN(n63496) );
  INV_X1 U51076 ( .A(ADD_RD1[2]), .ZN(n65099) );
  AND3_X1 U51077 ( .A1(ENABLE), .A2(n62958), .A3(WR), .ZN(n62492) );
  INV_X1 U51078 ( .A(ADD_WR[4]), .ZN(n62958) );
  CLKBUF_X1 U51079 ( .A(n65150), .Z(n67265) );
  CLKBUF_X1 U51080 ( .A(n65149), .Z(n67271) );
  CLKBUF_X1 U51081 ( .A(n65147), .Z(n67277) );
  CLKBUF_X1 U51082 ( .A(n65146), .Z(n67283) );
  CLKBUF_X1 U51083 ( .A(n65145), .Z(n67289) );
  CLKBUF_X1 U51084 ( .A(n65144), .Z(n67295) );
  CLKBUF_X1 U51085 ( .A(n65142), .Z(n67301) );
  CLKBUF_X1 U51086 ( .A(n65141), .Z(n67307) );
  CLKBUF_X1 U51087 ( .A(n65140), .Z(n67313) );
  CLKBUF_X1 U51088 ( .A(n65139), .Z(n67319) );
  CLKBUF_X1 U51089 ( .A(n65138), .Z(n67325) );
  CLKBUF_X1 U51090 ( .A(n65137), .Z(n67331) );
  CLKBUF_X1 U51091 ( .A(n65136), .Z(n67337) );
  CLKBUF_X1 U51092 ( .A(n65135), .Z(n67343) );
  CLKBUF_X1 U51093 ( .A(n65134), .Z(n67349) );
  CLKBUF_X1 U51094 ( .A(n65133), .Z(n67355) );
  CLKBUF_X1 U51095 ( .A(n65132), .Z(n67361) );
  CLKBUF_X1 U51096 ( .A(n65127), .Z(n67367) );
  CLKBUF_X1 U51097 ( .A(n65126), .Z(n67373) );
  CLKBUF_X1 U51098 ( .A(n65124), .Z(n67379) );
  CLKBUF_X1 U51099 ( .A(n65123), .Z(n67385) );
  CLKBUF_X1 U51100 ( .A(n65122), .Z(n67391) );
  CLKBUF_X1 U51101 ( .A(n65121), .Z(n67397) );
  CLKBUF_X1 U51102 ( .A(n65119), .Z(n67403) );
  CLKBUF_X1 U51103 ( .A(n65118), .Z(n67409) );
  CLKBUF_X1 U51104 ( .A(n65117), .Z(n67415) );
  CLKBUF_X1 U51105 ( .A(n65116), .Z(n67421) );
  CLKBUF_X1 U51106 ( .A(n65114), .Z(n67427) );
  CLKBUF_X1 U51107 ( .A(n65113), .Z(n67433) );
  CLKBUF_X1 U51108 ( .A(n65112), .Z(n67439) );
  CLKBUF_X1 U51109 ( .A(n65111), .Z(n67445) );
  CLKBUF_X1 U51110 ( .A(n65109), .Z(n67451) );
  CLKBUF_X1 U51111 ( .A(n65108), .Z(n67457) );
  CLKBUF_X1 U51112 ( .A(n63819), .Z(n67463) );
  CLKBUF_X1 U51113 ( .A(n63818), .Z(n67469) );
  CLKBUF_X1 U51114 ( .A(n63816), .Z(n67475) );
  CLKBUF_X1 U51115 ( .A(n63815), .Z(n67481) );
  CLKBUF_X1 U51116 ( .A(n63814), .Z(n67487) );
  CLKBUF_X1 U51117 ( .A(n63813), .Z(n67493) );
  CLKBUF_X1 U51118 ( .A(n63811), .Z(n67499) );
  CLKBUF_X1 U51119 ( .A(n63810), .Z(n67505) );
  CLKBUF_X1 U51120 ( .A(n63809), .Z(n67511) );
  CLKBUF_X1 U51121 ( .A(n63808), .Z(n67517) );
  CLKBUF_X1 U51122 ( .A(n63807), .Z(n67523) );
  CLKBUF_X1 U51123 ( .A(n63806), .Z(n67529) );
  CLKBUF_X1 U51124 ( .A(n63805), .Z(n67535) );
  CLKBUF_X1 U51125 ( .A(n63804), .Z(n67541) );
  CLKBUF_X1 U51126 ( .A(n63803), .Z(n67547) );
  CLKBUF_X1 U51127 ( .A(n63802), .Z(n67553) );
  CLKBUF_X1 U51128 ( .A(n63801), .Z(n67559) );
  CLKBUF_X1 U51129 ( .A(n63795), .Z(n67565) );
  CLKBUF_X1 U51130 ( .A(n63794), .Z(n67571) );
  CLKBUF_X1 U51131 ( .A(n63792), .Z(n67577) );
  CLKBUF_X1 U51132 ( .A(n63791), .Z(n67583) );
  CLKBUF_X1 U51133 ( .A(n63790), .Z(n67589) );
  CLKBUF_X1 U51134 ( .A(n63788), .Z(n67595) );
  CLKBUF_X1 U51135 ( .A(n63786), .Z(n67601) );
  CLKBUF_X1 U51136 ( .A(n63785), .Z(n67607) );
  CLKBUF_X1 U51137 ( .A(n63784), .Z(n67613) );
  CLKBUF_X1 U51138 ( .A(n63783), .Z(n67619) );
  CLKBUF_X1 U51139 ( .A(n63781), .Z(n67625) );
  CLKBUF_X1 U51140 ( .A(n63780), .Z(n67631) );
  CLKBUF_X1 U51141 ( .A(n63778), .Z(n67641) );
  CLKBUF_X1 U51142 ( .A(n63776), .Z(n67647) );
  CLKBUF_X1 U51143 ( .A(n63775), .Z(n67653) );
  CLKBUF_X1 U51144 ( .A(n63766), .Z(n67659) );
  CLKBUF_X1 U51145 ( .A(n63700), .Z(n67672) );
  CLKBUF_X1 U51146 ( .A(n63634), .Z(n67685) );
  CLKBUF_X1 U51147 ( .A(n63568), .Z(n67698) );
  CLKBUF_X1 U51148 ( .A(n63502), .Z(n67711) );
  CLKBUF_X1 U51149 ( .A(n63499), .Z(n67724) );
  CLKBUF_X1 U51150 ( .A(n63498), .Z(n67730) );
  CLKBUF_X1 U51151 ( .A(n63431), .Z(n67736) );
  CLKBUF_X1 U51152 ( .A(n63364), .Z(n67749) );
  CLKBUF_X1 U51153 ( .A(n63298), .Z(n67762) );
  CLKBUF_X1 U51154 ( .A(n63231), .Z(n67775) );
  CLKBUF_X1 U51155 ( .A(n63228), .Z(n67788) );
  CLKBUF_X1 U51156 ( .A(n63227), .Z(n67794) );
  CLKBUF_X1 U51157 ( .A(n63163), .Z(n67800) );
  CLKBUF_X1 U51158 ( .A(n63097), .Z(n67813) );
  CLKBUF_X1 U51159 ( .A(n63094), .Z(n67826) );
  CLKBUF_X1 U51160 ( .A(n63093), .Z(n67832) );
  CLKBUF_X1 U51161 ( .A(n63028), .Z(n67838) );
  CLKBUF_X1 U51162 ( .A(n62961), .Z(n67851) );
  CLKBUF_X1 U51163 ( .A(n62894), .Z(n67864) );
  CLKBUF_X1 U51164 ( .A(n62828), .Z(n67877) );
  CLKBUF_X1 U51165 ( .A(n62765), .Z(n67890) );
  CLKBUF_X1 U51166 ( .A(n62763), .Z(n67903) );
  CLKBUF_X1 U51167 ( .A(n62762), .Z(n67909) );
  CLKBUF_X1 U51168 ( .A(n62698), .Z(n67915) );
  CLKBUF_X1 U51169 ( .A(n62695), .Z(n67928) );
  CLKBUF_X1 U51170 ( .A(n62693), .Z(n67934) );
  CLKBUF_X1 U51171 ( .A(n62628), .Z(n67940) );
  CLKBUF_X1 U51172 ( .A(n62561), .Z(n67953) );
  CLKBUF_X1 U51173 ( .A(n62495), .Z(n67966) );
  CLKBUF_X1 U51174 ( .A(n62425), .Z(n67979) );
  CLKBUF_X1 U51175 ( .A(n62359), .Z(n67992) );
  CLKBUF_X1 U51176 ( .A(n62292), .Z(n68005) );
  CLKBUF_X1 U51177 ( .A(n62226), .Z(n68018) );
  CLKBUF_X1 U51178 ( .A(n62159), .Z(n68031) );
  CLKBUF_X1 U51179 ( .A(n62092), .Z(n68044) );
  CLKBUF_X1 U51180 ( .A(n62087), .Z(n68057) );
  CLKBUF_X1 U51181 ( .A(n61959), .Z(n68255) );
endmodule

