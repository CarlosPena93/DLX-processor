package CONSTANTS is
   constant IVDELAY : time := 0 ns;--0.1 ns;
   constant NDDELAY : time := 0 ns;--0.2 ns;
   constant NDDELAYRISE : time := 0 ns;--0.6 ns;
   constant NDDELAYFALL : time := 0 ns;--0.4 ns;
   constant NRDELAY : time := 0 ns;--0.2 ns;
   constant DRCAS : time := 0 ns;--1 ns;
   constant DRCAC : time := 0 ns;--2 ns;
   constant NumBit : integer := 32;	
   constant N_bit : integer := 4;
   constant CBIT : integer := 8; --division between Numbit and Cbit
   constant TP_MUX : time := 0 ns;--0 ns;	
end CONSTANTS;


package body CONSTANTS is

  function log2 ( arg: integer )  return integer is
    variable temp    : integer := arg;
    variable result : integer := 0;
  begin
    while temp > 1 loop
      result := result + 1;
      temp    := temp / 2;
    end loop;
    return result;
  end function log2 ;

end CONSTANTS;
