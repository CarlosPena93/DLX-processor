
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_registerfile_generic_n_bit32_data_bit64 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_registerfile_generic_n_bit32_data_bit64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerfile_generic_n_bit32_data_bit64.all;

entity registerfile_generic_n_bit32_data_bit64 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (5 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end registerfile_generic_n_bit32_data_bit64;

architecture SYN_A of registerfile_generic_n_bit32_data_bit64 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, OUT1_59_port,
      OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, OUT1_54_port, 
      OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, OUT1_49_port, 
      OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, OUT1_44_port, 
      OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, OUT1_39_port, 
      OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, OUT1_34_port, 
      OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, OUT1_29_port, 
      OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, 
      OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, 
      OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, 
      OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, 
      OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, 
      OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, OUT2_63_port, 
      OUT2_62_port, OUT2_61_port, OUT2_60_port, OUT2_59_port, OUT2_58_port, 
      OUT2_57_port, OUT2_56_port, OUT2_55_port, OUT2_54_port, OUT2_53_port, 
      OUT2_52_port, OUT2_51_port, OUT2_50_port, OUT2_49_port, OUT2_48_port, 
      OUT2_47_port, OUT2_46_port, OUT2_45_port, OUT2_44_port, OUT2_43_port, 
      OUT2_42_port, OUT2_41_port, OUT2_40_port, OUT2_39_port, OUT2_38_port, 
      OUT2_37_port, OUT2_36_port, OUT2_35_port, OUT2_34_port, OUT2_33_port, 
      OUT2_32_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port, n4159, n4160, n4161, n4162, n4163,
      n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
      n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, 
      n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, 
      n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, 
      n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4223, n4224, n4225, 
      n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, 
      n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, 
      n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, 
      n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, 
      n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, 
      n4276, n4277, n4278, n4279, n4280, n4281, n4282, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, 
      n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, 
      n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, 
      n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, 
      n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, 
      n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, 
      n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, 
      n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, 
      n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, 
      n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, 
      n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, 
      n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, 
      n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, 
      n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, 
      n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
      n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, 
      n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, 
      n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, 
      n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, 
      n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, 
      n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, 
      n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, 
      n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, 
      n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, 
      n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, 
      n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, 
      n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
      n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, 
      n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, 
      n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, 
      n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, 
      n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, 
      n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, 
      n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, 
      n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, 
      n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, 
      n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, 
      n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, 
      n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, 
      n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, 
      n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, 
      n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, 
      n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, 
      n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, 
      n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, 
      n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, 
      n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, 
      n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, 
      n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, 
      n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, 
      n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, 
      n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, 
      n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, 
      n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, 
      n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, 
      n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, 
      n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, 
      n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
      n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, 
      n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, 
      n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, 
      n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, 
      n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
      n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, 
      n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, 
      n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, 
      n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, 
      n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, 
      n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, 
      n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, 
      n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, 
      n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, 
      n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, 
      n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, 
      n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, 
      n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, 
      n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, 
      n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, 
      n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, 
      n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, 
      n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, 
      n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, 
      n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, 
      n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, 
      n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, 
      n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, 
      n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, 
      n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, 
      n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, 
      n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
      n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, 
      n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, 
      n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, 
      n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
      n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, 
      n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, 
      n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, 
      n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, 
      n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, 
      n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, 
      n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
      n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, 
      n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
      n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, 
      n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, 
      n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, 
      n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, 
      n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, 
      n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, 
      n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
      n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, 
      n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
      n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
      n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
      n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, 
      n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, 
      n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
      n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, 
      n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, 
      n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, 
      n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
      n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, 
      n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, 
      n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
      n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, 
      n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
      n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, 
      n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
      n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, 
      n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7489, n7505, n7521, n7537, n7553, n7569, n7585, 
      n7601, n7617, n7633, n7649, n7665, n7681, n7697, n7713, n7729, n7745, 
      n7761, n7777, n7793, n7809, n7825, n7841, n7857, n7873, n7889, n7905, 
      n7921, n7937, n7953, n7969, n7985, n8001, n8017, n8033, n8049, n8065, 
      n8081, n8097, n8113, n8129, n8145, n8161, n8177, n8193, n8209, n8225, 
      n8241, n8257, n8273, n8289, n8305, n8321, n8337, n8353, n8369, n8385, 
      n8401, n8417, n8433, n8449, n8461, n8465, n8477, n8481, n8493, n8497, 
      n8509, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, 
      n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, 
      n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
      n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, 
      n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8956, n8957, n8958, n8959, n8961, n8963, n8965, n8967, 
      n8969, n8971, n8973, n8975, n8977, n8979, n8981, n8983, n8985, n8987, 
      n8989, n8991, n8993, n8995, n8997, n8999, n9001, n9003, n9005, n9007, 
      n9009, n9011, n9013, n9015, n9017, n9019, n9021, n9023, n9025, n9027, 
      n9029, n9031, n9033, n9035, n9037, n9039, n9041, n9043, n9045, n9047, 
      n9049, n9051, n9053, n9055, n9057, n9059, n9061, n9063, n9065, n9067, 
      n9069, n9071, n9073, n9075, n9077, n9079, n9081, n9083, n9085, n41759, 
      n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768, 
      n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777, 
      n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786, 
      n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795, 
      n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804, 
      n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41813, 
      n41814, n41815, n41816, n41817, n41818, n42003, n42004, n42005, n42006, 
      n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235, n49236, 
      n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244, n49245, 
      n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254, 
      n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262, n49263, 
      n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272, 
      n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280, n49281, 
      n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290, 
      n49291, n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427, 
      n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436, 
      n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445, 
      n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454, 
      n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463, 
      n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472, 
      n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481, 
      n49482, n49483, n50517, n50518, n50519, n50520, n50521, n50522, n50523, 
      n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532, 
      n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540, n50541, 
      n50542, n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550, 
      n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558, n50559, 
      n50560, n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568, 
      n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576, n50577, 
      n50578, n50579, n50644, n50645, n50646, n50647, n50648, n50649, n50650, 
      n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659, 
      n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668, 
      n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676, n50677, 
      n50678, n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686, 
      n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695, 
      n50696, n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704, 
      n50705, n50706, n50707, n54184, n54185, n54186, n54187, n54188, n54189, 
      n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, 
      n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, 
      n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, 
      n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, 
      n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, 
      n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, 
      n54244, n54245, n54246, n54606, n54608, n54609, n54610, n54611, n54612, 
      n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, 
      n54622, n54623, n54624, n54625, n54626, n54627, n54628, n54629, n54630, 
      n54631, n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639, 
      n54640, n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648, 
      n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657, 
      n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666, 
      n54667, n54668, n54669, n54670, n56020, n56047, n56074, n56101, n56490, 
      n56531, n56555, n56579, n56597, n56603, n56609, n56611, n56621, n56627, 
      n56633, n56635, n56645, n56651, n56657, n56659, n56669, n56675, n56681, 
      n56683, n56693, n56699, n56705, n56707, n56717, n56723, n56729, n56731, 
      n56741, n56747, n56753, n56755, n56765, n56771, n56777, n56779, n56789, 
      n56791, n56795, n56801, n56803, n56813, n56815, n56819, n56825, n56827, 
      n56837, n56839, n56843, n56849, n56851, n56861, n56863, n56867, n56873, 
      n56875, n56885, n56887, n56891, n56897, n56899, n56909, n56911, n56915, 
      n56921, n56923, n56933, n56935, n56939, n56945, n56947, n56957, n56959, 
      n56963, n56969, n56971, n56981, n56983, n56987, n56993, n56995, n57005, 
      n57007, n57011, n57017, n57019, n57029, n57031, n57035, n57041, n57043, 
      n57053, n57055, n57059, n57065, n57067, n57077, n57079, n57083, n57089, 
      n57091, n57101, n57103, n57107, n57113, n57115, n57125, n57127, n57131, 
      n57137, n57139, n57149, n57151, n57155, n57161, n57163, n57173, n57175, 
      n57179, n57185, n57187, n57197, n57199, n57203, n57209, n57211, n57221, 
      n57223, n57227, n57233, n57235, n57245, n57247, n57251, n57257, n57259, 
      n57269, n57271, n57275, n57281, n57283, n57293, n57295, n57299, n57305, 
      n57307, n57317, n57319, n57323, n57329, n57331, n57341, n57343, n57347, 
      n57353, n57355, n57365, n57367, n57371, n57377, n57379, n57389, n57391, 
      n57395, n57401, n57403, n57413, n57415, n57419, n57425, n57427, n57437, 
      n57439, n57443, n57449, n57451, n57461, n57463, n57467, n57473, n57475, 
      n57485, n57487, n57491, n57497, n57499, n57509, n57511, n57515, n57521, 
      n57523, n57533, n57535, n57539, n57545, n57547, n57557, n57559, n57563, 
      n57569, n57571, n57581, n57583, n57587, n57593, n57595, n57605, n57607, 
      n57611, n57617, n57619, n57629, n57631, n57635, n57641, n57643, n57653, 
      n57659, n57665, n57667, n57677, n57683, n57689, n57691, n57701, n57707, 
      n57713, n57715, n57725, n57731, n57737, n57739, n57749, n57755, n57761, 
      n57763, n57773, n57779, n57785, n57787, n57797, n57803, n57809, n57811, 
      n57821, n57827, n57833, n57835, n57845, n57851, n57857, n57859, n57869, 
      n57875, n57881, n57883, n57893, n57899, n57905, n57907, n57917, n57923, 
      n57929, n57931, n57941, n57947, n57953, n57955, n57965, n57971, n57977, 
      n57979, n57989, n57995, n58001, n58003, n58013, n58028, n58036, n58041, 
      n58047, n58048, n58049, n58050, n58051, n58052, n58053, n58054, n58055, 
      n58056, n58057, n58058, n58059, n58060, n58061, n58062, n58063, n58064, 
      n58065, n58066, n58067, n58068, n58069, n58070, n58071, n58072, n58073, 
      n58074, n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082, 
      n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090, n58091, 
      n58092, n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100, 
      n58101, n58102, n58103, n58104, n58105, n58106, n58107, n58108, n58109, 
      n58110, n58112, n58114, n58116, n58118, n58120, n58122, n58124, n58126, 
      n58128, n58130, n58132, n58134, n58135, n58137, n58139, n58141, n58143, 
      n58145, n58147, n58149, n58151, n58153, n58155, n58157, n58159, n58161, 
      n58163, n58165, n58167, n58169, n58171, n58173, n58175, n58177, n58179, 
      n58181, n58183, n58185, n58187, n58189, n58191, n58193, n58195, n58197, 
      n58199, n58201, n58203, n58205, n58207, n58209, n58211, n58213, n58215, 
      n58217, n58219, n58221, n58223, n58225, n58227, n58229, n58231, n58232, 
      n58233, n58234, n58235, n58236, n58237, n58238, n58239, n58240, n58241, 
      n58242, n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250, 
      n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258, n58259, 
      n58260, n58261, n58262, n58263, n58264, n58265, n58266, n58267, n58268, 
      n58269, n58270, n58271, n58272, n58273, n58274, n58275, n58276, n58277, 
      n58278, n58279, n58280, n58281, n58282, n58283, n58284, n58285, n58286, 
      n58287, n58288, n58289, n58290, n58291, n58292, n58293, n58294, n58295, 
      n58297, n58299, n58301, n58303, n58304, n58305, n58306, n58307, n58308, 
      n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316, n58317, 
      n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325, n58326, 
      n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334, n58335, 
      n58336, n58337, n58338, n58339, n58340, n58341, n58342, n58343, n58344, 
      n58345, n58346, n58347, n58348, n58349, n58350, n58351, n58352, n58353, 
      n58354, n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362, 
      n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370, n58375, 
      n58376, n58377, n58378, n58379, n58380, n58381, n58382, n58383, n58384, 
      n58385, n58386, n58387, n58388, n58389, n58390, n58391, n58392, n58393, 
      n58394, n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402, 
      n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410, n58411, 
      n58412, n58413, n58414, n58415, n58416, n58417, n58418, n58419, n58420, 
      n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428, n58429, 
      n58430, n58431, n58432, n58433, n58434, n58435, n58436, n58437, n58438, 
      n58439, n58440, n58441, n58442, n58443, n58444, n58445, n58446, n58447, 
      n58448, n58449, n58450, n58451, n58452, n58453, n58454, n58455, n58456, 
      n58457, n58458, n58459, n58460, n58461, n58462, n58463, n58464, n58465, 
      n58466, n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474, 
      n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482, n58483, 
      n58484, n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492, 
      n58493, n58494, n58495, n58496, n58497, n58498, n58627, n58628, n58629, 
      n58630, n58631, n58632, n58633, n58634, n58635, n58636, n58637, n58638, 
      n58639, n58640, n58641, n58642, n58643, n58644, n58645, n58646, n58647, 
      n58648, n58649, n58650, n58651, n58652, n58653, n58654, n58667, n58668, 
      n58669, n58670, n58671, n58672, n58673, n58674, n58675, n58676, n58677, 
      n58678, n58679, n58680, n58681, n58682, n58683, n58684, n58685, n58686, 
      n58687, n58688, n58689, n58690, n58691, n58692, n58693, n58694, n58695, 
      n58696, n58697, n58698, n58699, n58700, n58701, n58702, n58703, n58704, 
      n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712, n58713, 
      n58714, n58715, n58716, n58717, n58718, n58731, n58732, n58733, n58734, 
      n58735, n58736, n58737, n58738, n58739, n58740, n58741, n58742, n58779, 
      n58780, n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788, 
      n58789, n58790, n58791, n58792, n58793, n58794, n58795, n58796, n58797, 
      n58798, n58799, n58800, n58801, n58802, n58803, n58804, n58805, n58806, 
      n58807, n58808, n58809, n58810, n58811, n58812, n58813, n58814, n58815, 
      n58816, n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824, 
      n58825, n58826, n58827, n58828, n58829, n58830, n58831, n58832, n58833, 
      n58834, n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842, 
      n58960, n59022, n59024, n59026, n59027, n59028, n59029, n59030, n59031, 
      n59032, n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040, 
      n59041, n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049, 
      n59050, n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058, 
      n59059, n59060, n59061, n59062, n59063, n59064, n59065, n59066, n59067, 
      n59068, n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076, 
      n59077, n59078, n59079, n59080, n59081, n59082, n59083, n59084, n59085, 
      n59086, n59087, n59088, n59089, n59090, n59091, n59092, n61957, n61958, 
      n61959, n61960, n61961, n61962, n61963, n61964, n61965, n61966, n61967, 
      n61968, n61969, n61970, n61971, n61972, n61973, n61974, n61975, n61976, 
      n61977, n61978, n61979, n61980, n61981, n61982, n61983, n61984, n61985, 
      n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993, n61994, 
      n61995, n61996, n61997, n61998, n61999, n62000, n62001, n62002, n62003, 
      n62004, n62005, n62006, n62007, n62008, n62009, n62010, n62011, n62012, 
      n62013, n62014, n62015, n62016, n62017, n62018, n62019, n62020, n62021, 
      n62022, n62023, n62024, n62025, n62026, n62027, n62028, n62029, n62030, 
      n62031, n62032, n62033, n62034, n62035, n62036, n62037, n62038, n62039, 
      n62040, n62041, n62042, n62043, n62044, n62045, n62046, n62047, n62048, 
      n62049, n62050, n62051, n62052, n62053, n62054, n62055, n62056, n62057, 
      n62058, n62059, n62060, n62061, n62062, n62063, n62064, n62065, n62066, 
      n62067, n62068, n62069, n62070, n62071, n62072, n62073, n62074, n62075, 
      n62076, n62077, n62078, n62079, n62080, n62081, n62082, n62083, n62084, 
      n62085, n62086, n62087, n62088, n62089, n62090, n62091, n62092, n62093, 
      n62094, n62095, n62096, n62097, n62098, n62099, n62100, n62101, n62102, 
      n62103, n62104, n62105, n62106, n62107, n62108, n62109, n62110, n62111, 
      n62112, n62113, n62114, n62115, n62116, n62117, n62118, n62119, n62120, 
      n62121, n62122, n62123, n62124, n62125, n62126, n62127, n62128, n62129, 
      n62130, n62131, n62132, n62133, n62134, n62135, n62136, n62137, n62138, 
      n62139, n62140, n62141, n62142, n62143, n62144, n62145, n62146, n62147, 
      n62148, n62149, n62150, n62151, n62152, n62153, n62154, n62155, n62156, 
      n62157, n62158, n62159, n62160, n62161, n62162, n62163, n62164, n62165, 
      n62166, n62167, n62168, n62169, n62170, n62171, n62172, n62173, n62174, 
      n62175, n62176, n62177, n62178, n62179, n62180, n62181, n62182, n62183, 
      n62184, n62185, n62186, n62187, n62188, n62189, n62190, n62191, n62192, 
      n62193, n62194, n62195, n62196, n62197, n62198, n62199, n62200, n62201, 
      n62202, n62203, n62204, n62205, n62206, n62207, n62208, n62209, n62210, 
      n62211, n62212, n62213, n62214, n62215, n62216, n62217, n62218, n62219, 
      n62220, n62221, n62222, n62223, n62224, n62225, n62226, n62227, n62228, 
      n62229, n62230, n62231, n62232, n62233, n62234, n62235, n62236, n62237, 
      n62238, n62239, n62240, n62241, n62242, n62243, n62244, n62245, n62246, 
      n62247, n62248, n62249, n62250, n62251, n62252, n62253, n62254, n62255, 
      n62256, n62257, n62258, n62259, n62260, n62261, n62262, n62263, n62264, 
      n62265, n62266, n62267, n62268, n62269, n62270, n62271, n62272, n62273, 
      n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281, n62282, 
      n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290, n62291, 
      n62292, n62293, n62294, n62295, n62296, n62297, n62298, n62299, n62300, 
      n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62308, n62309, 
      n62310, n62311, n62312, n62313, n62314, n62315, n62316, n62317, n62318, 
      n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326, n62327, 
      n62328, n62329, n62330, n62331, n62332, n62333, n62334, n62335, n62336, 
      n62337, n62338, n62339, n62340, n62341, n62342, n62343, n62344, n62345, 
      n62346, n62347, n62348, n62349, n62350, n62351, n62352, n62353, n62354, 
      n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362, n62363, 
      n62364, n62365, n62366, n62367, n62368, n62369, n62370, n62371, n62372, 
      n62373, n62374, n62375, n62376, n62377, n62378, n62379, n62380, n62381, 
      n62382, n62383, n62384, n62385, n62386, n62387, n62388, n62389, n62390, 
      n62391, n62392, n62393, n62394, n62395, n62396, n62397, n62398, n62399, 
      n62400, n62401, n62402, n62403, n62404, n62405, n62406, n62407, n62408, 
      n62409, n62410, n62411, n62412, n62413, n62414, n62415, n62416, n62417, 
      n62418, n62419, n62420, n62421, n62422, n62423, n62424, n62425, n62426, 
      n62427, n62428, n62429, n62430, n62431, n62432, n62433, n62434, n62435, 
      n62436, n62437, n62438, n62439, n62440, n62441, n62442, n62443, n62444, 
      n62445, n62446, n62447, n62448, n62449, n62450, n62451, n62452, n62453, 
      n62454, n62455, n62456, n62457, n62458, n62459, n62460, n62461, n62462, 
      n62463, n62464, n62465, n62466, n62467, n62468, n62469, n62470, n62471, 
      n62472, n62473, n62474, n62475, n62476, n62477, n62478, n62479, n62480, 
      n62481, n62482, n62483, n62484, n62485, n62486, n62487, n62488, n62489, 
      n62490, n62491, n62492, n62493, n62494, n62495, n62496, n62497, n62498, 
      n62499, n62500, n62501, n62502, n62503, n62504, n62505, n62506, n62507, 
      n62508, n62509, n62510, n62511, n62512, n62513, n62514, n62515, n62516, 
      n62517, n62518, n62519, n62520, n62521, n62522, n62523, n62524, n62525, 
      n62526, n62527, n62528, n62529, n62530, n62531, n62532, n62533, n62534, 
      n62535, n62536, n62537, n62538, n62539, n62540, n62541, n62542, n62543, 
      n62544, n62545, n62546, n62547, n62548, n62549, n62550, n62551, n62552, 
      n62553, n62554, n62555, n62556, n62557, n62558, n62559, n62560, n62561, 
      n62562, n62563, n62564, n62565, n62566, n62567, n62568, n62569, n62570, 
      n62571, n62572, n62573, n62574, n62575, n62576, n62577, n62578, n62579, 
      n62580, n62581, n62582, n62583, n62584, n62585, n62586, n62587, n62588, 
      n62589, n62590, n62591, n62592, n62593, n62594, n62595, n62596, n62597, 
      n62598, n62599, n62600, n62601, n62602, n62603, n62604, n62605, n62606, 
      n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614, n62615, 
      n62616, n62617, n62618, n62619, n62620, n62621, n62622, n62623, n62624, 
      n62625, n62626, n62627, n62628, n62629, n62630, n62631, n62632, n62633, 
      n62634, n62635, n62636, n62637, n62638, n62639, n62640, n62641, n62642, 
      n62643, n62644, n62645, n62646, n62647, n62648, n62649, n62650, n62651, 
      n62652, n62653, n62654, n62655, n62656, n62657, n62658, n62659, n62660, 
      n62661, n62662, n62663, n62664, n62665, n62666, n62667, n62668, n62669, 
      n62670, n62671, n62672, n62673, n62674, n62675, n62676, n62677, n62678, 
      n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686, n62687, 
      n62688, n62689, n62690, n62691, n62692, n62693, n62694, n62695, n62696, 
      n62697, n62698, n62699, n62700, n62701, n62702, n62703, n62704, n62705, 
      n62706, n62707, n62708, n62709, n62710, n62711, n62712, n62713, n62714, 
      n62715, n62716, n62717, n62718, n62719, n62720, n62721, n62722, n62723, 
      n62724, n62725, n62726, n62727, n62728, n62729, n62730, n62731, n62732, 
      n62733, n62734, n62735, n62736, n62737, n62738, n62739, n62740, n62741, 
      n62742, n62743, n62744, n62745, n62746, n62747, n62748, n62749, n62750, 
      n62751, n62752, n62753, n62754, n62755, n62756, n62757, n62758, n62759, 
      n62760, n62761, n62762, n62763, n62764, n62765, n62766, n62767, n62768, 
      n62769, n62770, n62771, n62772, n62773, n62774, n62775, n62776, n62777, 
      n62778, n62779, n62780, n62781, n62782, n62783, n62784, n62785, n62786, 
      n62787, n62788, n62789, n62790, n62791, n62792, n62793, n62794, n62795, 
      n62796, n62797, n62798, n62799, n62800, n62801, n62802, n62803, n62804, 
      n62805, n62806, n62807, n62808, n62809, n62810, n62811, n62812, n62813, 
      n62814, n62815, n62816, n62817, n62818, n62819, n62820, n62821, n62822, 
      n62823, n62824, n62825, n62826, n62827, n62828, n62829, n62830, n62831, 
      n62832, n62833, n62834, n62835, n62836, n62837, n62838, n62839, n62840, 
      n62841, n62842, n62843, n62844, n62845, n62846, n62847, n62848, n62849, 
      n62850, n62851, n62852, n62853, n62854, n62855, n62856, n62857, n62858, 
      n62859, n62860, n62861, n62862, n62863, n62864, n62865, n62866, n62867, 
      n62868, n62869, n62870, n62871, n62872, n62873, n62874, n62875, n62876, 
      n62877, n62878, n62879, n62880, n62881, n62882, n62883, n62884, n62885, 
      n62886, n62887, n62888, n62889, n62890, n62891, n62892, n62893, n62894, 
      n62895, n62896, n62897, n62898, n62899, n62900, n62901, n62902, n62903, 
      n62904, n62905, n62906, n62907, n62908, n62909, n62910, n62911, n62912, 
      n62913, n62914, n62915, n62916, n62917, n62918, n62919, n62920, n62921, 
      n62922, n62923, n62924, n62925, n62926, n62927, n62928, n62929, n62930, 
      n62931, n62932, n62933, n62934, n62935, n62936, n62937, n62938, n62939, 
      n62940, n62941, n62942, n62943, n62944, n62945, n62946, n62947, n62948, 
      n62949, n62950, n62951, n62952, n62953, n62954, n62955, n62956, n62957, 
      n62958, n62959, n62960, n62961, n62962, n62963, n62964, n62965, n62966, 
      n62967, n62968, n62969, n62970, n62971, n62972, n62973, n62974, n62975, 
      n62976, n62977, n62978, n62979, n62980, n62981, n62982, n62983, n62984, 
      n62985, n62986, n62987, n62988, n62989, n62990, n62991, n62992, n62993, 
      n62994, n62995, n62996, n62997, n62998, n62999, n63000, n63001, n63002, 
      n63003, n63004, n63005, n63006, n63007, n63008, n63009, n63010, n63011, 
      n63012, n63013, n63014, n63015, n63016, n63017, n63018, n63019, n63020, 
      n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028, n63029, 
      n63030, n63031, n63032, n63033, n63034, n63035, n63036, n63037, n63038, 
      n63039, n63040, n63041, n63042, n63043, n63044, n63045, n63046, n63047, 
      n63048, n63049, n63050, n63051, n63052, n63053, n63054, n63055, n63056, 
      n63057, n63058, n63059, n63060, n63061, n63062, n63063, n63064, n63065, 
      n63066, n63067, n63068, n63069, n63070, n63071, n63072, n63073, n63074, 
      n63075, n63076, n63077, n63078, n63079, n63080, n63081, n63082, n63083, 
      n63084, n63085, n63086, n63087, n63088, n63089, n63090, n63091, n63092, 
      n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100, n63101, 
      n63102, n63103, n63104, n63105, n63106, n63107, n63108, n63109, n63110, 
      n63111, n63112, n63113, n63114, n63115, n63116, n63117, n63118, n63119, 
      n63120, n63121, n63122, n63123, n63124, n63125, n63126, n63127, n63128, 
      n63129, n63130, n63131, n63132, n63133, n63134, n63135, n63136, n63137, 
      n63138, n63139, n63140, n63141, n63142, n63143, n63144, n63145, n63146, 
      n63147, n63148, n63149, n63150, n63151, n63152, n63153, n63154, n63155, 
      n63156, n63157, n63158, n63159, n63160, n63161, n63162, n63163, n63164, 
      n63165, n63166, n63167, n63168, n63169, n63170, n63171, n63172, n63173, 
      n63174, n63175, n63176, n63177, n63178, n63179, n63180, n63181, n63182, 
      n63183, n63184, n63185, n63186, n63187, n63188, n63189, n63190, n63191, 
      n63192, n63193, n63194, n63195, n63196, n63197, n63198, n63199, n63200, 
      n63201, n63202, n63203, n63204, n63205, n63206, n63207, n63208, n63209, 
      n63210, n63211, n63212, n63213, n63214, n63215, n63216, n63217, n63218, 
      n63219, n63220, n63221, n63222, n63223, n63224, n63225, n63226, n63227, 
      n63228, n63229, n63230, n63231, n63232, n63233, n63234, n63235, n63236, 
      n63237, n63238, n63239, n63240, n63241, n63242, n63243, n63244, n63245, 
      n63246, n63247, n63248, n63249, n63250, n63251, n63252, n63253, n63254, 
      n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262, n63263, 
      n63264, n63265, n63266, n63267, n63268, n63269, n63270, n63271, n63272, 
      n63273, n63274, n63275, n63276, n63277, n63278, n63279, n63280, n63281, 
      n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289, n63290, 
      n63291, n63292, n63293, n63294, n63295, n63296, n63297, n63298, n63299, 
      n63300, n63301, n63302, n63303, n63304, n63305, n63306, n63307, n63308, 
      n63309, n63310, n63311, n63312, n63313, n63314, n63315, n63316, n63317, 
      n63318, n63319, n63320, n63321, n63322, n63323, n63324, n63325, n63326, 
      n63327, n63328, n63329, n63330, n63331, n63332, n63333, n63334, n63335, 
      n63336, n63337, n63338, n63339, n63340, n63341, n63342, n63343, n63344, 
      n63345, n63346, n63347, n63348, n63349, n63350, n63351, n63352, n63353, 
      n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361, n63362, 
      n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370, n63371, 
      n63372, n63373, n63374, n63375, n63376, n63377, n63378, n63379, n63380, 
      n63381, n63382, n63383, n63384, n63385, n63386, n63387, n63388, n63389, 
      n63390, n63391, n63392, n63393, n63394, n63395, n63396, n63397, n63398, 
      n63399, n63400, n63401, n63402, n63403, n63404, n63405, n63406, n63407, 
      n63408, n63409, n63410, n63411, n63412, n63413, n63414, n63415, n63416, 
      n63417, n63418, n63419, n63420, n63421, n63422, n63423, n63424, n63425, 
      n63426, n63427, n63428, n63429, n63430, n63431, n63432, n63433, n63434, 
      n63435, n63436, n63437, n63438, n63439, n63440, n63441, n63442, n63443, 
      n63444, n63445, n63446, n63447, n63448, n63449, n63450, n63451, n63452, 
      n63453, n63454, n63455, n63456, n63457, n63458, n63459, n63460, n63461, 
      n63462, n63463, n63464, n63465, n63466, n63467, n63468, n63469, n63470, 
      n63471, n63472, n63473, n63474, n63475, n63476, n63477, n63478, n63479, 
      n63480, n63481, n63482, n63483, n63484, n63485, n63486, n63487, n63488, 
      n63489, n63490, n63491, n63492, n63493, n63494, n63495, n63496, n63497, 
      n63498, n63499, n63500, n63501, n63502, n63503, n63504, n63505, n63506, 
      n63507, n63508, n63509, n63510, n63511, n63512, n63513, n63514, n63515, 
      n63516, n63517, n63518, n63519, n63520, n63521, n63522, n63523, n63524, 
      n63525, n63526, n63527, n63528, n63529, n63530, n63531, n63532, n63533, 
      n63534, n63535, n63536, n63537, n63538, n63539, n63540, n63541, n63542, 
      n63543, n63544, n63545, n63546, n63547, n63548, n63549, n63550, n63551, 
      n63552, n63553, n63554, n63555, n63556, n63557, n63558, n63559, n63560, 
      n63561, n63562, n63563, n63564, n63565, n63566, n63567, n63568, n63569, 
      n63570, n63571, n63572, n63573, n63574, n63575, n63576, n63577, n63578, 
      n63579, n63580, n63581, n63582, n63583, n63584, n63585, n63586, n63587, 
      n63588, n63589, n63590, n63591, n63592, n63593, n63594, n63595, n63596, 
      n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604, n63605, 
      n63606, n63607, n63608, n63609, n63610, n63611, n63612, n63613, n63614, 
      n63615, n63616, n63617, n63618, n63619, n63620, n63621, n63622, n63623, 
      n63624, n63625, n63626, n63627, n63628, n63629, n63630, n63631, n63632, 
      n63633, n63634, n63635, n63636, n63637, n63638, n63639, n63640, n63641, 
      n63642, n63643, n63644, n63645, n63646, n63647, n63648, n63649, n63650, 
      n63651, n63652, n63653, n63654, n63655, n63656, n63657, n63658, n63659, 
      n63660, n63661, n63662, n63663, n63664, n63665, n63666, n63667, n63668, 
      n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676, n63677, 
      n63678, n63679, n63680, n63681, n63682, n63683, n63684, n63685, n63686, 
      n63687, n63688, n63689, n63690, n63691, n63692, n63693, n63694, n63695, 
      n63696, n63697, n63698, n63699, n63700, n63701, n63702, n63703, n63704, 
      n63705, n63706, n63707, n63708, n63709, n63710, n63711, n63712, n63713, 
      n63714, n63715, n63716, n63717, n63718, n63719, n63720, n63721, n63722, 
      n63723, n63724, n63725, n63726, n63727, n63728, n63729, n63730, n63731, 
      n63732, n63733, n63734, n63735, n63736, n63737, n63738, n63739, n63740, 
      n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748, n63749, 
      n63750, n63751, n63752, n63753, n63754, n63755, n63756, n63757, n63758, 
      n63759, n63760, n63761, n63762, n63763, n63764, n63765, n63766, n63767, 
      n63768, n63769, n63770, n63771, n63772, n63773, n63774, n63775, n63776, 
      n63777, n63778, n63780, n63781, n63782, n63783, n63784, n63785, n63786, 
      n63787, n63788, n63790, n63791, n63792, n63793, n63794, n63795, n63797, 
      n63798, n63799, n63800, n63801, n63802, n63803, n63804, n63805, n63806, 
      n63807, n63808, n63809, n63810, n63811, n63812, n63813, n63814, n63815, 
      n63816, n63817, n63818, n63819, n63820, n63821, n63822, n63823, n63824, 
      n63825, n63826, n63827, n63828, n63829, n63830, n63831, n63833, n63835, 
      n63836, n63837, n63838, n63839, n63840, n63841, n63842, n63843, n63844, 
      n63845, n63846, n63847, n63848, n63849, n63850, n63851, n63852, n63854, 
      n63856, n63857, n63858, n63859, n63860, n63861, n63862, n63863, n63864, 
      n63865, n63866, n63867, n63868, n63869, n63870, n63871, n63872, n63873, 
      n63875, n63877, n63878, n63879, n63880, n63881, n63882, n63883, n63884, 
      n63885, n63886, n63887, n63888, n63889, n63890, n63891, n63892, n63893, 
      n63894, n63896, n63897, n63898, n63899, n63900, n63901, n63902, n63903, 
      n63904, n63905, n63906, n63907, n63908, n63909, n63910, n63911, n63912, 
      n63913, n63914, n63916, n63917, n63918, n63919, n63920, n63921, n63922, 
      n63923, n63924, n63925, n63926, n63927, n63928, n63929, n63930, n63931, 
      n63932, n63933, n63934, n63936, n63937, n63938, n63939, n63940, n63941, 
      n63942, n63943, n63944, n63945, n63946, n63947, n63948, n63949, n63950, 
      n63951, n63952, n63953, n63954, n63956, n63957, n63958, n63959, n63960, 
      n63961, n63962, n63963, n63964, n63965, n63966, n63967, n63968, n63969, 
      n63970, n63971, n63972, n63973, n63974, n63976, n63977, n63978, n63979, 
      n63980, n63981, n63982, n63983, n63984, n63985, n63986, n63987, n63988, 
      n63989, n63990, n63991, n63992, n63993, n63994, n63996, n63997, n63998, 
      n63999, n64000, n64001, n64002, n64003, n64004, n64005, n64006, n64007, 
      n64008, n64009, n64010, n64011, n64012, n64013, n64014, n64016, n64017, 
      n64018, n64019, n64020, n64021, n64022, n64023, n64024, n64025, n64026, 
      n64027, n64028, n64029, n64030, n64031, n64032, n64033, n64034, n64036, 
      n64037, n64038, n64039, n64040, n64041, n64042, n64043, n64044, n64045, 
      n64046, n64047, n64048, n64049, n64050, n64051, n64052, n64053, n64054, 
      n64056, n64057, n64058, n64059, n64060, n64061, n64062, n64063, n64064, 
      n64065, n64066, n64067, n64068, n64069, n64070, n64071, n64072, n64073, 
      n64074, n64076, n64077, n64078, n64079, n64080, n64081, n64082, n64083, 
      n64084, n64085, n64086, n64087, n64088, n64089, n64090, n64091, n64092, 
      n64093, n64094, n64096, n64097, n64098, n64099, n64100, n64101, n64102, 
      n64103, n64104, n64105, n64106, n64107, n64108, n64109, n64110, n64111, 
      n64112, n64113, n64114, n64116, n64117, n64118, n64119, n64120, n64121, 
      n64122, n64123, n64124, n64125, n64126, n64127, n64128, n64129, n64130, 
      n64131, n64132, n64133, n64134, n64136, n64137, n64138, n64139, n64140, 
      n64141, n64142, n64143, n64144, n64145, n64146, n64147, n64148, n64149, 
      n64150, n64151, n64152, n64153, n64154, n64156, n64157, n64158, n64159, 
      n64160, n64161, n64162, n64163, n64164, n64165, n64166, n64167, n64168, 
      n64169, n64170, n64171, n64172, n64173, n64174, n64176, n64177, n64178, 
      n64179, n64180, n64181, n64182, n64183, n64184, n64185, n64186, n64187, 
      n64188, n64189, n64190, n64191, n64192, n64193, n64194, n64196, n64197, 
      n64198, n64199, n64200, n64201, n64202, n64203, n64204, n64205, n64206, 
      n64207, n64208, n64209, n64210, n64211, n64212, n64213, n64214, n64216, 
      n64217, n64218, n64219, n64220, n64221, n64222, n64223, n64224, n64225, 
      n64226, n64227, n64228, n64229, n64230, n64231, n64232, n64233, n64234, 
      n64236, n64237, n64238, n64239, n64240, n64241, n64242, n64243, n64244, 
      n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64252, n64253, 
      n64254, n64256, n64257, n64258, n64259, n64260, n64261, n64262, n64263, 
      n64264, n64265, n64266, n64267, n64268, n64269, n64270, n64271, n64272, 
      n64273, n64274, n64276, n64277, n64278, n64279, n64280, n64281, n64282, 
      n64283, n64284, n64285, n64286, n64287, n64288, n64289, n64290, n64291, 
      n64292, n64293, n64294, n64296, n64297, n64298, n64299, n64300, n64301, 
      n64302, n64303, n64304, n64305, n64306, n64307, n64308, n64309, n64310, 
      n64311, n64312, n64313, n64314, n64316, n64317, n64318, n64319, n64320, 
      n64321, n64322, n64323, n64324, n64325, n64326, n64327, n64328, n64329, 
      n64330, n64331, n64332, n64333, n64334, n64336, n64337, n64338, n64339, 
      n64340, n64341, n64342, n64343, n64344, n64345, n64346, n64347, n64348, 
      n64349, n64350, n64351, n64352, n64353, n64354, n64356, n64357, n64358, 
      n64359, n64360, n64361, n64362, n64363, n64364, n64365, n64366, n64367, 
      n64368, n64369, n64370, n64371, n64372, n64373, n64374, n64376, n64377, 
      n64378, n64379, n64380, n64381, n64382, n64383, n64384, n64385, n64386, 
      n64387, n64388, n64389, n64390, n64391, n64392, n64393, n64394, n64396, 
      n64397, n64398, n64399, n64400, n64401, n64402, n64403, n64404, n64405, 
      n64406, n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414, 
      n64416, n64417, n64418, n64419, n64420, n64421, n64422, n64423, n64424, 
      n64425, n64426, n64427, n64428, n64429, n64430, n64431, n64432, n64433, 
      n64434, n64436, n64437, n64438, n64439, n64440, n64441, n64442, n64443, 
      n64444, n64445, n64446, n64447, n64448, n64449, n64450, n64451, n64452, 
      n64453, n64454, n64456, n64457, n64458, n64459, n64460, n64461, n64462, 
      n64463, n64464, n64465, n64466, n64467, n64468, n64469, n64470, n64471, 
      n64472, n64473, n64474, n64476, n64477, n64478, n64479, n64480, n64481, 
      n64482, n64483, n64484, n64485, n64486, n64487, n64488, n64489, n64490, 
      n64491, n64492, n64493, n64494, n64496, n64497, n64498, n64499, n64500, 
      n64501, n64502, n64503, n64504, n64505, n64506, n64507, n64508, n64509, 
      n64510, n64511, n64512, n64513, n64514, n64516, n64517, n64518, n64519, 
      n64520, n64521, n64522, n64523, n64524, n64525, n64526, n64527, n64528, 
      n64529, n64530, n64531, n64532, n64533, n64534, n64536, n64537, n64538, 
      n64539, n64540, n64541, n64542, n64543, n64544, n64545, n64546, n64547, 
      n64548, n64549, n64550, n64551, n64552, n64553, n64554, n64556, n64557, 
      n64558, n64559, n64560, n64561, n64562, n64563, n64564, n64565, n64566, 
      n64567, n64568, n64569, n64570, n64571, n64572, n64573, n64574, n64576, 
      n64577, n64578, n64579, n64580, n64581, n64582, n64583, n64584, n64585, 
      n64586, n64587, n64588, n64589, n64590, n64591, n64592, n64593, n64594, 
      n64596, n64597, n64598, n64599, n64600, n64601, n64602, n64603, n64604, 
      n64605, n64606, n64607, n64608, n64609, n64610, n64611, n64612, n64613, 
      n64614, n64616, n64617, n64618, n64619, n64620, n64621, n64622, n64623, 
      n64624, n64625, n64626, n64627, n64628, n64629, n64630, n64631, n64632, 
      n64633, n64634, n64636, n64637, n64638, n64639, n64640, n64641, n64642, 
      n64643, n64644, n64645, n64646, n64647, n64648, n64649, n64650, n64651, 
      n64652, n64653, n64654, n64656, n64657, n64658, n64659, n64660, n64661, 
      n64662, n64663, n64664, n64665, n64666, n64667, n64668, n64669, n64670, 
      n64671, n64672, n64673, n64674, n64676, n64677, n64678, n64679, n64680, 
      n64681, n64682, n64683, n64684, n64685, n64686, n64687, n64688, n64689, 
      n64690, n64691, n64692, n64693, n64694, n64696, n64697, n64698, n64699, 
      n64700, n64701, n64702, n64703, n64704, n64705, n64706, n64707, n64708, 
      n64709, n64710, n64711, n64712, n64713, n64714, n64716, n64717, n64718, 
      n64719, n64720, n64721, n64722, n64723, n64724, n64725, n64726, n64727, 
      n64728, n64729, n64730, n64731, n64732, n64733, n64734, n64736, n64737, 
      n64738, n64739, n64740, n64741, n64742, n64743, n64744, n64745, n64746, 
      n64747, n64748, n64749, n64750, n64751, n64752, n64753, n64754, n64756, 
      n64757, n64758, n64759, n64760, n64761, n64762, n64763, n64764, n64765, 
      n64766, n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774, 
      n64776, n64777, n64778, n64779, n64780, n64781, n64782, n64783, n64784, 
      n64785, n64786, n64787, n64788, n64789, n64790, n64791, n64792, n64793, 
      n64794, n64796, n64797, n64798, n64799, n64800, n64801, n64802, n64803, 
      n64804, n64805, n64806, n64807, n64808, n64809, n64810, n64811, n64812, 
      n64813, n64814, n64816, n64817, n64818, n64819, n64820, n64821, n64822, 
      n64823, n64824, n64825, n64826, n64827, n64828, n64829, n64830, n64831, 
      n64832, n64833, n64834, n64836, n64837, n64838, n64839, n64840, n64841, 
      n64842, n64843, n64844, n64845, n64846, n64847, n64848, n64849, n64850, 
      n64851, n64852, n64853, n64854, n64855, n64856, n64857, n64858, n64859, 
      n64860, n64861, n64862, n64863, n64864, n64865, n64866, n64867, n64868, 
      n64869, n64870, n64871, n64872, n64873, n64874, n64875, n64876, n64877, 
      n64878, n64879, n64880, n64881, n64882, n64883, n64884, n64885, n64886, 
      n64887, n64888, n64889, n64890, n64891, n64892, n64893, n64894, n64895, 
      n64896, n64897, n64898, n64899, n64900, n64901, n64902, n64903, n64904, 
      n64905, n64906, n64907, n64908, n64909, n64910, n64911, n64912, n64913, 
      n64914, n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922, 
      n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930, n64931, 
      n64932, n64933, n64934, n64935, n64936, n64937, n64938, n64939, n64940, 
      n64941, n64942, n64943, n64944, n64945, n64946, n64947, n64948, n64949, 
      n64950, n64951, n64952, n64953, n64954, n64955, n64956, n64957, n64958, 
      n64959, n64960, n64961, n64962, n64963, n64964, n64965, n64966, n64967, 
      n64968, n64969, n64970, n64971, n64972, n64973, n64974, n64975, n64976, 
      n64977, n64978, n64979, n64980, n64981, n64982, n64983, n64984, n64985, 
      n64986, n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994, 
      n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002, n65003, 
      n65004, n65005, n65006, n65007, n65008, n65009, n65010, n65011, n65012, 
      n65013, n65014, n65015, n65016, n65017, n65018, n65019, n65020, n65021, 
      n65022, n65023, n65024, n65025, n65026, n65027, n65028, n65029, n65030, 
      n65031, n65032, n65033, n65034, n65035, n65036, n65037, n65038, n65039, 
      n65040, n65041, n65042, n65043, n65044, n65045, n65046, n65047, n65048, 
      n65049, n65050, n65051, n65052, n65053, n65054, n65055, n65056, n65057, 
      n65058, n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066, 
      n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074, n65075, 
      n65076, n65077, n65078, n65079, n65080, n65081, n65082, n65083, n65084, 
      n65085, n65086, n65087, n65088, n65089, n65090, n65091, n65092, n65093, 
      n65094, n65095, n65096, n65098, n65099, n65100, n65101, n65102, n65103, 
      n65104, n65105, n65106, n65107, n65108, n65109, n65110, n65111, n65112, 
      n65113, n65114, n65115, n65116, n65117, n65118, n65119, n65120, n65121, 
      n65122, n65123, n65124, n65125, n65126, n65127, n65128, n65129, n65130, 
      n65131, n65132, n65133, n65134, n65135, n65136, n65137, n65138, n65139, 
      n65140, n65141, n65142, n65143, n65144, n65145, n65146, n65147, n65148, 
      n65149, n65150, n65151, n65152, n65153, n65154, n65155, n65156, n65157, 
      n65158, n65159, n65160, n65161, n65162, n65163, n65164, n65165, n65166, 
      n65167, n65168, n65169, n65170, n65171, n65172, n65173, n65174, n65175, 
      n65176, n65177, n65178, n65179, n65180, n65181, n65182, n65183, n65184, 
      n65185, n65186, n65187, n65188, n65189, n65190, n65191, n65192, n65193, 
      n65194, n65195, n65196, n65197, n65198, n65199, n65200, n65201, n65202, 
      n65203, n65204, n65205, n65206, n65207, n65208, n65209, n65210, n65211, 
      n65212, n65213, n65214, n65215, n65216, n65217, n65218, n65219, n65220, 
      n65221, n65222, n65223, n65224, n65225, n65226, n65227, n65228, n65229, 
      n65230, n65231, n65232, n65233, n65234, n65235, n65236, n65237, n65238, 
      n65239, n65240, n65241, n65242, n65243, n65244, n65245, n65246, n65247, 
      n65248, n65249, n65250, n65251, n65252, n65253, n65254, n65255, n65256, 
      n65257, n65258, n65259, n65260, n65261, n65262, n65263, n65264, n65265, 
      n65266, n65267, n65268, n65269, n65270, n65271, n65272, n65273, n65274, 
      n65275, n65276, n65277, n65278, n65279, n65280, n65281, n65282, n65283, 
      n65284, n65285, n65286, n65287, n65288, n65289, n65290, n65291, n65292, 
      n65293, n65294, n65295, n65296, n65297, n65298, n65299, n65300, n65301, 
      n65302, n65303, n65304, n65305, n65306, n65307, n65308, n65309, n65310, 
      n65311, n65312, n65313, n65314, n65315, n65316, n65317, n65318, n65319, 
      n65320, n65321, n65322, n65323, n65324, n65325, n65326, n65327, n65328, 
      n65329, n65330, n65331, n65332, n65333, n65334, n65335, n65336, n65337, 
      n65338, n65339, n65340, n65341, n65342, n65343, n65344, n65345, n65346, 
      n65347, n65348, n65349, n65350, n65351, n65352, n65353, n65354, n65355, 
      n65356, n65357, n65358, n65359, n65360, n65361, n65362, n65363, n65364, 
      n65365, n65366, n65367, n65368, n65369, n65370, n65371, n65372, n65373, 
      n65374, n65375, n65376, n65377, n65378, n65379, n65380, n65381, n65382, 
      n65383, n65384, n65385, n65386, n65387, n65388, n65389, n65390, n65391, 
      n65392, n65393, n65394, n65395, n65396, n65397, n65398, n65399, n65400, 
      n65401, n65402, n65403, n65404, n65405, n65406, n65407, n65408, n65409, 
      n65410, n65411, n65412, n65413, n65414, n65415, n65416, n65417, n65418, 
      n65419, n65420, n65421, n65422, n65423, n65424, n65425, n65426, n65427, 
      n65428, n65429, n65430, n65431, n65432, n65433, n65434, n65435, n65436, 
      n65437, n65438, n65439, n65440, n65441, n65442, n65443, n65444, n65445, 
      n65446, n65447, n65448, n65449, n65450, n65451, n65452, n65453, n65454, 
      n65455, n65456, n65457, n65458, n65459, n65460, n65461, n65462, n65463, 
      n65464, n65465, n65466, n65467, n65468, n65469, n65470, n65471, n65472, 
      n65473, n65474, n65475, n65476, n65477, n65478, n65479, n65480, n65481, 
      n65482, n65483, n65484, n65485, n65486, n65487, n65488, n65489, n65490, 
      n65491, n65492, n65493, n65494, n65495, n65496, n65497, n65498, n65499, 
      n65500, n65501, n65502, n65503, n65504, n65505, n65506, n65507, n65508, 
      n65509, n65510, n65511, n65512, n65513, n65514, n65515, n65516, n65517, 
      n65518, n65519, n65520, n65521, n65522, n65523, n65524, n65525, n65526, 
      n65527, n65528, n65529, n65530, n65531, n65532, n65533, n65534, n65535, 
      n65536, n65537, n65538, n65539, n65540, n65541, n65542, n65543, n65544, 
      n65545, n65546, n65547, n65548, n65549, n65550, n65551, n65552, n65553, 
      n65554, n65555, n65556, n65557, n65558, n65559, n65560, n65561, n65562, 
      n65563, n65564, n65565, n65566, n65567, n65568, n65569, n65570, n65571, 
      n65572, n65573, n65574, n65575, n65576, n65577, n65578, n65579, n65580, 
      n65581, n65582, n65583, n65584, n65585, n65586, n65587, n65588, n65589, 
      n65590, n65591, n65592, n65593, n65594, n65595, n65596, n65597, n65598, 
      n65599, n65600, n65601, n65602, n65603, n65604, n65605, n65606, n65607, 
      n65608, n65609, n65610, n65611, n65612, n65613, n65614, n65615, n65616, 
      n65617, n65618, n65619, n65620, n65621, n65622, n65623, n65624, n65625, 
      n65626, n65627, n65628, n65629, n65630, n65631, n65632, n65633, n65634, 
      n65635, n65636, n65637, n65638, n65639, n65640, n65641, n65642, n65643, 
      n65644, n65645, n65646, n65647, n65648, n65649, n65650, n65651, n65652, 
      n65653, n65654, n65655, n65656, n65657, n65658, n65659, n65660, n65661, 
      n65662, n65663, n65664, n65665, n65666, n65667, n65668, n65669, n65670, 
      n65671, n65672, n65673, n65674, n65675, n65676, n65677, n65678, n65679, 
      n65680, n65681, n65682, n65683, n65684, n65685, n65686, n65687, n65688, 
      n65689, n65690, n65691, n65692, n65693, n65694, n65695, n65696, n65697, 
      n65698, n65699, n65700, n65701, n65702, n65703, n65704, n65705, n65706, 
      n65707, n65708, n65709, n65710, n65711, n65712, n65713, n65714, n65715, 
      n65716, n65717, n65718, n65719, n65720, n65721, n65722, n65723, n65724, 
      n65725, n65726, n65727, n65728, n65729, n65730, n65731, n65732, n65733, 
      n65734, n65735, n65736, n65737, n65738, n65739, n65740, n65741, n65742, 
      n65743, n65744, n65745, n65746, n65747, n65748, n65749, n65750, n65751, 
      n65752, n65753, n65754, n65755, n65756, n65757, n65758, n65759, n65760, 
      n65761, n65762, n65763, n65764, n65765, n65766, n65767, n65768, n65769, 
      n65770, n65771, n65772, n65773, n65774, n65775, n65776, n65777, n65778, 
      n65779, n65780, n65781, n65782, n65783, n65784, n65785, n65786, n65787, 
      n65788, n65789, n65790, n65791, n65792, n65793, n65794, n65795, n65796, 
      n65797, n65798, n65799, n65800, n65801, n65802, n65803, n65804, n65805, 
      n65806, n65807, n65808, n65809, n65810, n65811, n65812, n65813, n65814, 
      n65815, n65816, n65817, n65818, n65819, n65820, n65821, n65822, n65823, 
      n65824, n65825, n65826, n65827, n65828, n65829, n65830, n65831, n65832, 
      n65833, n65834, n65835, n65836, n65837, n65838, n65839, n65840, n65841, 
      n65842, n65843, n65844, n65845, n65846, n65847, n65848, n65849, n65850, 
      n65851, n65852, n65853, n65854, n65855, n65856, n65857, n65858, n65859, 
      n65860, n65861, n65862, n65863, n65864, n65865, n65866, n65867, n65868, 
      n65869, n65870, n65871, n65872, n65873, n65874, n65875, n65876, n65877, 
      n65878, n65879, n65880, n65881, n65882, n65883, n65884, n65885, n65886, 
      n65887, n65888, n65889, n65890, n65891, n65892, n65893, n65894, n65895, 
      n65896, n65897, n65898, n65899, n65900, n65901, n65902, n65903, n65904, 
      n65905, n65906, n65907, n65908, n65909, n65910, n65911, n65912, n65913, 
      n65914, n65915, n65916, n65917, n65918, n65919, n65920, n65921, n65922, 
      n65923, n65924, n65925, n65926, n65927, n65928, n65929, n65930, n65931, 
      n65932, n65933, n65934, n65935, n65936, n65937, n65938, n65939, n65940, 
      n65941, n65942, n65943, n65944, n65945, n65946, n65947, n65948, n65949, 
      n65950, n65951, n65952, n65953, n65954, n65955, n65956, n65957, n65958, 
      n65959, n65960, n65961, n65962, n65963, n65964, n65965, n65966, n65967, 
      n65968, n65969, n65970, n65971, n65972, n65973, n65974, n65975, n65976, 
      n65977, n65978, n65979, n65980, n65981, n65982, n65983, n65984, n65985, 
      n65986, n65987, n65988, n65989, n65990, n65991, n65992, n65993, n65994, 
      n65995, n65996, n65997, n65998, n65999, n66000, n66001, n66002, n66003, 
      n66004, n66005, n66006, n66007, n66008, n66009, n66010, n66011, n66012, 
      n66013, n66014, n66015, n66016, n66017, n66018, n66019, n66020, n66021, 
      n66022, n66023, n66024, n66025, n66026, n66027, n66028, n66029, n66030, 
      n66031, n66032, n66033, n66034, n66035, n66036, n66037, n66038, n66039, 
      n66040, n66041, n66042, n66043, n66044, n66045, n66046, n66047, n66048, 
      n66049, n66050, n66051, n66052, n66053, n66054, n66055, n66056, n66057, 
      n66058, n66059, n66060, n66061, n66062, n66063, n66064, n66065, n66066, 
      n66067, n66068, n66069, n66070, n66071, n66072, n66073, n66074, n66075, 
      n66076, n66077, n66078, n66079, n66080, n66081, n66082, n66083, n66084, 
      n66085, n66086, n66087, n66088, n66089, n66090, n66091, n66092, n66093, 
      n66094, n66095, n66096, n66097, n66098, n66099, n66100, n66101, n66102, 
      n66103, n66104, n66105, n66106, n66107, n66108, n66109, n66110, n66111, 
      n66112, n66113, n66114, n66115, n66116, n66117, n66118, n66119, n66120, 
      n66121, n66122, n66123, n66124, n66125, n66126, n66127, n66128, n66129, 
      n66130, n66131, n66132, n66133, n66134, n66135, n66136, n66137, n66138, 
      n66139, n66140, n66141, n66142, n66143, n66144, n66145, n66146, n66147, 
      n66148, n66149, n66150, n66151, n66152, n66153, n66154, n66155, n66156, 
      n66157, n66158, n66159, n66160, n66161, n66162, n66163, n66164, n66165, 
      n66166, n66167, n66168, n66169, n66170, n66171, n66172, n66173, n66174, 
      n66175, n66176, n66177, n66178, n66179, n66180, n66181, n66182, n66183, 
      n66184, n66185, n66186, n66187, n66188, n66189, n66190, n66191, n66192, 
      n66193, n66194, n66195, n66196, n66197, n66198, n66199, n66200, n66201, 
      n66202, n66203, n66204, n66205, n66206, n66207, n66208, n66209, n66210, 
      n66211, n66212, n66213, n66214, n66215, n66216, n66217, n66218, n66219, 
      n66220, n66221, n66222, n66223, n66224, n66225, n66226, n66227, n66228, 
      n66229, n66230, n66231, n66232, n66233, n66234, n66235, n66236, n66237, 
      n66238, n66239, n66240, n66241, n66242, n66243, n66244, n66245, n66246, 
      n66247, n66248, n66249, n66250, n66251, n66252, n66253, n66254, n66255, 
      n66256, n66257, n66258, n66259, n66260, n66261, n66262, n66263, n66264, 
      n66265, n66266, n66267, n66268, n66269, n66270, n66271, n66272, n66273, 
      n66274, n66275, n66276, n66277, n66278, n66279, n66280, n66281, n66282, 
      n66283, n66284, n66285, n66286, n66287, n66288, n66289, n66290, n66291, 
      n66292, n66293, n66294, n66295, n66296, n66297, n66298, n66299, n66300, 
      n66301, n66305, n66306, n66307, n66308, n66313, n66314, n66315, n66316, 
      n66317, n66318, n66319, n66320, n66321, n66322, n66323, n66324, n66325, 
      n66326, n66327, n66328, n66329, n66330, n66331, n66332, n66333, n66334, 
      n66335, n66336, n66337, n66338, n66339, n66340, n66341, n66342, n66343, 
      n66344, n66345, n66346, n66347, n66348, n66349, n66350, n66351, n66352, 
      n66353, n66354, n66355, n66356, n66357, n66358, n66359, n66360, n66361, 
      n66362, n66363, n66364, n66365, n66366, n66367, n66368, n66369, n66370, 
      n66371, n66372, n66494, n66495, n66496, n66497, n66498, n66499, n66500, 
      n66501, n66502, n66503, n66504, n66505, n66506, n66507, n66508, n66509, 
      n66510, n66511, n66512, n66513, n66514, n66515, n66516, n66517, n66518, 
      n66519, n66520, n66521, n66522, n66523, n66524, n66525, n66526, n66527, 
      n66528, n66529, n66530, n66531, n66532, n66533, n66534, n66535, n66536, 
      n66537, n66538, n66539, n66540, n66541, n66542, n66543, n66544, n66545, 
      n66546, n66547, n66548, n66549, n66550, n66551, n66552, n66553, n66554, 
      n66555, n66556, n66557, n66558, n66559, n66560, n66561, n66562, n66563, 
      n66564, n66565, n66566, n66567, n66568, n66569, n66570, n66571, n66572, 
      n66573, n66574, n66575, n66576, n66577, n66578, n66579, n66580, n66581, 
      n66582, n66583, n66584, n66585, n66586, n66587, n66588, n66589, n66590, 
      n66591, n66592, n66593, n66594, n66595, n66596, n66597, n66598, n66599, 
      n66600, n66601, n66602, n66603, n66604, n66605, n66606, n66607, n66608, 
      n66609, n66610, n66611, n66612, n66613, n66614, n66615, n66616, n66617, 
      n66618, n66619, n66620, n66621, n66622, n66623, n66624, n66625, n66626, 
      n66627, n66628, n66629, n66630, n66631, n66632, n66633, n66634, n66635, 
      n66636, n66637, n66638, n66639, n66640, n66641, n66642, n66643, n66644, 
      n66645, n66646, n66647, n66648, n66649, n66650, n66651, n66652, n66653, 
      n66654, n66655, n66656, n66657, n66658, n66659, n66660, n66661, n66662, 
      n66663, n66664, n66665, n66666, n66667, n66668, n66669, n66670, n66671, 
      n66672, n66673, n66674, n66675, n66676, n66677, n66678, n66679, n66680, 
      n66681, n66682, n66683, n66684, n66685, n66686, n66687, n66688, n66689, 
      n66690, n66691, n66692, n66693, n66694, n66695, n66696, n66697, n66698, 
      n66699, n66700, n66701, n66702, n66703, n66704, n66705, n66706, n66707, 
      n66708, n66709, n66710, n66711, n66712, n66713, n66714, n66715, n66716, 
      n66717, n66718, n66719, n66720, n66721, n66722, n66723, n66724, n66725, 
      n66726, n66727, n66728, n66729, n66730, n66731, n66732, n66733, n66734, 
      n66735, n66736, n66737, n66738, n66739, n66740, n66741, n66742, n66743, 
      n66744, n66745, n66746, n66747, n66748, n66749, n66750, n66751, n66752, 
      n66753, n66754, n66755, n66756, n66757, n66758, n66759, n66760, n66761, 
      n66762, n66763, n66764, n66765, n66766, n66767, n66768, n66769, n66770, 
      n66771, n66772, n66773, n66774, n66775, n66776, n66777, n66778, n66779, 
      n66780, n66781, n66782, n66783, n66784, n66785, n66786, n66787, n66788, 
      n66789, n66790, n66791, n66792, n66793, n66794, n66795, n66796, n66797, 
      n66798, n66799, n66800, n66801, n66802, n66803, n66804, n66805, n66806, 
      n66807, n66808, n66809, n66810, n66811, n66812, n66813, n66814, n66815, 
      n66816, n66817, n66818, n66819, n66820, n66821, n66822, n66823, n66824, 
      n66825, n66826, n66827, n66828, n66829, n66830, n66831, n66832, n66833, 
      n66834, n66835, n66836, n66837, n66838, n66839, n66840, n66841, n66842, 
      n66843, n66844, n66845, n66846, n66847, n66848, n66849, n66850, n66851, 
      n66852, n66853, n66854, n66855, n66856, n66857, n66858, n66859, n66860, 
      n66861, n66862, n66863, n66864, n66865, n66866, n66867, n66868, n66869, 
      n66870, n66871, n66872, n66873, n66874, n66875, n66876, n66877, n66878, 
      n66879, n66880, n66881, n66882, n66883, n66884, n66885, n66886, n66887, 
      n66888, n66889, n66890, n66891, n66892, n66893, n66894, n66895, n66896, 
      n66897, n66898, n66899, n66900, n66901, n66902, n66903, n66904, n66905, 
      n66906, n66907, n66908, n66909, n66910, n66911, n66912, n66913, n66914, 
      n66915, n66916, n66917, n66918, n66919, n66920, n66921, n66922, n66923, 
      n66924, n66925, n66926, n66927, n66928, n66929, n66930, n66931, n66932, 
      n66933, n66934, n66935, n66936, n66937, n66938, n66939, n66940, n66941, 
      n66942, n66943, n66944, n66945, n66946, n66947, n66948, n66949, n66950, 
      n66951, n66952, n66953, n66954, n66955, n66956, n66957, n66958, n66959, 
      n66960, n66961, n66962, n66963, n66964, n66965, n66966, n66967, n66968, 
      n66969, n66970, n66971, n66972, n66973, n66974, n66975, n66976, n66977, 
      n66978, n66979, n66980, n66981, n66982, n66983, n66984, n66985, n66986, 
      n66987, n66988, n66989, n66990, n66991, n66992, n66993, n66994, n66995, 
      n66996, n66997, n66998, n66999, n67000, n67001, n67002, n67003, n67004, 
      n67005, n67006, n67007, n67008, n67009, n67010, n67011, n67012, n67013, 
      n67014, n67015, n67016, n67017, n67018, n67019, n67020, n67021, n67022, 
      n67023, n67024, n67025, n67026, n67027, n67028, n67029, n67030, n67031, 
      n67032, n67033, n67034, n67035, n67036, n67037, n67038, n67039, n67040, 
      n67041, n67042, n67043, n67044, n67045, n67046, n67047, n67048, n67049, 
      n67050, n67051, n67052, n67053, n67054, n67055, n67056, n67057, n67058, 
      n67059, n67060, n67061, n67062, n67063, n67064, n67065, n67066, n67067, 
      n67068, n67069, n67070, n67071, n67072, n67073, n67074, n67075, n67076, 
      n67077, n67078, n67079, n67080, n67081, n67082, n67083, n67084, n67085, 
      n67086, n67087, n67088, n67089, n67090, n67091, n67092, n67093, n67094, 
      n67095, n67096, n67097, n67098, n67099, n67100, n67101, n67102, n67103, 
      n67104, n67105, n67106, n67107, n67108, n67109, n67110, n67111, n67112, 
      n67113, n67114, n67115, n67116, n67117, n67118, n67119, n67120, n67121, 
      n67122, n67123, n67124, n67125, n67126, n67127, n67128, n67129, n67130, 
      n67131, n67132, n67133, n67134, n67135, n67136, n67137, n67138, n67139, 
      n67140, n67141, n67142, n67143, n67144, n67145, n67146, n67147, n67148, 
      n67149, n67150, n67151, n67152, n67153, n67154, n67155, n67156, n67157, 
      n67158, n67159, n67160, n67161, n67162, n67163, n67164, n67165, n67166, 
      n67167, n67168, n67169, n67170, n67171, n67172, n67173, n67174, n67175, 
      n67176, n67177, n67178, n67179, n67180, n67181, n67182, n67183, n67184, 
      n67185, n67186, n67187, n67188, n67189, n67190, n67191, n67192, n67193, 
      n67194, n67195, n67196, n67197, n67198, n67199, n67200, n67201, n67202, 
      n67203, n67204, n67205, n67206, n67207, n67208, n67209, n67210, n67211, 
      n67212, n67213, n67214, n67215, n67216, n67217, n67218, n67219, n67220, 
      n67221, n67222, n67223, n67224, n67225, n67226, n67227, n67228, n67229, 
      n67230, n67231, n67232, n67233, n67234, n67235, n67236, n67237, n67238, 
      n67239, n67240, n67241, n67242, n67243, n67244, n67245, n67246, n67247, 
      n67248, n67249, n67250, n67251, n67252, n67253, n67254, n67255, n67256, 
      n67257, n67258, n67259, n67260, n67261, n67262, n67263, n67264, n67265, 
      n67266, n67267, n67268, n67269, n67270, n67271, n67272, n67273, n67274, 
      n67275, n67276, n67277, n67278, n67279, n67280, n67281, n67282, n67283, 
      n67284, n67285, n67286, n67287, n67288, n67289, n67290, n67291, n67292, 
      n67293, n67294, n67295, n67296, n67297, n67298, n67299, n67300, n67301, 
      n67302, n67303, n67304, n67305, n67306, n67307, n67308, n67309, n67310, 
      n67311, n67312, n67313, n67314, n67315, n67316, n67317, n67318, n67319, 
      n67320, n67321, n67322, n67323, n67324, n67325, n67326, n67327, n67328, 
      n67329, n67330, n67331, n67332, n67333, n67334, n67335, n67336, n67337, 
      n67338, n67339, n67340, n67341, n67342, n67343, n67344, n67345, n67346, 
      n67347, n67348, n67349, n67350, n67351, n67352, n67353, n67354, n67355, 
      n67356, n67357, n67358, n67359, n67360, n67361, n67362, n67363, n67364, 
      n67365, n67366, n67367, n67368, n67369, n67370, n67371, n67372, n67373, 
      n67374, n67375, n67376, n67377, n67378, n67379, n67380, n67381, n67382, 
      n67383, n67384, n67385, n67386, n67387, n67388, n67389, n67390, n67391, 
      n67392, n67393, n67394, n67395, n67396, n67397, n67398, n67399, n67400, 
      n67401, n67402, n67403, n67404, n67405, n67406, n67407, n67408, n67409, 
      n67410, n67411, n67412, n67413, n67414, n67415, n67416, n67417, n67418, 
      n67419, n67420, n67421, n67422, n67423, n67424, n67425, n67426, n67427, 
      n67428, n67429, n67430, n67431, n67432, n67433, n67434, n67435, n67436, 
      n67437, n67438, n67439, n67440, n67441, n67442, n67443, n67444, n67445, 
      n67446, n67447, n67448, n67449, n67450, n67451, n67452, n67453, n67454, 
      n67455, n67456, n67457, n67458, n67459, n67460, n67461, n67462, n67463, 
      n67464, n67465, n67466, n67467, n67468, n67469, n67470, n67471, n67472, 
      n67473, n67474, n67475, n67476, n67477, n67478, n67479, n67480, n67481, 
      n67482, n67483, n67484, n67485, n67486, n67487, n67488, n67489, n67490, 
      n67491, n67492, n67493, n67494, n67495, n67496, n67497, n67498, n67499, 
      n67500, n67501, n67502, n67503, n67504, n67505, n67506, n67507, n67508, 
      n67509, n67510, n67511, n67512, n67513, n67514, n67515, n67516, n67517, 
      n67518, n67519, n67520, n67521, n67522, n67523, n67524, n67525, n67526, 
      n67527, n67528, n67529, n67530, n67531, n67532, n67533, n67534, n67535, 
      n67536, n67537, n67538, n67539, n67540, n67541, n67542, n67543, n67544, 
      n67545, n67546, n67547, n67548, n67549, n67550, n67551, n67552, n67553, 
      n67554, n67555, n67556, n67557, n67558, n67559, n67560, n67561, n67562, 
      n67563, n67564, n67565, n67566, n67567, n67568, n67569, n67570, n67571, 
      n67572, n67573, n67574, n67575, n67576, n67577, n67578, n67579, n67580, 
      n67581, n67582, n67583, n67584, n67585, n67586, n67587, n67588, n67589, 
      n67590, n67591, n67592, n67593, n67594, n67595, n67596, n67597, n67598, 
      n67599, n67600, n67601, n67602, n67603, n67604, n67605, n67606, n67607, 
      n67608, n67609, n67610, n67611, n67612, n67613, n67614, n67615, n67616, 
      n67617, n67618, n67619, n67620, n67621, n67622, n67623, n67624, n67625, 
      n67626, n67627, n67628, n67629, n67630, n67631, n67632, n67633, n67634, 
      n67635, n67636, n67637, n67638, n67639, n67640, n67641, n67642, n67643, 
      n67644, n67645, n67646, n67647, n67648, n67649, n67650, n67651, n67652, 
      n67653, n67654, n67655, n67656, n67657, n67658, n67659, n67660, n67661, 
      n67662, n67663, n67664, n67665, n67666, n67667, n67668, n67669, n67670, 
      n67671, n67672, n67673, n67674, n67675, n67676, n67677, n67678, n67679, 
      n67680, n67681, n67682, n67683, n67684, n67685, n67686, n67687, n67688, 
      n67689, n67690, n67691, n67692, n67693, n67694, n67695, n67696, n67697, 
      n67698, n67699, n67700, n67701, n67702, n67703, n67704, n67705, n67706, 
      n67707, n67708, n67709, n67710, n67711, n67712, n67713, n67714, n67715, 
      n67716, n67717, n67718, n67719, n67720, n67721, n67722, n67723, n67724, 
      n67725, n67726, n67727, n67728, n67729, n67730, n67731, n67732, n67733, 
      n67734, n67735, n67736, n67737, n67738, n67739, n67740, n67741, n67742, 
      n67743, n67744, n67745, n67746, n67747, n67748, n67749, n67750, n67751, 
      n67752, n67753, n67754, n67755, n67756, n67757, n67758, n67759, n67760, 
      n67761, n67762, n67763, n67764, n67765, n67766, n67767, n67768, n67769, 
      n67770, n67771, n67772, n67773, n67774, n67775, n67776, n67777, n67778, 
      n67779, n67780, n67781, n67782, n67783, n67784, n67785, n67786, n67787, 
      n67788, n67789, n67790, n67791, n67792, n67793, n67794, n67795, n67796, 
      n67797, n67798, n67799, n67800, n67801, n67802, n67803, n67804, n67805, 
      n67806, n67807, n67808, n67809, n67810, n67811, n67812, n67813, n67814, 
      n67815, n67816, n67817, n67818, n67819, n67820, n67821, n67822, n67823, 
      n67824, n67825, n67826, n67827, n67828, n67829, n67830, n67831, n67832, 
      n67833, n67834, n67835, n67836, n67837, n67838, n67839, n67840, n67841, 
      n67842, n67843, n67844, n67845, n67846, n67847, n67848, n67849, n67850, 
      n67851, n67852, n67853, n67854, n67855, n67856, n67857, n67858, n67859, 
      n67860, n67861, n67862, n67863, n67864, n67865, n67866, n67867, n67868, 
      n67869, n67870, n67871, n67872, n67873, n67874, n67875, n67876, n67877, 
      n67878, n67879, n67880, n67881, n67882, n67883, n67884, n67885, n67886, 
      n67887, n67888, n67889, n67890, n67891, n67892, n67893, n67894, n67895, 
      n67896, n67897, n67898, n67899, n67900, n67901, n67902, n67903, n67904, 
      n67905, n67906, n67907, n67908, n67909, n67910, n67911, n67912, n67913, 
      n67914, n67915, n67916, n67917, n67918, n67919, n67920, n67921, n67922, 
      n67923, n67924, n67925, n67926, n67927, n67928, n67929, n67930, n67931, 
      n67932, n67933, n67934, n67935, n67936, n67937, n67938, n67939, n67940, 
      n67941, n67942, n67943, n67944, n67945, n67946, n67947, n67948, n67949, 
      n67950, n67951, n67952, n67953, n67954, n67955, n67956, n67957, n67958, 
      n67959, n67960, n67961, n67962, n67963, n67964, n67965, n67966, n67967, 
      n67968, n67969, n67970, n67971, n67972, n67973, n67974, n67975, n67976, 
      n67977, n67978, n67979, n67980, n67981, n67982, n67983, n67984, n67985, 
      n67986, n67987, n67988, n67989, n67990, n67991, n67992, n67993, n67994, 
      n67995, n67996, n67997, n67998, n67999, n68000, n68001, n68002, n68003, 
      n68004, n68005, n68006, n68007, n68008, n68009, n68010, n68011, n68012, 
      n68013, n68014, n68015, n68016, n68017, n68018, n68019, n68020, n68021, 
      n68022, n68023, n68024, n68025, n68026, n68027, n68028, n68029, n68030, 
      n68031, n68032, n68033, n68034, n68035, n68036, n68037, n68038, n68039, 
      n68040, n68041, n68042, n68043, n68044, n68045, n68046, n68047, n68048, 
      n68049, n68050, n68051, n68052, n68053, n68054, n68055, n68056, n68057, 
      n68058, n68059, n68060, n68061, n68062, n68063, n68064, n68065, n68066, 
      n68067, n68068, n68069, n68070, n68071, n68072, n68073, n68074, n68075, 
      n68076, n68077, n68078, n68079, n68080, n68081, n68082, n68083, n68084, 
      n68085, n68086, n68087, n68088, n68089, n68090, n68091, n68092, n68093, 
      n68094, n68095, n68096, n68097, n68098, n68099, n68100, n68101, n68102, 
      n68103, n68104, n68105, n68106, n68107, n68108, n68109, n68110, n68111, 
      n68112, n68113, n68114, n68115, n68116, n68117, n68118, n68119, n68120, 
      n68121, n68122, n68123, n68124, n68125, n68126, n68127, n68128, n68129, 
      n68130, n68131, n68132, n68133, n68134, n68135, n68136, n68137, n68138, 
      n68139, n68140, n68141, n68142, n68143, n68144, n68145, n68146, n68147, 
      n68148, n68149, n68150, n68151, n68152, n68153, n68154, n68155, n68156, 
      n68157, n68158, n68159, n68160, n68161, n68162, n68163, n68164, n68165, 
      n68166, n68167, n68168, n68169, n68170, n68171, n68172, n68173, n68174, 
      n68175, n68176, n68177, n68178, n68179, n68180, n68181, n68182, n68183, 
      n68184, n68185, n68186, n68187, n68188, n68189, n68190, n68191, n68192, 
      n68193, n68194, n68195, n68196, n68197, n68198, n68199, n68200, n68201, 
      n68202, n68203, n68204, n68205, n68206, n68207, n68208, n68209, n68210, 
      n68211, n68212, n68213, n68214, n68215, n68216, n68217, n68218, n68219, 
      n68220, n68221, n68222, n68223, n68224, n68225, n68226, n68227, n68228, 
      n68229, n68230, n68231, n68232, n68233, n68234, n68235, n68236, n68237, 
      n68238, n68239, n68240, n68241, n68242, n68243, n68244, n68245, n68246, 
      n68247, n68248, n68249, n68250, n68251, n68252, n68253, n68254, n68255, 
      n68256, n68257, n68258, n68259, n68260, n68261, n68262 : std_logic;

begin
   OUT1 <= ( OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, 
      OUT1_59_port, OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, 
      OUT1_54_port, OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, 
      OUT1_49_port, OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, 
      OUT1_44_port, OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, 
      OUT1_39_port, OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, 
      OUT1_34_port, OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, 
      OUT1_29_port, OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, 
      OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, 
      OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, 
      OUT1_14_port, OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, 
      OUT1_9_port, OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, 
      OUT1_4_port, OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_63_port, OUT2_62_port, OUT2_61_port, OUT2_60_port, 
      OUT2_59_port, OUT2_58_port, OUT2_57_port, OUT2_56_port, OUT2_55_port, 
      OUT2_54_port, OUT2_53_port, OUT2_52_port, OUT2_51_port, OUT2_50_port, 
      OUT2_49_port, OUT2_48_port, OUT2_47_port, OUT2_46_port, OUT2_45_port, 
      OUT2_44_port, OUT2_43_port, OUT2_42_port, OUT2_41_port, OUT2_40_port, 
      OUT2_39_port, OUT2_38_port, OUT2_37_port, OUT2_36_port, OUT2_35_port, 
      OUT2_34_port, OUT2_33_port, OUT2_32_port, OUT2_31_port, OUT2_30_port, 
      OUT2_29_port, OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, 
      OUT2_24_port, OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, 
      OUT2_19_port, OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, 
      OUT2_14_port, OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, 
      OUT2_9_port, OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, 
      OUT2_4_port, OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   OUT1_reg_59_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => OUT1_59_port
                           , QN => n4282);
   OUT1_reg_58_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => OUT1_58_port
                           , QN => n4281);
   OUT1_reg_57_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => OUT1_57_port
                           , QN => n4280);
   OUT1_reg_56_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => OUT1_56_port
                           , QN => n4279);
   OUT1_reg_55_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => OUT1_55_port
                           , QN => n4278);
   OUT1_reg_54_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => OUT1_54_port
                           , QN => n4277);
   OUT1_reg_53_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => OUT1_53_port
                           , QN => n4276);
   OUT1_reg_52_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => OUT1_52_port
                           , QN => n4275);
   OUT1_reg_51_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => OUT1_51_port
                           , QN => n4274);
   OUT1_reg_50_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => OUT1_50_port
                           , QN => n4273);
   OUT1_reg_49_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => OUT1_49_port
                           , QN => n4272);
   OUT1_reg_48_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => OUT1_48_port
                           , QN => n4271);
   OUT1_reg_47_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => OUT1_47_port
                           , QN => n4270);
   OUT1_reg_46_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => OUT1_46_port
                           , QN => n4269);
   OUT1_reg_45_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => OUT1_45_port
                           , QN => n4268);
   OUT1_reg_44_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => OUT1_44_port
                           , QN => n4267);
   OUT1_reg_43_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => OUT1_43_port
                           , QN => n4266);
   OUT1_reg_42_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => OUT1_42_port
                           , QN => n4265);
   OUT1_reg_41_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => OUT1_41_port
                           , QN => n4264);
   OUT1_reg_40_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => OUT1_40_port
                           , QN => n4263);
   OUT1_reg_39_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => OUT1_39_port
                           , QN => n4262);
   OUT1_reg_38_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => OUT1_38_port
                           , QN => n4261);
   OUT1_reg_37_inst : DFF_X1 port map( D => n5449, CK => CLK, Q => OUT1_37_port
                           , QN => n4260);
   OUT1_reg_36_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => OUT1_36_port
                           , QN => n4259);
   OUT1_reg_35_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => OUT1_35_port
                           , QN => n4258);
   OUT1_reg_34_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => OUT1_34_port
                           , QN => n4257);
   OUT1_reg_33_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => OUT1_33_port
                           , QN => n4256);
   OUT1_reg_32_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => OUT1_32_port
                           , QN => n4255);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => OUT1_31_port
                           , QN => n4254);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => OUT1_30_port
                           , QN => n4253);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => OUT1_29_port
                           , QN => n4252);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => OUT1_28_port
                           , QN => n4251);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => OUT1_27_port
                           , QN => n4250);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => OUT1_26_port
                           , QN => n4249);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => OUT1_25_port
                           , QN => n4248);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => OUT1_24_port
                           , QN => n4247);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => OUT1_23_port
                           , QN => n4246);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => OUT1_22_port
                           , QN => n4245);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5417, CK => CLK, Q => OUT1_21_port
                           , QN => n4244);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5415, CK => CLK, Q => OUT1_20_port
                           , QN => n4243);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => OUT1_19_port
                           , QN => n4242);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => OUT1_18_port
                           , QN => n4241);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => OUT1_17_port
                           , QN => n4240);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => OUT1_16_port
                           , QN => n4239);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => OUT1_15_port
                           , QN => n4238);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => OUT1_14_port
                           , QN => n4237);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => OUT1_13_port
                           , QN => n4236);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => OUT1_12_port
                           , QN => n4235);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => OUT1_11_port
                           , QN => n4234);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => OUT1_10_port
                           , QN => n4233);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => OUT1_9_port, 
                           QN => n4232);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => OUT1_8_port, 
                           QN => n4231);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => OUT1_7_port, 
                           QN => n4230);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => OUT1_6_port, 
                           QN => n4229);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => OUT1_5_port, 
                           QN => n4228);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => OUT1_4_port, 
                           QN => n4227);
   OUT1_reg_3_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => OUT1_3_port, 
                           QN => n4226);
   OUT1_reg_2_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => OUT1_2_port, 
                           QN => n4225);
   OUT1_reg_1_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => OUT1_1_port, 
                           QN => n4224);
   OUT1_reg_0_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => OUT1_0_port, 
                           QN => n4223);
   OUT2_reg_61_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => OUT2_61_port
                           , QN => n4220);
   OUT2_reg_60_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => OUT2_60_port
                           , QN => n4219);
   OUT2_reg_59_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => OUT2_59_port
                           , QN => n4218);
   OUT2_reg_58_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => OUT2_58_port
                           , QN => n4217);
   OUT2_reg_57_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => OUT2_57_port
                           , QN => n4216);
   OUT2_reg_56_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => OUT2_56_port
                           , QN => n4215);
   OUT2_reg_55_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => OUT2_55_port
                           , QN => n4214);
   OUT2_reg_54_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => OUT2_54_port
                           , QN => n4213);
   OUT2_reg_53_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => OUT2_53_port
                           , QN => n4212);
   OUT2_reg_52_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => OUT2_52_port
                           , QN => n4211);
   OUT2_reg_51_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => OUT2_51_port
                           , QN => n4210);
   OUT2_reg_50_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => OUT2_50_port
                           , QN => n4209);
   OUT2_reg_49_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => OUT2_49_port
                           , QN => n4208);
   OUT2_reg_48_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => OUT2_48_port
                           , QN => n4207);
   OUT2_reg_47_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => OUT2_47_port
                           , QN => n4206);
   OUT2_reg_46_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => OUT2_46_port
                           , QN => n4205);
   OUT2_reg_45_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => OUT2_45_port
                           , QN => n4204);
   OUT2_reg_44_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => OUT2_44_port
                           , QN => n4203);
   OUT2_reg_43_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => OUT2_43_port
                           , QN => n4202);
   OUT2_reg_42_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => OUT2_42_port
                           , QN => n4201);
   OUT2_reg_41_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => OUT2_41_port
                           , QN => n4200);
   OUT2_reg_40_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => OUT2_40_port
                           , QN => n4199);
   OUT2_reg_39_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => OUT2_39_port
                           , QN => n4198);
   OUT2_reg_38_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => OUT2_38_port
                           , QN => n4197);
   OUT2_reg_37_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => OUT2_37_port
                           , QN => n4196);
   OUT2_reg_36_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => OUT2_36_port
                           , QN => n4195);
   OUT2_reg_35_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => OUT2_35_port
                           , QN => n4194);
   OUT2_reg_34_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => OUT2_34_port
                           , QN => n4193);
   OUT2_reg_33_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => OUT2_33_port
                           , QN => n4192);
   OUT2_reg_32_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => OUT2_32_port
                           , QN => n4191);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => OUT2_31_port
                           , QN => n4190);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5341, CK => CLK, Q => OUT2_30_port
                           , QN => n4189);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5340, CK => CLK, Q => OUT2_29_port
                           , QN => n4188);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5339, CK => CLK, Q => OUT2_28_port
                           , QN => n4187);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5338, CK => CLK, Q => OUT2_27_port
                           , QN => n4186);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5337, CK => CLK, Q => OUT2_26_port
                           , QN => n4185);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5336, CK => CLK, Q => OUT2_25_port
                           , QN => n4184);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5335, CK => CLK, Q => OUT2_24_port
                           , QN => n4183);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5334, CK => CLK, Q => OUT2_23_port
                           , QN => n4182);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5333, CK => CLK, Q => OUT2_22_port
                           , QN => n4181);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5332, CK => CLK, Q => OUT2_21_port
                           , QN => n4180);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5331, CK => CLK, Q => OUT2_20_port
                           , QN => n4179);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5330, CK => CLK, Q => OUT2_19_port
                           , QN => n4178);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5329, CK => CLK, Q => OUT2_18_port
                           , QN => n4177);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5328, CK => CLK, Q => OUT2_17_port
                           , QN => n4176);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5327, CK => CLK, Q => OUT2_16_port
                           , QN => n4175);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5326, CK => CLK, Q => OUT2_15_port
                           , QN => n4174);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5325, CK => CLK, Q => OUT2_14_port
                           , QN => n4173);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5324, CK => CLK, Q => OUT2_13_port
                           , QN => n4172);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5323, CK => CLK, Q => OUT2_12_port
                           , QN => n4171);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5322, CK => CLK, Q => OUT2_11_port
                           , QN => n4170);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5321, CK => CLK, Q => OUT2_10_port
                           , QN => n4169);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5320, CK => CLK, Q => OUT2_9_port, 
                           QN => n4168);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5319, CK => CLK, Q => OUT2_8_port, 
                           QN => n4167);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5318, CK => CLK, Q => OUT2_7_port, 
                           QN => n4166);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5317, CK => CLK, Q => OUT2_6_port, 
                           QN => n4165);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5316, CK => CLK, Q => OUT2_5_port, 
                           QN => n4164);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5315, CK => CLK, Q => OUT2_4_port, 
                           QN => n4163);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5314, CK => CLK, Q => OUT2_3_port, 
                           QN => n4162);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5313, CK => CLK, Q => OUT2_2_port, 
                           QN => n4161);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5312, CK => CLK, Q => OUT2_1_port, 
                           QN => n4160);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5311, CK => CLK, Q => OUT2_0_port, 
                           QN => n4159);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n58960, QN => n8497);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n59026, QN => n8481);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n59024, QN => n8465);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n59022, QN => n8449);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n42006, QN => n49483);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n42005, QN => n49482);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n42004, QN => n49481);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n42003, QN => n49480);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n56611, QN => n8433);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n56635, QN => n8417);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n56659, QN => n8401);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n56683, QN => n8385);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n56707, QN => n8369);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n56731, QN => n8353);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n56755, QN => n8337);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n56779, QN => n8321);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n56803, QN => n8305);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n56827, QN => n8289);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n56851, QN => n8273);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n56875, QN => n8257);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n56899, QN => n8241);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n56923, QN => n8225);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n56947, QN => n8209);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n56971, QN => n8193);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n56995, QN => n8177);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n57019, QN => n8161);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n57043, QN => n8145);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n57067, QN => n8129);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n57091, QN => n8113);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n57115, QN => n8097);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n57139, QN => n8081);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n57163, QN => n8065);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n57187, QN => n8049);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n57211, QN => n8033);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n57235, QN => n8017);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n57259, QN => n8001);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n57283, QN => n7985);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n57307, QN => n7969);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n57331, QN => n7953);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n57355, QN => n7937);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n57379, QN => n7921);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n57403, QN => n7905);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n57427, QN => n7889);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n57451, QN => n7873);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n57475, QN => n7857);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n57499, QN => n7841);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n57523, QN => n7825);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n57547, QN => n7809);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n57571, QN => n7793);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n57595, QN => n7777);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n57619, QN => n7761);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n57643, QN => n7745);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n57667, QN => n7729);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n57691, QN => n7713);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n57715, QN => n7697);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n57739, QN => n7681);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n57763, QN => n7665);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n57787, QN => n7649);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n57811, QN => n7633);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n57835, QN => n7617);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n57859, QN => n7601);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n57883, QN => n7585);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n57907, QN => n7569);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n57931, QN => n7553);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n57955, QN => n7537);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n57979, QN => n7521);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n58003, QN => n7505);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n58041, QN => n7489);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n41818, QN => n49479);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n41817, QN => n49478);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n41816, QN => n49477);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n41815, QN => n49476);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n41814, QN => n49475);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n41813, QN => n49474);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n41812, QN => n49473);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n41811, QN => n49472);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n41810, QN => n49471);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n41809, QN => n49470);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n41808, QN => n49469);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n41807, QN => n49468);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n41806, QN => n49467);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n41805, QN => n49466);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n41804, QN => n49465);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n41803, QN => n49464);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n41802, QN => n49463);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n41801, QN => n49462);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n41800, QN => n49461);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n41799, QN => n49460);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n41798, QN => n49459);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n41797, QN => n49458);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n41796, QN => n49457);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n41795, QN => n49456);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n41794, QN => n49455);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n41793, QN => n49454);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n41792, QN => n49453);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n41791, QN => n49452);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n41790, QN => n49451);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n41789, QN => n49450);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n41788, QN => n49449);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n41787, QN => n49448);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n41786, QN => n49447);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n41785, QN => n49446);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n41784, QN => n49445);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n41783, QN => n49444);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n41782, QN => n49443);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n41781, QN => n49442);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n41780, QN => n49441);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n41779, QN => n49440);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n41778, QN => n49439);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n41777, QN => n49438);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n41776, QN => n49437);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n41775, QN => n49436);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n41774, QN => n49435);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n41773, QN => n49434);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n41772, QN => n49433);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n41771, QN => n49432);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n41770, QN => n49431);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n41769, QN => n49430);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n41768, QN => n49429);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n41767, QN => n49428);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n41766, QN => n49427);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n41765, QN => n49426);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n41764, QN => n49425);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n41763, QN => n49424);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n41762, QN => n49423);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n41761, QN => n49422);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n41760, QN => n49421);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n41759, QN => n49420);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n66498, QN => n8509);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n66497, QN => n8493);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n66496, QN => n8477);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n66495, QN => n8461);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => 
                           n66550, QN => n49228);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n66501, QN => n49231);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n66500, QN => n49230);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n66499, QN => n49229);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n66513, QN => n49291);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n66512, QN => n49290);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n66511, QN => n49289);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n66510, QN => n49288);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n66509, QN => n49287);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n66508, QN => n49286);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n66507, QN => n49285);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n66506, QN => n49284);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n66505, QN => n49283);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n66504, QN => n49282);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n66503, QN => n49281);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n66502, QN => n49280);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n66549, QN => n49279);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n66548, QN => n49278);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n66547, QN => n49277);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n66546, QN => n49276);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n66545, QN => n49275);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n66544, QN => n49274);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n66543, QN => n49273);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n66542, QN => n49272);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n66541, QN => n49271);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n66540, QN => n49270);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n66539, QN => n49269);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n66538, QN => n49268);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n66537, QN => n49267);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n66536, QN => n49266);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n66535, QN => n49265);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n66534, QN => n49264);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n66533, QN => n49263);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n66532, QN => n49262);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n66531, QN => n49261);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n66530, QN => n49260);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n66529, QN => n49259);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n66528, QN => n49258);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n66527, QN => n49257);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n66526, QN => n49256);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n66525, QN => n49255);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n66524, QN => n49254);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n66523, QN => n49253);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n66522, QN => n49252);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n66521, QN => n49251);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n66520, QN => n49250);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n66519, QN => n49249);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n66518, QN => n49248);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n66517, QN => n49247);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n66516, QN => n49246);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n66515, QN => n49245);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n66514, QN => n49244);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n64855, QN => n49243);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n64875, QN => n49242);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n64895, QN => n49241);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => 
                           n64915, QN => n49240);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => 
                           n64935, QN => n49239);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => 
                           n64955, QN => n49238);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => 
                           n64975, QN => n49237);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n64995, QN => n49236);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n65015, QN => n49235);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n65035, QN => n49234);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n65055, QN => n49233);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n65084, QN => n49232);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => 
                           n50647, QN => n54606);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => 
                           n50646, QN => n54608);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n50645, QN => n54609);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => 
                           n50644, QN => n54610);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => 
                           n50579, QN => n54184);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => 
                           n50578, QN => n54185);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => 
                           n50577, QN => n54186);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n50707, QN => n54611);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => 
                           n50706, QN => n54612);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n50705, QN => n54613);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => 
                           n50704, QN => n54614);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n50703, QN => n54615);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => 
                           n50702, QN => n54616);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n50701, QN => n54617);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => 
                           n50700, QN => n54618);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n50699, QN => n54619);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => 
                           n50698, QN => n54620);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n50697, QN => n54621);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => 
                           n50696, QN => n54622);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n50695, QN => n54623);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => 
                           n50694, QN => n54624);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n50693, QN => n54625);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => 
                           n50692, QN => n54626);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n50691, QN => n54627);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => 
                           n50690, QN => n54628);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n50689, QN => n54629);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => 
                           n50688, QN => n54630);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n50687, QN => n54631);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => 
                           n50686, QN => n54632);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n50685, QN => n54633);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => 
                           n50684, QN => n54634);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n50683, QN => n54635);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => 
                           n50682, QN => n54636);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n50681, QN => n54637);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => 
                           n50680, QN => n54638);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n50679, QN => n54639);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => 
                           n50678, QN => n54640);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n50677, QN => n54641);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => 
                           n50676, QN => n54642);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n50675, QN => n54643);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => 
                           n50674, QN => n54644);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n50673, QN => n54645);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => 
                           n50672, QN => n54646);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n50671, QN => n54647);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => 
                           n50670, QN => n54648);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n50669, QN => n54649);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => 
                           n50668, QN => n54650);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n50667, QN => n54651);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => 
                           n50666, QN => n54652);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n50665, QN => n54653);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => 
                           n50664, QN => n54654);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n50663, QN => n54655);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => 
                           n50662, QN => n54656);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n50661, QN => n54657);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => 
                           n50660, QN => n54658);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n50659, QN => n54659);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => 
                           n50658, QN => n54660);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => 
                           n50657, QN => n54661);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => 
                           n50656, QN => n54662);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => 
                           n50655, QN => n54663);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => 
                           n50654, QN => n54664);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => 
                           n50653, QN => n54665);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => 
                           n50652, QN => n54666);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => 
                           n50651, QN => n54667);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => 
                           n50650, QN => n54668);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => 
                           n50649, QN => n54669);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => 
                           n50648, QN => n54670);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => 
                           n50576, QN => n54187);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => 
                           n50575, QN => n54188);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => 
                           n50574, QN => n54189);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => 
                           n50573, QN => n54190);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => 
                           n50572, QN => n54191);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => 
                           n50571, QN => n54192);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => 
                           n50570, QN => n54193);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => 
                           n50569, QN => n54194);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => 
                           n50568, QN => n54195);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => 
                           n50567, QN => n54196);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => 
                           n50566, QN => n54197);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => 
                           n50565, QN => n54198);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => 
                           n50564, QN => n54199);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => 
                           n50563, QN => n54200);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => 
                           n50562, QN => n54201);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => 
                           n50561, QN => n54202);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => 
                           n50560, QN => n54203);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => 
                           n50559, QN => n54204);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => 
                           n50558, QN => n54205);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => 
                           n50557, QN => n54206);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => 
                           n50556, QN => n54207);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => 
                           n50555, QN => n54208);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => 
                           n50554, QN => n54209);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => 
                           n50553, QN => n54210);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => 
                           n50552, QN => n54211);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => 
                           n50551, QN => n54212);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => 
                           n50550, QN => n54213);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => 
                           n50549, QN => n54214);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => 
                           n50548, QN => n54215);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => 
                           n50547, QN => n54216);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => 
                           n50546, QN => n54217);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => 
                           n50545, QN => n54218);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => 
                           n50544, QN => n54219);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => 
                           n50543, QN => n54220);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => 
                           n50542, QN => n54221);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => 
                           n50541, QN => n54222);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => 
                           n50540, QN => n54223);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => 
                           n50539, QN => n54224);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => 
                           n50538, QN => n54225);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => 
                           n50537, QN => n54226);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => 
                           n50536, QN => n54227);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => 
                           n50535, QN => n54228);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => 
                           n50534, QN => n54229);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => 
                           n50533, QN => n54230);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => 
                           n50532, QN => n54231);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => 
                           n50531, QN => n54232);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => 
                           n50530, QN => n54233);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => 
                           n50529, QN => n54234);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => 
                           n50528, QN => n54235);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => 
                           n50527, QN => n54236);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => 
                           n50526, QN => n54237);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => 
                           n50525, QN => n54238);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => 
                           n50524, QN => n54239);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => 
                           n50523, QN => n54240);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => 
                           n50522, QN => n54241);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => 
                           n50521, QN => n54242);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => 
                           n50520, QN => n54243);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => 
                           n50519, QN => n54244);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => 
                           n50518, QN => n54245);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => 
                           n50517, QN => n54246);
   OUT2_reg_63_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => OUT2_63_port
                           , QN => n59028);
   OUT2_reg_62_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => OUT2_62_port
                           , QN => n59027);
   U45435 : NOR3_X2 port map( A1 => n67434, A2 => ADD_RD2(2), A3 => n66301, ZN 
                           => n66283);
   U45452 : NAND3_X1 port map( A1 => n62490, A2 => n62491, A3 => n62492, ZN => 
                           n62088);
   U45453 : NAND3_X1 port map( A1 => n62492, A2 => n62491, A3 => ADD_WR(0), ZN 
                           => n62156);
   U45454 : NAND3_X1 port map( A1 => n62492, A2 => n62490, A3 => ADD_WR(3), ZN 
                           => n62625);
   U45455 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n62492, A3 => ADD_WR(3), 
                           ZN => n62692);
   U45456 : NAND3_X1 port map( A1 => n62490, A2 => n62491, A3 => n63295, ZN => 
                           n63025);
   U45457 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n62491, A3 => n63295, ZN 
                           => n63092);
   U45458 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n62490, A3 => n63295, ZN 
                           => n63428);
   U45459 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(0), A3 => n63295, 
                           ZN => n63495);
   U45461 : NAND3_X1 port map( A1 => ENABLE, A2 => n68057, A3 => RD2, ZN => 
                           n65112);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => 
                           n58378, QN => n63765);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => 
                           n58377, QN => n63820);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => 
                           n58376, QN => n63841);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => 
                           n58375, QN => n63862);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n5566, CK => CLK, Q => 
                           n66308, QN => n63699);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n5565, CK => CLK, Q => 
                           n66307, QN => n63701);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n5564, CK => CLK, Q => 
                           n66306, QN => n63702);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n5563, CK => CLK, Q => 
                           n66305, QN => n63703);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => 
                           n67259, QN => n63633);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => 
                           n67258, QN => n63635);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => 
                           n67257, QN => n63636);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => 
                           n67256, QN => n63637);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => 
                           n67255, QN => n63567);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n67254, QN => n63569);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => 
                           n67253, QN => n63570);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n67252, QN => n63571);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => 
                           n67251, QN => n63501);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => 
                           n67250, QN => n63503);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => 
                           n67249, QN => n63504);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n67248, QN => n63505);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => 
                           n8959, QN => n63430);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => 
                           n8961, QN => n63432);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n8963, QN => n63433);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => 
                           n8965, QN => n63434);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => 
                           n67247, QN => n63297);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n67246, QN => n63299);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n67245, QN => n63300);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n67244, QN => n63301);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n67243, QN => n63096);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n67242, QN => n63098);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n67241, QN => n63099);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n67240, QN => n63100);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => 
                           n67239, QN => n63363);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n67238, QN => n63365);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n67237, QN => n63366);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n67236, QN => n63367);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => 
                           n58234, QN => n63027);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n58233, QN => n63029);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n58232, QN => n63030);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n58231, QN => n63031);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => 
                           n58370, QN => n62960);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n58369, QN => n62962);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n58368, QN => n62963);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n58367, QN => n62964);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n58718, QN => n63230);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n58717, QN => n63232);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n58716, QN => n63233);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n58715, QN => n63234);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => 
                           n58301, QN => n63162);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n58299, QN => n63164);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n58297, QN => n63165);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n58295, QN => n63166);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => 
                           n67235, QN => n62694);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7486, CK => CLK, Q => 
                           n56490, QN => n61958);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7485, CK => CLK, Q => 
                           n56531, QN => n61961);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7484, CK => CLK, Q => 
                           n56555, QN => n61963);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7483, CK => CLK, Q => 
                           n56579, QN => n61965);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => 
                           n58050, QN => n62494);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => 
                           n58049, QN => n62496);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n58048, QN => n62497);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n58047, QN => n62498);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => 
                           n58782, QN => n62358);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => 
                           n58781, QN => n62360);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => 
                           n58780, QN => n62361);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => 
                           n58779, QN => n62362);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => 
                           n67234, QN => n62225);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => 
                           n67233, QN => n62227);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => 
                           n67232, QN => n62228);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => 
                           n67231, QN => n62229);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => 
                           n67230, QN => n62158);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => 
                           n67229, QN => n62160);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => 
                           n67228, QN => n62161);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => 
                           n67227, QN => n62162);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => 
                           n58438, QN => n63883);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => 
                           n58437, QN => n63903);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => 
                           n58436, QN => n63923);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => 
                           n58435, QN => n63943);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => 
                           n58434, QN => n63963);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => 
                           n58433, QN => n63983);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => 
                           n58432, QN => n64003);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => 
                           n58431, QN => n64023);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => 
                           n58430, QN => n64043);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => 
                           n58429, QN => n64063);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => 
                           n58428, QN => n64083);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => 
                           n58427, QN => n64103);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => 
                           n58426, QN => n64123);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => 
                           n58425, QN => n64143);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => 
                           n58424, QN => n64163);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => 
                           n58423, QN => n64183);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => 
                           n58422, QN => n64203);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => 
                           n58421, QN => n64223);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => 
                           n58420, QN => n64243);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => 
                           n58419, QN => n64263);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => 
                           n58418, QN => n64283);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => 
                           n58417, QN => n64303);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => 
                           n58416, QN => n64323);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => 
                           n58415, QN => n64343);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => 
                           n58414, QN => n64363);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => 
                           n58413, QN => n64383);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => 
                           n58412, QN => n64403);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => 
                           n58411, QN => n64423);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => 
                           n58410, QN => n64443);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => 
                           n58409, QN => n64463);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => 
                           n58408, QN => n64483);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => 
                           n58407, QN => n64503);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => 
                           n58406, QN => n64523);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => 
                           n58405, QN => n64543);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => 
                           n58404, QN => n64563);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => 
                           n58403, QN => n64583);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => 
                           n58402, QN => n64603);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => 
                           n58401, QN => n64623);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => 
                           n58400, QN => n64643);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => 
                           n58399, QN => n64663);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => 
                           n58398, QN => n64683);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => 
                           n58397, QN => n64703);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => 
                           n58396, QN => n64723);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => 
                           n58395, QN => n64743);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => 
                           n58394, QN => n64763);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => 
                           n58393, QN => n64783);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => 
                           n58392, QN => n64803);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => 
                           n58391, QN => n64823);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => 
                           n58390, QN => n64843);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => 
                           n58389, QN => n64863);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => 
                           n58388, QN => n64883);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => 
                           n58387, QN => n64903);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => 
                           n58386, QN => n64923);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => 
                           n58385, QN => n64943);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => 
                           n58384, QN => n64963);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => 
                           n58383, QN => n64983);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => 
                           n58382, QN => n65003);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => 
                           n58381, QN => n65023);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => 
                           n58380, QN => n65043);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => 
                           n58379, QN => n65063);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => 
                           n67226, QN => n62424);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => 
                           n67225, QN => n62426);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n67224, QN => n62427);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n67223, QN => n62428);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => 
                           n59092, QN => n62291);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => 
                           n59091, QN => n62293);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => 
                           n59090, QN => n62294);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => 
                           n59089, QN => n62295);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n7422, CK => CLK, Q => 
                           n67222, QN => n62091);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n7421, CK => CLK, Q => 
                           n67221, QN => n62093);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => 
                           n67220, QN => n62094);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => 
                           n67219, QN => n62095);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => 
                           n58303, QN => n62560);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n58306, QN => n62562);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n58305, QN => n62563);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n58304, QN => n62564);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => 
                           n58783, QN => n62827);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n58786, QN => n62829);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n58785, QN => n62830);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n58784, QN => n62831);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n5562, CK => CLK, Q => 
                           n66372, QN => n63704);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n5561, CK => CLK, Q => 
                           n66371, QN => n63705);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n5560, CK => CLK, Q => 
                           n66370, QN => n63706);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n5559, CK => CLK, Q => 
                           n66369, QN => n63707);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n5558, CK => CLK, Q => 
                           n66368, QN => n63708);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n5557, CK => CLK, Q => 
                           n66367, QN => n63709);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n5556, CK => CLK, Q => 
                           n66366, QN => n63710);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n5555, CK => CLK, Q => 
                           n66365, QN => n63711);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n5554, CK => CLK, Q => 
                           n66364, QN => n63712);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n5553, CK => CLK, Q => 
                           n66363, QN => n63713);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n5552, CK => CLK, Q => 
                           n66362, QN => n63714);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n5551, CK => CLK, Q => 
                           n66361, QN => n63715);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n5550, CK => CLK, Q => 
                           n66360, QN => n63716);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n5549, CK => CLK, Q => 
                           n66359, QN => n63717);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n5548, CK => CLK, Q => 
                           n66358, QN => n63718);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n5547, CK => CLK, Q => 
                           n66357, QN => n63719);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n5546, CK => CLK, Q => 
                           n66356, QN => n63720);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n5545, CK => CLK, Q => 
                           n66355, QN => n63721);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n5544, CK => CLK, Q => 
                           n66354, QN => n63722);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n5543, CK => CLK, Q => 
                           n66353, QN => n63723);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n5542, CK => CLK, Q => 
                           n66352, QN => n63724);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n5541, CK => CLK, Q => 
                           n66351, QN => n63725);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n5540, CK => CLK, Q => 
                           n66350, QN => n63726);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n5539, CK => CLK, Q => 
                           n66349, QN => n63727);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n5538, CK => CLK, Q => 
                           n66348, QN => n63728);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n5537, CK => CLK, Q => 
                           n66347, QN => n63729);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n5536, CK => CLK, Q => 
                           n66346, QN => n63730);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n5535, CK => CLK, Q => 
                           n66345, QN => n63731);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n5534, CK => CLK, Q => 
                           n66344, QN => n63732);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n5533, CK => CLK, Q => 
                           n66343, QN => n63733);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n5532, CK => CLK, Q => 
                           n66342, QN => n63734);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n5531, CK => CLK, Q => 
                           n66341, QN => n63735);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n5530, CK => CLK, Q => 
                           n66340, QN => n63736);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n5529, CK => CLK, Q => 
                           n66339, QN => n63737);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n5528, CK => CLK, Q => 
                           n66338, QN => n63738);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n5527, CK => CLK, Q => 
                           n66337, QN => n63739);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n5526, CK => CLK, Q => 
                           n66336, QN => n63740);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n5525, CK => CLK, Q => 
                           n66335, QN => n63741);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n5524, CK => CLK, Q => 
                           n66334, QN => n63742);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n5523, CK => CLK, Q => 
                           n66333, QN => n63743);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n5522, CK => CLK, Q => 
                           n66332, QN => n63744);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n5521, CK => CLK, Q => 
                           n66331, QN => n63745);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n5520, CK => CLK, Q => 
                           n66330, QN => n63746);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n5519, CK => CLK, Q => 
                           n66329, QN => n63747);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n5518, CK => CLK, Q => 
                           n66328, QN => n63748);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n5517, CK => CLK, Q => 
                           n66327, QN => n63749);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n5516, CK => CLK, Q => 
                           n66326, QN => n63750);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n5515, CK => CLK, Q => 
                           n66325, QN => n63751);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n5514, CK => CLK, Q => 
                           n66324, QN => n63752);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => 
                           n66323, QN => n63753);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => 
                           n66322, QN => n63754);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => 
                           n66321, QN => n63755);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => 
                           n66320, QN => n63756);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => 
                           n66319, QN => n63757);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => 
                           n66318, QN => n63758);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => 
                           n66317, QN => n63759);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => 
                           n66316, QN => n63760);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => 
                           n66315, QN => n63761);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => 
                           n66314, QN => n63762);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => 
                           n66313, QN => n63763);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => 
                           n67218, QN => n63638);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => 
                           n67217, QN => n63639);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => 
                           n67216, QN => n63640);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => 
                           n67215, QN => n63641);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => 
                           n67214, QN => n63642);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => 
                           n67213, QN => n63643);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => 
                           n67212, QN => n63644);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => 
                           n67211, QN => n63645);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => 
                           n67210, QN => n63646);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => 
                           n67209, QN => n63647);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => 
                           n67208, QN => n63648);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => 
                           n67207, QN => n63649);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => 
                           n67206, QN => n63650);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => 
                           n67205, QN => n63651);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => 
                           n67204, QN => n63652);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => 
                           n67203, QN => n63653);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => 
                           n67202, QN => n63654);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => 
                           n67201, QN => n63655);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n5608, CK => CLK, Q => 
                           n67200, QN => n63656);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n5607, CK => CLK, Q => 
                           n67199, QN => n63657);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n5606, CK => CLK, Q => 
                           n67198, QN => n63658);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n5605, CK => CLK, Q => 
                           n67197, QN => n63659);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n5604, CK => CLK, Q => 
                           n67196, QN => n63660);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n5603, CK => CLK, Q => 
                           n67195, QN => n63661);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n5602, CK => CLK, Q => 
                           n67194, QN => n63662);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n5601, CK => CLK, Q => 
                           n67193, QN => n63663);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n5600, CK => CLK, Q => 
                           n67192, QN => n63664);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n5599, CK => CLK, Q => 
                           n67191, QN => n63665);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n5598, CK => CLK, Q => 
                           n67190, QN => n63666);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n5597, CK => CLK, Q => 
                           n67189, QN => n63667);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n5596, CK => CLK, Q => 
                           n67188, QN => n63668);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n5595, CK => CLK, Q => 
                           n67187, QN => n63669);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n5594, CK => CLK, Q => 
                           n67186, QN => n63670);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n5593, CK => CLK, Q => 
                           n67185, QN => n63671);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n5592, CK => CLK, Q => 
                           n67184, QN => n63672);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n5591, CK => CLK, Q => 
                           n67183, QN => n63673);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n5590, CK => CLK, Q => 
                           n67182, QN => n63674);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n5589, CK => CLK, Q => 
                           n67181, QN => n63675);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n5588, CK => CLK, Q => 
                           n67180, QN => n63676);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n5587, CK => CLK, Q => 
                           n67179, QN => n63677);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n5586, CK => CLK, Q => 
                           n67178, QN => n63678);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n5585, CK => CLK, Q => 
                           n67177, QN => n63679);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n5584, CK => CLK, Q => 
                           n67176, QN => n63680);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n5583, CK => CLK, Q => 
                           n67175, QN => n63681);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n5582, CK => CLK, Q => 
                           n67174, QN => n63682);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n5581, CK => CLK, Q => 
                           n67173, QN => n63683);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n5580, CK => CLK, Q => 
                           n67172, QN => n63684);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n5579, CK => CLK, Q => 
                           n67171, QN => n63685);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n5578, CK => CLK, Q => 
                           n67170, QN => n63686);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n5577, CK => CLK, Q => 
                           n67169, QN => n63687);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n5576, CK => CLK, Q => 
                           n67168, QN => n63688);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n5575, CK => CLK, Q => 
                           n67167, QN => n63689);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n5574, CK => CLK, Q => 
                           n67166, QN => n63690);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n5573, CK => CLK, Q => 
                           n67165, QN => n63691);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n5572, CK => CLK, Q => 
                           n67164, QN => n63692);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n5571, CK => CLK, Q => 
                           n67163, QN => n63693);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n5570, CK => CLK, Q => 
                           n67162, QN => n63694);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n5569, CK => CLK, Q => 
                           n67161, QN => n63695);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n5568, CK => CLK, Q => 
                           n67160, QN => n63696);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n5567, CK => CLK, Q => 
                           n67159, QN => n63697);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => 
                           n67158, QN => n63572);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n67157, QN => n63573);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => 
                           n67156, QN => n63574);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n67155, QN => n63575);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => 
                           n67154, QN => n63576);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n67153, QN => n63577);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => 
                           n67152, QN => n63578);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n67151, QN => n63579);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => 
                           n67150, QN => n63580);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n67149, QN => n63581);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => 
                           n67148, QN => n63582);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n67147, QN => n63583);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => 
                           n67146, QN => n63584);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n67145, QN => n63585);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => 
                           n67144, QN => n63586);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n67143, QN => n63587);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => 
                           n67142, QN => n63588);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n67141, QN => n63589);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => 
                           n67140, QN => n63590);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => 
                           n67139, QN => n63591);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => 
                           n67138, QN => n63592);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => 
                           n67137, QN => n63593);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => 
                           n67136, QN => n63594);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => 
                           n67135, QN => n63595);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => 
                           n67134, QN => n63596);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => 
                           n67133, QN => n63597);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => 
                           n67132, QN => n63598);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => 
                           n67131, QN => n63599);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => 
                           n67130, QN => n63600);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n67129, QN => n63601);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => 
                           n67128, QN => n63602);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n67127, QN => n63603);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => 
                           n67126, QN => n63604);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n67125, QN => n63605);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => 
                           n67124, QN => n63606);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n67123, QN => n63607);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => 
                           n67122, QN => n63608);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n67121, QN => n63609);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => 
                           n67120, QN => n63610);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n67119, QN => n63611);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => 
                           n67118, QN => n63612);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n67117, QN => n63613);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => 
                           n67116, QN => n63614);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n67115, QN => n63615);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => 
                           n67114, QN => n63616);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n67113, QN => n63617);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => 
                           n67112, QN => n63618);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n67111, QN => n63619);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => 
                           n67110, QN => n63620);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n67109, QN => n63621);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n5640, CK => CLK, Q => 
                           n67108, QN => n63622);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => 
                           n67107, QN => n63623);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => 
                           n67106, QN => n63624);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => 
                           n67105, QN => n63625);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => 
                           n67104, QN => n63626);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => 
                           n67103, QN => n63627);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => 
                           n67102, QN => n63628);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => 
                           n67101, QN => n63629);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => 
                           n67100, QN => n63630);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => 
                           n67099, QN => n63631);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => 
                           n67098, QN => n63506);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n67097, QN => n63507);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => 
                           n67096, QN => n63508);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n67095, QN => n63509);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => 
                           n67094, QN => n63510);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n67093, QN => n63511);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => 
                           n67092, QN => n63512);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n67091, QN => n63513);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => 
                           n67090, QN => n63514);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n67089, QN => n63515);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => 
                           n67088, QN => n63516);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n67087, QN => n63517);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => 
                           n67086, QN => n63518);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n67085, QN => n63519);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => 
                           n67084, QN => n63520);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n67083, QN => n63521);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => 
                           n67082, QN => n63522);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n67081, QN => n63523);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => 
                           n67080, QN => n63524);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n67079, QN => n63525);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => 
                           n67078, QN => n63526);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n67077, QN => n63527);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => 
                           n67076, QN => n63528);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n67075, QN => n63529);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => 
                           n67074, QN => n63530);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n67073, QN => n63531);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => 
                           n67072, QN => n63532);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n67071, QN => n63533);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => 
                           n67070, QN => n63534);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n67069, QN => n63535);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => 
                           n67068, QN => n63536);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n67067, QN => n63537);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => 
                           n67066, QN => n63538);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n67065, QN => n63539);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => 
                           n67064, QN => n63540);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n67063, QN => n63541);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => 
                           n67062, QN => n63542);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n67061, QN => n63543);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => 
                           n67060, QN => n63544);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n67059, QN => n63545);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => 
                           n67058, QN => n63546);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n67057, QN => n63547);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => 
                           n67056, QN => n63548);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n67055, QN => n63549);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => 
                           n67054, QN => n63550);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => 
                           n67053, QN => n63551);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => 
                           n67052, QN => n63552);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => 
                           n67051, QN => n63553);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => 
                           n67050, QN => n63554);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => 
                           n67049, QN => n63555);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => 
                           n67048, QN => n63556);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => 
                           n67047, QN => n63557);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => 
                           n67046, QN => n63558);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => 
                           n67045, QN => n63559);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => 
                           n67044, QN => n63560);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n67043, QN => n63561);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => 
                           n67042, QN => n63562);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n67041, QN => n63563);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => 
                           n67040, QN => n63564);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n67039, QN => n63565);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n8967, QN => n63435);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => 
                           n8969, QN => n63436);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n8971, QN => n63437);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => 
                           n8973, QN => n63438);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n8975, QN => n63439);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => 
                           n8977, QN => n63440);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n8979, QN => n63441);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => 
                           n8981, QN => n63442);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n8983, QN => n63443);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => 
                           n8985, QN => n63444);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n8987, QN => n63445);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => 
                           n8989, QN => n63446);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n8991, QN => n63447);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => 
                           n8993, QN => n63448);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n8995, QN => n63449);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => 
                           n8997, QN => n63450);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n8999, QN => n63451);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => 
                           n9001, QN => n63452);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n9003, QN => n63453);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => 
                           n9005, QN => n63454);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n9007, QN => n63455);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => 
                           n9009, QN => n63456);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n9011, QN => n63457);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => 
                           n9013, QN => n63458);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n9015, QN => n63459);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => 
                           n9017, QN => n63460);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n9019, QN => n63461);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => 
                           n9021, QN => n63462);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n9023, QN => n63463);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => 
                           n9025, QN => n63464);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n9027, QN => n63465);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => 
                           n9029, QN => n63466);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n9031, QN => n63467);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => 
                           n9033, QN => n63468);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n9035, QN => n63469);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => 
                           n9037, QN => n63470);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n9039, QN => n63471);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => 
                           n9041, QN => n63472);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n9043, QN => n63473);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => 
                           n9045, QN => n63474);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n9047, QN => n63475);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => 
                           n9049, QN => n63476);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n9051, QN => n63477);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => 
                           n9053, QN => n63478);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n9055, QN => n63479);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => 
                           n9057, QN => n63480);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n9059, QN => n63481);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => 
                           n9061, QN => n63482);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n9063, QN => n63483);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => 
                           n9065, QN => n63484);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => n9067
                           , QN => n63485);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => n9069
                           , QN => n63486);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => n9071
                           , QN => n63487);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => n9073
                           , QN => n63488);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => n9075
                           , QN => n63489);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => n9077
                           , QN => n63490);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => n9079
                           , QN => n63491);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => n9081
                           , QN => n63492);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => n9083
                           , QN => n63493);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => n9085
                           , QN => n63494);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n67038, QN => n63302);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n67037, QN => n63303);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n67036, QN => n63304);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n67035, QN => n63305);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n67034, QN => n63306);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n67033, QN => n63307);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n67032, QN => n63308);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n67031, QN => n63309);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n67030, QN => n63310);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n67029, QN => n63311);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n67028, QN => n63312);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n67027, QN => n63313);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n67026, QN => n63314);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n67025, QN => n63315);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n67024, QN => n63316);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n67023, QN => n63317);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n67022, QN => n63318);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n67021, QN => n63319);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n67020, QN => n63320);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => 
                           n67019, QN => n63321);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => 
                           n67018, QN => n63322);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => 
                           n67017, QN => n63323);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => 
                           n67016, QN => n63324);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => 
                           n67015, QN => n63325);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => 
                           n67014, QN => n63326);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => 
                           n67013, QN => n63327);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => 
                           n67012, QN => n63328);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => 
                           n67011, QN => n63329);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => 
                           n67010, QN => n63330);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n67009, QN => n63331);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n67008, QN => n63332);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n67007, QN => n63333);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n67006, QN => n63334);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n67005, QN => n63335);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n67004, QN => n63336);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n67003, QN => n63337);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n67002, QN => n63338);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n67001, QN => n63339);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n67000, QN => n63340);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n66999, QN => n63341);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n66998, QN => n63342);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n66997, QN => n63343);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n66996, QN => n63344);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n66995, QN => n63345);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n66994, QN => n63346);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n66993, QN => n63347);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n66992, QN => n63348);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n66991, QN => n63349);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n66990, QN => n63350);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n66989, QN => n63351);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n66988, QN => n63352);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => 
                           n66987, QN => n63353);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => 
                           n66986, QN => n63354);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => 
                           n66985, QN => n63355);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => 
                           n66984, QN => n63356);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => 
                           n66983, QN => n63357);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => 
                           n66982, QN => n63358);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => 
                           n66981, QN => n63359);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => 
                           n66980, QN => n63360);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => 
                           n66979, QN => n63361);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n66978, QN => n63101);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n66977, QN => n63102);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n66976, QN => n63103);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n66975, QN => n63104);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n66974, QN => n63105);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n66973, QN => n63106);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n66972, QN => n63107);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n66971, QN => n63108);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n66970, QN => n63109);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n66969, QN => n63110);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n66968, QN => n63111);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n66967, QN => n63112);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n66966, QN => n63113);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n66965, QN => n63114);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n66964, QN => n63115);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n66963, QN => n63116);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n66962, QN => n63117);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n66961, QN => n63118);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n66960, QN => n63119);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n66959, QN => n63120);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n66958, QN => n63121);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n66957, QN => n63122);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n66956, QN => n63123);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n66955, QN => n63124);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n66954, QN => n63125);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n66953, QN => n63126);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n66952, QN => n63127);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n66951, QN => n63128);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n66950, QN => n63129);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n66949, QN => n63130);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n66948, QN => n63131);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n66947, QN => n63132);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n66946, QN => n63133);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n66945, QN => n63134);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n66944, QN => n63135);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n66943, QN => n63136);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n66942, QN => n63137);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n66941, QN => n63138);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n66940, QN => n63139);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n66939, QN => n63140);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n66938, QN => n63141);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n66937, QN => n63142);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n66936, QN => n63143);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n66935, QN => n63144);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n66934, QN => n63145);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n66933, QN => n63146);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n66932, QN => n63147);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n66931, QN => n63148);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n66930, QN => n63149);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n66929, QN => n63150);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n66928, QN => n63151);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => 
                           n66927, QN => n63152);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => 
                           n66926, QN => n63153);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => 
                           n66925, QN => n63154);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => 
                           n66924, QN => n63155);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => 
                           n66923, QN => n63156);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => 
                           n66922, QN => n63157);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => 
                           n66921, QN => n63158);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => 
                           n66920, QN => n63159);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => 
                           n66919, QN => n63160);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n66918, QN => n63368);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n66917, QN => n63369);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n66916, QN => n63370);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n66915, QN => n63371);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n66914, QN => n63372);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n66913, QN => n63373);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n66912, QN => n63374);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n66911, QN => n63375);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n66910, QN => n63376);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n66909, QN => n63377);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n66908, QN => n63378);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n66907, QN => n63379);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n66906, QN => n63380);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n66905, QN => n63381);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n66904, QN => n63382);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n66903, QN => n63383);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n66902, QN => n63384);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n66901, QN => n63385);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n66900, QN => n63386);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n66899, QN => n63387);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n66898, QN => n63388);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n66897, QN => n63389);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n66896, QN => n63390);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n66895, QN => n63391);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n66894, QN => n63392);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n66893, QN => n63393);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n66892, QN => n63394);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n66891, QN => n63395);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n66890, QN => n63396);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n66889, QN => n63397);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n66888, QN => n63398);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n66887, QN => n63399);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n66886, QN => n63400);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n66885, QN => n63401);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n66884, QN => n63402);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n66883, QN => n63403);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n66882, QN => n63404);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n66881, QN => n63405);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n66880, QN => n63406);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n66879, QN => n63407);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n66878, QN => n63408);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n66877, QN => n63409);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n66876, QN => n63410);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n66875, QN => n63411);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n66874, QN => n63412);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n66873, QN => n63413);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n66872, QN => n63414);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n66871, QN => n63415);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n66870, QN => n63416);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n66869, QN => n63417);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n66868, QN => n63418);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => 
                           n66867, QN => n63419);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => 
                           n66866, QN => n63420);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => 
                           n66865, QN => n63421);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => 
                           n66864, QN => n63422);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => 
                           n66863, QN => n63423);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => 
                           n66862, QN => n63424);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => 
                           n66861, QN => n63425);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => 
                           n66860, QN => n63426);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => 
                           n66859, QN => n63427);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n58229, QN => n63032);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n58227, QN => n63033);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n58225, QN => n63034);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n58223, QN => n63035);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n58221, QN => n63036);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n58219, QN => n63037);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n58217, QN => n63038);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n58215, QN => n63039);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n58213, QN => n63040);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n58211, QN => n63041);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n58209, QN => n63042);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n58207, QN => n63043);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n58205, QN => n63044);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n58203, QN => n63045);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n58201, QN => n63046);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n58199, QN => n63047);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n58197, QN => n63048);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n58195, QN => n63049);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n58193, QN => n63050);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n58191, QN => n63051);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n58189, QN => n63052);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n58187, QN => n63053);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n58185, QN => n63054);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n58183, QN => n63055);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n58181, QN => n63056);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n58179, QN => n63057);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n58177, QN => n63058);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n58175, QN => n63059);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n58173, QN => n63060);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n58171, QN => n63061);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n58169, QN => n63062);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n58167, QN => n63063);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n58165, QN => n63064);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n58163, QN => n63065);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n58161, QN => n63066);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n58159, QN => n63067);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n58157, QN => n63068);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n58155, QN => n63069);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n58153, QN => n63070);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n58151, QN => n63071);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n58149, QN => n63072);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n58147, QN => n63073);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n58145, QN => n63074);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n58143, QN => n63075);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n58141, QN => n63076);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n58139, QN => n63077);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n58137, QN => n63078);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n58135, QN => n63079);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n58134, QN => n63080);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n58132, QN => n63081);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n58130, QN => n63082);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n58128, QN => n63083);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n58126, QN => n63084);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n58124, QN => n63085);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n58122, QN => n63086);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n58120, QN => n63087);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n58118, QN => n63088);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n58116, QN => n63089);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n58114, QN => n63090);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n58112, QN => n63091);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n58498, QN => n62965);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n58497, QN => n62966);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n58496, QN => n62967);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n58495, QN => n62968);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n58494, QN => n62969);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n58493, QN => n62970);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n58492, QN => n62971);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n58491, QN => n62972);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n58490, QN => n62973);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n58489, QN => n62974);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n58488, QN => n62975);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n58487, QN => n62976);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n58486, QN => n62977);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n58485, QN => n62978);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n58484, QN => n62979);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n58483, QN => n62980);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n58482, QN => n62981);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n58481, QN => n62982);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n58480, QN => n62983);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n58479, QN => n62984);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n58478, QN => n62985);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n58477, QN => n62986);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n58476, QN => n62987);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n58475, QN => n62988);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n58474, QN => n62989);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n58473, QN => n62990);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n58472, QN => n62991);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n58471, QN => n62992);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n58470, QN => n62993);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n58469, QN => n62994);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n58468, QN => n62995);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n58467, QN => n62996);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n58466, QN => n62997);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n58465, QN => n62998);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n58464, QN => n62999);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n58463, QN => n63000);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n58462, QN => n63001);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n58461, QN => n63002);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n58460, QN => n63003);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n58459, QN => n63004);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n58458, QN => n63005);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n58457, QN => n63006);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n58456, QN => n63007);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n58455, QN => n63008);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n58454, QN => n63009);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n58453, QN => n63010);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n58452, QN => n63011);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n58451, QN => n63012);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n58450, QN => n63013);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n58449, QN => n63014);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n58448, QN => n63015);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => 
                           n58447, QN => n63016);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => 
                           n58446, QN => n63017);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => 
                           n58445, QN => n63018);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => 
                           n58444, QN => n63019);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => 
                           n58443, QN => n63020);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => 
                           n58442, QN => n63021);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => 
                           n58441, QN => n63022);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => 
                           n58440, QN => n63023);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => 
                           n58439, QN => n63024);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n58714, QN => n63235);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n58713, QN => n63236);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n58712, QN => n63237);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n58711, QN => n63238);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n58710, QN => n63239);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n58709, QN => n63240);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n58708, QN => n63241);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n58707, QN => n63242);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n58706, QN => n63243);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n58705, QN => n63244);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n58704, QN => n63245);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n58703, QN => n63246);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n58702, QN => n63247);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n58701, QN => n63248);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n58700, QN => n63249);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n58699, QN => n63250);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n58698, QN => n63251);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n58697, QN => n63252);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n58696, QN => n63253);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n58695, QN => n63254);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n58694, QN => n63255);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n58693, QN => n63256);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n58692, QN => n63257);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n58691, QN => n63258);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n58690, QN => n63259);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n58689, QN => n63260);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n58688, QN => n63261);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n58687, QN => n63262);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n58686, QN => n63263);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n58685, QN => n63264);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n58684, QN => n63265);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n58683, QN => n63266);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n58682, QN => n63267);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n58681, QN => n63268);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n58680, QN => n63269);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n58679, QN => n63270);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n58678, QN => n63271);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n58677, QN => n63272);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n58676, QN => n63273);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n58675, QN => n63274);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n58674, QN => n63275);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n58673, QN => n63276);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n58672, QN => n63277);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n58671, QN => n63278);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n58670, QN => n63279);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n58669, QN => n63280);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n58668, QN => n63281);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n58667, QN => n63282);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n58742, QN => n63283);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n58741, QN => n63284);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n58740, QN => n63285);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => 
                           n58739, QN => n63286);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => 
                           n58738, QN => n63287);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => 
                           n58737, QN => n63288);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => 
                           n58736, QN => n63289);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n58735, QN => n63290);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n58734, QN => n63291);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => 
                           n58733, QN => n63292);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => 
                           n58732, QN => n63293);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => 
                           n58731, QN => n63294);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n58282, QN => n63167);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n58281, QN => n63168);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n58280, QN => n63169);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n58279, QN => n63170);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n58278, QN => n63171);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n58277, QN => n63172);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n58276, QN => n63173);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n58275, QN => n63174);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n58274, QN => n63175);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n58273, QN => n63176);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n58272, QN => n63177);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n58271, QN => n63178);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n58270, QN => n63179);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n58269, QN => n63180);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n58268, QN => n63181);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n58267, QN => n63182);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n58266, QN => n63183);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n58265, QN => n63184);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n58264, QN => n63185);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n58263, QN => n63186);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n58262, QN => n63187);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n58261, QN => n63188);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n58260, QN => n63189);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n58259, QN => n63190);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n58258, QN => n63191);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n58257, QN => n63192);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n58256, QN => n63193);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n58255, QN => n63194);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n58254, QN => n63195);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n58253, QN => n63196);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n58252, QN => n63197);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n58251, QN => n63198);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n58250, QN => n63199);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n58249, QN => n63200);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n58248, QN => n63201);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n58247, QN => n63202);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n58246, QN => n63203);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n58245, QN => n63204);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n58244, QN => n63205);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n58243, QN => n63206);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n58242, QN => n63207);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n58241, QN => n63208);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n58240, QN => n63209);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n58239, QN => n63210);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n58238, QN => n63211);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n58237, QN => n63212);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n58236, QN => n63213);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => 
                           n58235, QN => n63214);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => 
                           n58294, QN => n63215);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => 
                           n58293, QN => n63216);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n58292, QN => n63217);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n58291, QN => n63218);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n58290, QN => n63219);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n58289, QN => n63220);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n58288, QN => n63221);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n58287, QN => n63222);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n58286, QN => n63223);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n58285, QN => n63224);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n58284, QN => n63225);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n58283, QN => n63226);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => 
                           n66858, QN => n62697);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n66857, QN => n62699);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n66856, QN => n62700);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n66855, QN => n62701);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => n8895
                           , QN => n62627);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => n8896
                           , QN => n62629);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => n8897
                           , QN => n62630);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => n8898
                           , QN => n62631);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => 
                           n58654, QN => n62893);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n58653, QN => n62895);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n58652, QN => n62896);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n58651, QN => n62897);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7482, CK => CLK, Q => 
                           n56603, QN => n61967);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7481, CK => CLK, Q => 
                           n56627, QN => n61969);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7480, CK => CLK, Q => 
                           n56651, QN => n61971);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7479, CK => CLK, Q => 
                           n56675, QN => n61973);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7478, CK => CLK, Q => 
                           n56699, QN => n61975);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7477, CK => CLK, Q => 
                           n56723, QN => n61977);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7476, CK => CLK, Q => 
                           n56747, QN => n61979);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7475, CK => CLK, Q => 
                           n56771, QN => n61981);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7474, CK => CLK, Q => 
                           n56795, QN => n61983);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7473, CK => CLK, Q => 
                           n56819, QN => n61985);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7472, CK => CLK, Q => 
                           n56843, QN => n61987);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7471, CK => CLK, Q => 
                           n56867, QN => n61989);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7470, CK => CLK, Q => 
                           n56891, QN => n61991);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7469, CK => CLK, Q => 
                           n56915, QN => n61993);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7468, CK => CLK, Q => 
                           n56939, QN => n61995);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7467, CK => CLK, Q => 
                           n56963, QN => n61997);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7466, CK => CLK, Q => 
                           n56987, QN => n61999);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7465, CK => CLK, Q => 
                           n57011, QN => n62001);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7464, CK => CLK, Q => 
                           n57035, QN => n62003);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7463, CK => CLK, Q => 
                           n57059, QN => n62005);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7462, CK => CLK, Q => 
                           n57083, QN => n62007);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7461, CK => CLK, Q => 
                           n57107, QN => n62009);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7460, CK => CLK, Q => 
                           n57131, QN => n62011);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7459, CK => CLK, Q => 
                           n57155, QN => n62013);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7458, CK => CLK, Q => 
                           n57179, QN => n62015);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7457, CK => CLK, Q => 
                           n57203, QN => n62017);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7456, CK => CLK, Q => 
                           n57227, QN => n62019);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7455, CK => CLK, Q => 
                           n57251, QN => n62021);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7454, CK => CLK, Q => 
                           n57275, QN => n62023);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7453, CK => CLK, Q => 
                           n57299, QN => n62025);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7452, CK => CLK, Q => 
                           n57323, QN => n62027);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7451, CK => CLK, Q => 
                           n57347, QN => n62029);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7450, CK => CLK, Q => 
                           n57371, QN => n62031);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7449, CK => CLK, Q => 
                           n57395, QN => n62033);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7448, CK => CLK, Q => 
                           n57419, QN => n62035);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7447, CK => CLK, Q => 
                           n57443, QN => n62037);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7446, CK => CLK, Q => 
                           n57467, QN => n62039);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7445, CK => CLK, Q => 
                           n57491, QN => n62041);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7444, CK => CLK, Q => 
                           n57515, QN => n62043);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7443, CK => CLK, Q => 
                           n57539, QN => n62045);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7442, CK => CLK, Q => 
                           n57563, QN => n62047);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7441, CK => CLK, Q => 
                           n57587, QN => n62049);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7440, CK => CLK, Q => 
                           n57611, QN => n62051);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7439, CK => CLK, Q => 
                           n57635, QN => n62053);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7438, CK => CLK, Q => 
                           n57659, QN => n62055);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7437, CK => CLK, Q => 
                           n57683, QN => n62057);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7436, CK => CLK, Q => 
                           n57707, QN => n62059);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7435, CK => CLK, Q => 
                           n57731, QN => n62061);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7434, CK => CLK, Q => 
                           n57755, QN => n62063);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7433, CK => CLK, Q => 
                           n57779, QN => n62065);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7432, CK => CLK, Q => n57803
                           , QN => n62067);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7431, CK => CLK, Q => n57827
                           , QN => n62069);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7430, CK => CLK, Q => n57851
                           , QN => n62071);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7429, CK => CLK, Q => n57875
                           , QN => n62073);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7428, CK => CLK, Q => n57899
                           , QN => n62075);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7427, CK => CLK, Q => n57923
                           , QN => n62077);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7426, CK => CLK, Q => n57947
                           , QN => n62079);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7425, CK => CLK, Q => n57971
                           , QN => n62081);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7424, CK => CLK, Q => n57995
                           , QN => n62083);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7423, CK => CLK, Q => n58028
                           , QN => n62085);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n58110, QN => n62499);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n58109, QN => n62500);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n58108, QN => n62501);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n58107, QN => n62502);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n58106, QN => n62503);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n58105, QN => n62504);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n58104, QN => n62505);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n58103, QN => n62506);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n58102, QN => n62507);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n58101, QN => n62508);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n58100, QN => n62509);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n58099, QN => n62510);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n58098, QN => n62511);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n58097, QN => n62512);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n58096, QN => n62513);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n58095, QN => n62514);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n58094, QN => n62515);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n58093, QN => n62516);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n58092, QN => n62517);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n58091, QN => n62518);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n58090, QN => n62519);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n58089, QN => n62520);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n58088, QN => n62521);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n58087, QN => n62522);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n58086, QN => n62523);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n58085, QN => n62524);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => 
                           n58084, QN => n62525);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => 
                           n58083, QN => n62526);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => 
                           n58082, QN => n62527);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n58081, QN => n62528);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n58080, QN => n62529);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n58079, QN => n62530);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n58078, QN => n62531);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n58077, QN => n62532);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n58076, QN => n62533);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n58075, QN => n62534);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n58074, QN => n62535);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n58073, QN => n62536);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n58072, QN => n62537);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n58071, QN => n62538);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n58070, QN => n62539);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n58069, QN => n62540);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n58068, QN => n62541);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n58067, QN => n62542);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n58066, QN => n62543);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n58065, QN => n62544);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n58064, QN => n62545);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n58063, QN => n62546);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n58062, QN => n62547);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n58061, QN => n62548);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => n58060
                           , QN => n62549);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => n58059
                           , QN => n62550);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => n58058
                           , QN => n62551);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => n58057
                           , QN => n62552);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => n58056
                           , QN => n62553);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => n58055
                           , QN => n62554);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => n58054
                           , QN => n62555);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => n58053
                           , QN => n62556);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => n58052
                           , QN => n62557);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => n58051
                           , QN => n62558);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => 
                           n58842, QN => n62363);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => 
                           n58841, QN => n62364);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => 
                           n58840, QN => n62365);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => 
                           n58839, QN => n62366);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => 
                           n58838, QN => n62367);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => 
                           n58837, QN => n62368);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => 
                           n58836, QN => n62369);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => 
                           n58835, QN => n62370);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => 
                           n58834, QN => n62371);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => 
                           n58833, QN => n62372);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => 
                           n58832, QN => n62373);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => 
                           n58831, QN => n62374);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => 
                           n58830, QN => n62375);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => 
                           n58829, QN => n62376);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => 
                           n58828, QN => n62377);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => 
                           n58827, QN => n62378);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => 
                           n58826, QN => n62379);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => 
                           n58825, QN => n62380);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => 
                           n58824, QN => n62381);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => 
                           n58823, QN => n62382);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => 
                           n58822, QN => n62383);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => 
                           n58821, QN => n62384);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => 
                           n58820, QN => n62385);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => 
                           n58819, QN => n62386);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => 
                           n58818, QN => n62387);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n7137, CK => CLK, Q => 
                           n58817, QN => n62388);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n7136, CK => CLK, Q => 
                           n58816, QN => n62389);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n7135, CK => CLK, Q => 
                           n58815, QN => n62390);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7134, CK => CLK, Q => 
                           n58814, QN => n62391);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7133, CK => CLK, Q => 
                           n58813, QN => n62392);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7132, CK => CLK, Q => 
                           n58812, QN => n62393);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7131, CK => CLK, Q => 
                           n58811, QN => n62394);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7130, CK => CLK, Q => 
                           n58810, QN => n62395);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7129, CK => CLK, Q => 
                           n58809, QN => n62396);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7128, CK => CLK, Q => 
                           n58808, QN => n62397);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7127, CK => CLK, Q => 
                           n58807, QN => n62398);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7126, CK => CLK, Q => 
                           n58806, QN => n62399);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7125, CK => CLK, Q => 
                           n58805, QN => n62400);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7124, CK => CLK, Q => 
                           n58804, QN => n62401);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7123, CK => CLK, Q => 
                           n58803, QN => n62402);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7122, CK => CLK, Q => 
                           n58802, QN => n62403);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7121, CK => CLK, Q => 
                           n58801, QN => n62404);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7120, CK => CLK, Q => 
                           n58800, QN => n62405);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7119, CK => CLK, Q => 
                           n58799, QN => n62406);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           n56020, QN => n62407);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7117, CK => CLK, Q => 
                           n56047, QN => n62408);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7116, CK => CLK, Q => 
                           n56074, QN => n62409);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7115, CK => CLK, Q => 
                           n56101, QN => n62410);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7114, CK => CLK, Q => 
                           n58798, QN => n62411);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7113, CK => CLK, Q => 
                           n58797, QN => n62412);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7112, CK => CLK, Q => n58796
                           , QN => n62413);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7111, CK => CLK, Q => n58795
                           , QN => n62414);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7110, CK => CLK, Q => n58794
                           , QN => n62415);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7109, CK => CLK, Q => n58793
                           , QN => n62416);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7108, CK => CLK, Q => n58792
                           , QN => n62417);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => n58791
                           , QN => n62418);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => n58790
                           , QN => n62419);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => n58789
                           , QN => n62420);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => n58788
                           , QN => n62421);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => n58787
                           , QN => n62422);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => 
                           n66854, QN => n62230);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => 
                           n66853, QN => n62231);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => 
                           n66852, QN => n62232);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => 
                           n66851, QN => n62233);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => 
                           n66850, QN => n62234);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => 
                           n66849, QN => n62235);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => 
                           n66848, QN => n62236);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => 
                           n66847, QN => n62237);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => 
                           n66846, QN => n62238);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => 
                           n66845, QN => n62239);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => 
                           n66844, QN => n62240);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => 
                           n66843, QN => n62241);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => 
                           n66842, QN => n62242);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => 
                           n66841, QN => n62243);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => 
                           n66840, QN => n62244);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => 
                           n66839, QN => n62245);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => 
                           n66838, QN => n62246);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => 
                           n66837, QN => n62247);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => 
                           n66836, QN => n62248);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => 
                           n66835, QN => n62249);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => 
                           n66834, QN => n62250);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => 
                           n66833, QN => n62251);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => 
                           n66832, QN => n62252);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => 
                           n66831, QN => n62253);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => 
                           n66830, QN => n62254);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => 
                           n66829, QN => n62255);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => 
                           n66828, QN => n62256);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => 
                           n66827, QN => n62257);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => 
                           n66826, QN => n62258);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => 
                           n66825, QN => n62259);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => 
                           n66824, QN => n62260);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => 
                           n66823, QN => n62261);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => 
                           n66822, QN => n62262);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => 
                           n66821, QN => n62263);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => 
                           n66820, QN => n62264);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => 
                           n66819, QN => n62265);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => 
                           n66818, QN => n62266);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => 
                           n66817, QN => n62267);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => 
                           n66816, QN => n62268);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => 
                           n66815, QN => n62269);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => 
                           n66814, QN => n62270);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => 
                           n66813, QN => n62271);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => 
                           n66812, QN => n62272);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => 
                           n66811, QN => n62273);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => 
                           n66810, QN => n62274);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => 
                           n66809, QN => n62275);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => 
                           n66808, QN => n62276);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => 
                           n66807, QN => n62277);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => 
                           n66806, QN => n62278);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => 
                           n66805, QN => n62279);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => n66804
                           , QN => n62280);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => n66803
                           , QN => n62281);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => n66802
                           , QN => n62282);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => n66801
                           , QN => n62283);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => n66800
                           , QN => n62284);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => n66799
                           , QN => n62285);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => n66798
                           , QN => n62286);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => n66797
                           , QN => n62287);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => n66796
                           , QN => n62288);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => n66795
                           , QN => n62289);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => 
                           n66794, QN => n62163);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => 
                           n66793, QN => n62164);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => 
                           n66792, QN => n62165);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => 
                           n66791, QN => n62166);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => 
                           n66790, QN => n62167);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => 
                           n66789, QN => n62168);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => 
                           n66788, QN => n62169);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => 
                           n66787, QN => n62170);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => 
                           n66786, QN => n62171);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => 
                           n66785, QN => n62172);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => 
                           n66784, QN => n62173);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => 
                           n66783, QN => n62174);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => 
                           n66782, QN => n62175);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => 
                           n66781, QN => n62176);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => 
                           n66780, QN => n62177);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => 
                           n66779, QN => n62178);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => 
                           n66778, QN => n62179);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => 
                           n66777, QN => n62180);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => 
                           n66776, QN => n62181);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => 
                           n66775, QN => n62182);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => 
                           n66774, QN => n62183);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => 
                           n66773, QN => n62184);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => 
                           n66772, QN => n62185);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => 
                           n66771, QN => n62186);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => 
                           n66770, QN => n62187);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => 
                           n66769, QN => n62188);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => 
                           n66768, QN => n62189);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => 
                           n66767, QN => n62190);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => 
                           n66766, QN => n62191);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => 
                           n66765, QN => n62192);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => 
                           n66764, QN => n62193);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => 
                           n66763, QN => n62194);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => 
                           n66762, QN => n62195);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => 
                           n66761, QN => n62196);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => 
                           n66760, QN => n62197);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => 
                           n66759, QN => n62198);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => 
                           n66758, QN => n62199);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => 
                           n66757, QN => n62200);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => 
                           n66756, QN => n62201);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => 
                           n66755, QN => n62202);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => 
                           n66754, QN => n62203);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => 
                           n66753, QN => n62204);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => 
                           n66752, QN => n62205);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => 
                           n66751, QN => n62206);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => 
                           n66750, QN => n62207);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => 
                           n66749, QN => n62208);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => 
                           n66748, QN => n62209);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => 
                           n66747, QN => n62210);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => 
                           n66746, QN => n62211);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => 
                           n66745, QN => n62212);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => n66744
                           , QN => n62213);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => n66743
                           , QN => n62214);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => n66742
                           , QN => n62215);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => n66741
                           , QN => n62216);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => n66740
                           , QN => n62217);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => n66739
                           , QN => n62218);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => n66738
                           , QN => n62219);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => n66737
                           , QN => n62220);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => n66736
                           , QN => n62221);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => n66735
                           , QN => n62222);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n66734, QN => n62429);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n66733, QN => n62430);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n66732, QN => n62431);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n66731, QN => n62432);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n66730, QN => n62433);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n66729, QN => n62434);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n66728, QN => n62435);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n66727, QN => n62436);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n66726, QN => n62437);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n66725, QN => n62438);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n66724, QN => n62439);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n66723, QN => n62440);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n66722, QN => n62441);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n66721, QN => n62442);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n66720, QN => n62443);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n66719, QN => n62444);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n66718, QN => n62445);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n66717, QN => n62446);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n66716, QN => n62447);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n66715, QN => n62448);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           n66714, QN => n62449);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           n66713, QN => n62450);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           n66712, QN => n62451);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           n66711, QN => n62452);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           n66710, QN => n62453);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => 
                           n66709, QN => n62454);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           n66708, QN => n62455);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           n66707, QN => n62456);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => 
                           n66706, QN => n62457);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n66705, QN => n62458);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n66704, QN => n62459);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n66703, QN => n62460);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n66702, QN => n62461);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n66701, QN => n62462);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n66700, QN => n62463);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n66699, QN => n62464);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n66698, QN => n62465);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n66697, QN => n62466);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n66696, QN => n62467);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n66695, QN => n62468);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => 
                           n66694, QN => n62469);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => 
                           n66693, QN => n62470);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => 
                           n66692, QN => n62471);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => 
                           n66691, QN => n62472);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => 
                           n66690, QN => n62473);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => 
                           n66689, QN => n62474);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => 
                           n66688, QN => n62475);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => 
                           n66687, QN => n62476);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => 
                           n66686, QN => n62477);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => 
                           n66685, QN => n62478);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => n66684
                           , QN => n62479);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => n66683
                           , QN => n62480);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => n66682
                           , QN => n62481);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => n66681
                           , QN => n62482);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => n66680
                           , QN => n62483);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => n66679
                           , QN => n62484);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => n66678
                           , QN => n62485);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => n66677
                           , QN => n62486);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => n66676
                           , QN => n62487);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => n66675
                           , QN => n62488);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => 
                           n59088, QN => n62296);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => 
                           n59087, QN => n62297);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => 
                           n59086, QN => n62298);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => 
                           n59085, QN => n62299);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => 
                           n59084, QN => n62300);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => 
                           n59083, QN => n62301);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => 
                           n59082, QN => n62302);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => 
                           n59081, QN => n62303);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => 
                           n59080, QN => n62304);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => 
                           n59079, QN => n62305);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => 
                           n59078, QN => n62306);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => 
                           n59077, QN => n62307);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => 
                           n59076, QN => n62308);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => 
                           n59075, QN => n62309);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => 
                           n59074, QN => n62310);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => 
                           n59073, QN => n62311);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => 
                           n59072, QN => n62312);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => 
                           n59071, QN => n62313);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => 
                           n59070, QN => n62314);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => 
                           n59069, QN => n62315);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => 
                           n59068, QN => n62316);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => 
                           n59067, QN => n62317);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => 
                           n59066, QN => n62318);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => 
                           n59065, QN => n62319);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n7202, CK => CLK, Q => 
                           n59064, QN => n62320);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => 
                           n59063, QN => n62321);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => 
                           n59062, QN => n62322);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => 
                           n59061, QN => n62323);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => 
                           n59060, QN => n62324);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => 
                           n59059, QN => n62325);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => 
                           n59058, QN => n62326);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => 
                           n59057, QN => n62327);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => 
                           n59056, QN => n62328);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => 
                           n59055, QN => n62329);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => 
                           n59054, QN => n62330);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => 
                           n59053, QN => n62331);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => 
                           n59052, QN => n62332);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => 
                           n59051, QN => n62333);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => 
                           n59050, QN => n62334);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => 
                           n59049, QN => n62335);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => 
                           n59048, QN => n62336);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => 
                           n59047, QN => n62337);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => 
                           n59046, QN => n62338);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => 
                           n59045, QN => n62339);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => 
                           n59044, QN => n62340);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => 
                           n59043, QN => n62341);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => 
                           n59042, QN => n62342);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => 
                           n59041, QN => n62343);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => 
                           n59040, QN => n62344);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => 
                           n59039, QN => n62345);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => n59038
                           , QN => n62346);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => n59037
                           , QN => n62347);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => n59036
                           , QN => n62348);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => n59035
                           , QN => n62349);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => n59034
                           , QN => n62350);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => n59033
                           , QN => n62351);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => n59032
                           , QN => n62352);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => n59031
                           , QN => n62353);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => n59030
                           , QN => n62354);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => n59029
                           , QN => n62355);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => 
                           n66674, QN => n62096);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => 
                           n66673, QN => n62097);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => 
                           n66672, QN => n62098);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => 
                           n66671, QN => n62099);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => 
                           n66670, QN => n62100);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => 
                           n66669, QN => n62101);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => 
                           n66668, QN => n62102);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => 
                           n66667, QN => n62103);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => 
                           n66666, QN => n62104);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => 
                           n66665, QN => n62105);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => 
                           n66664, QN => n62106);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => 
                           n66663, QN => n62107);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => 
                           n66662, QN => n62108);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => 
                           n66661, QN => n62109);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => 
                           n66660, QN => n62110);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => 
                           n66659, QN => n62111);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => 
                           n66658, QN => n62112);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => 
                           n66657, QN => n62113);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => 
                           n66656, QN => n62114);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => 
                           n66655, QN => n62115);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => 
                           n66654, QN => n62116);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => 
                           n66653, QN => n62117);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => 
                           n66652, QN => n62118);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => 
                           n66651, QN => n62119);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => 
                           n66650, QN => n62120);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => 
                           n66649, QN => n62121);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => 
                           n66648, QN => n62122);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => 
                           n66647, QN => n62123);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => 
                           n66646, QN => n62124);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => 
                           n66645, QN => n62125);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => 
                           n66644, QN => n62126);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => 
                           n66643, QN => n62127);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => 
                           n66642, QN => n62128);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => 
                           n66641, QN => n62129);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => 
                           n66640, QN => n62130);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => 
                           n66639, QN => n62131);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => 
                           n66638, QN => n62132);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => 
                           n66637, QN => n62133);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => 
                           n66636, QN => n62134);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => 
                           n66635, QN => n62135);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => 
                           n66634, QN => n62136);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => 
                           n66633, QN => n62137);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => 
                           n66632, QN => n62138);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => 
                           n66631, QN => n62139);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => 
                           n66630, QN => n62140);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => 
                           n66629, QN => n62141);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => 
                           n66628, QN => n62142);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => 
                           n66627, QN => n62143);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => 
                           n66626, QN => n62144);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => 
                           n66625, QN => n62145);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => n66624
                           , QN => n62146);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => n66623
                           , QN => n62147);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => n66622
                           , QN => n62148);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => n66621
                           , QN => n62149);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => n66620
                           , QN => n62150);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => n66619
                           , QN => n62151);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => n66618
                           , QN => n62152);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => n66617
                           , QN => n62153);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => n66616
                           , QN => n62154);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => n66615
                           , QN => n62155);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n58366, QN => n62565);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n58365, QN => n62566);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n58364, QN => n62567);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n58363, QN => n62568);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n58362, QN => n62569);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n58361, QN => n62570);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n58360, QN => n62571);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n58359, QN => n62572);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n58358, QN => n62573);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n58357, QN => n62574);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n58356, QN => n62575);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n58355, QN => n62576);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n58354, QN => n62577);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n58353, QN => n62578);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n58352, QN => n62579);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n58351, QN => n62580);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n58350, QN => n62581);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n58349, QN => n62582);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n58348, QN => n62583);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n58347, QN => n62584);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n58346, QN => n62585);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n58345, QN => n62586);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n58344, QN => n62587);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n58343, QN => n62588);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n58342, QN => n62589);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n58341, QN => n62590);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n58340, QN => n62591);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n58339, QN => n62592);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n58338, QN => n62593);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n58337, QN => n62594);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n58336, QN => n62595);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n58335, QN => n62596);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n58334, QN => n62597);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n58333, QN => n62598);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n58332, QN => n62599);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n58331, QN => n62600);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n58330, QN => n62601);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n58329, QN => n62602);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n58328, QN => n62603);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n58327, QN => n62604);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n58326, QN => n62605);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n58325, QN => n62606);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n58324, QN => n62607);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n58323, QN => n62608);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n58322, QN => n62609);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n58321, QN => n62610);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n58320, QN => n62611);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n58319, QN => n62612);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n58318, QN => n62613);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n58317, QN => n62614);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => n58316
                           , QN => n62615);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => n58315
                           , QN => n62616);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => n58314
                           , QN => n62617);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => n58313
                           , QN => n62618);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => n58312
                           , QN => n62619);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => n58311
                           , QN => n62620);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => n58310
                           , QN => n62621);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => n58309
                           , QN => n62622);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => n58308
                           , QN => n62623);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => n58307
                           , QN => n62624);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n56597, QN => n62832);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n56621, QN => n62833);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n56645, QN => n62834);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n56669, QN => n62835);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n56693, QN => n62836);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n56717, QN => n62837);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n56741, QN => n62838);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n56765, QN => n62839);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n56789, QN => n62840);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n56813, QN => n62841);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n56837, QN => n62842);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n56861, QN => n62843);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n56885, QN => n62844);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n56909, QN => n62845);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n56933, QN => n62846);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n56957, QN => n62847);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n56981, QN => n62848);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n57005, QN => n62849);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n57029, QN => n62850);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => 
                           n57053, QN => n62851);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => 
                           n57077, QN => n62852);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => 
                           n57101, QN => n62853);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => 
                           n57125, QN => n62854);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => 
                           n57149, QN => n62855);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => 
                           n57173, QN => n62856);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => 
                           n57197, QN => n62857);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => 
                           n57221, QN => n62858);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => 
                           n57245, QN => n62859);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => 
                           n57269, QN => n62860);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n57293, QN => n62861);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n57317, QN => n62862);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n57341, QN => n62863);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n57365, QN => n62864);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n57389, QN => n62865);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n57413, QN => n62866);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n57437, QN => n62867);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n57461, QN => n62868);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n57485, QN => n62869);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n57509, QN => n62870);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n57533, QN => n62871);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n57557, QN => n62872);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n57581, QN => n62873);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n57605, QN => n62874);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n57629, QN => n62875);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n57653, QN => n62876);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n57677, QN => n62877);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n57701, QN => n62878);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n57725, QN => n62879);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n57749, QN => n62880);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n57773, QN => n62881);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n57797, QN => n62882);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => 
                           n57821, QN => n62883);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => 
                           n57845, QN => n62884);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => 
                           n57869, QN => n62885);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => 
                           n57893, QN => n62886);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => 
                           n57917, QN => n62887);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => 
                           n57941, QN => n62888);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => 
                           n57965, QN => n62889);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => 
                           n57989, QN => n62890);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => 
                           n58013, QN => n62891);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n56609, QN => n62766);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n56633, QN => n62767);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n56657, QN => n62768);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n56681, QN => n62769);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n56705, QN => n62770);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n56729, QN => n62771);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n56753, QN => n62772);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n56777, QN => n62773);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n56801, QN => n62774);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n56825, QN => n62775);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n56849, QN => n62776);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n56873, QN => n62777);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n56897, QN => n62778);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n56921, QN => n62779);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n56945, QN => n62780);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n56969, QN => n62781);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n56993, QN => n62782);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n57017, QN => n62783);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n57041, QN => n62784);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n57065, QN => n62785);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n57089, QN => n62786);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n57113, QN => n62787);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n57137, QN => n62788);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n57161, QN => n62789);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n57185, QN => n62790);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n57209, QN => n62791);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n57233, QN => n62792);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n57257, QN => n62793);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n57281, QN => n62794);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n57305, QN => n62795);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n57329, QN => n62796);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n57353, QN => n62797);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n57377, QN => n62798);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n57401, QN => n62799);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n57425, QN => n62800);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n57449, QN => n62801);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n57473, QN => n62802);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n57497, QN => n62803);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n57521, QN => n62804);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n57545, QN => n62805);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n57569, QN => n62806);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n57593, QN => n62807);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n57617, QN => n62808);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n57641, QN => n62809);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n57665, QN => n62810);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n57689, QN => n62811);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n57713, QN => n62812);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n57737, QN => n62813);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n57761, QN => n62814);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n57785, QN => n62815);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n57809, QN => n62816);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => 
                           n57833, QN => n62817);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => 
                           n57857, QN => n62818);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => 
                           n57881, QN => n62819);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => 
                           n57905, QN => n62820);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => 
                           n57929, QN => n62821);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => 
                           n57953, QN => n62822);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => 
                           n57977, QN => n62823);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => 
                           n58001, QN => n62824);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => 
                           n58036, QN => n62825);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n66614, QN => n62702);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n66613, QN => n62703);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n66612, QN => n62704);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n66611, QN => n62705);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n66610, QN => n62706);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n66609, QN => n62707);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n66608, QN => n62708);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n66607, QN => n62709);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n66606, QN => n62710);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n66605, QN => n62711);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n66604, QN => n62712);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n66603, QN => n62713);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n66602, QN => n62714);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n66601, QN => n62715);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n66600, QN => n62716);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n66599, QN => n62717);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n66598, QN => n62718);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n66597, QN => n62719);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n66596, QN => n62720);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n66595, QN => n62721);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n66594, QN => n62722);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n66593, QN => n62723);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n66592, QN => n62724);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n66591, QN => n62725);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n66590, QN => n62726);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n66589, QN => n62727);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n66588, QN => n62728);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n66587, QN => n62729);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n66586, QN => n62730);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n66585, QN => n62731);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n66584, QN => n62732);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n66583, QN => n62733);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n66582, QN => n62734);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n66581, QN => n62735);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n66580, QN => n62736);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n66579, QN => n62737);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n66578, QN => n62738);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n66577, QN => n62739);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n66576, QN => n62740);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n66575, QN => n62741);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n66574, QN => n62742);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n66573, QN => n62743);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n66572, QN => n62744);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n66571, QN => n62745);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n66570, QN => n62746);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n66569, QN => n62747);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n66568, QN => n62748);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n66567, QN => n62749);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n66566, QN => n62750);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n66565, QN => n62751);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n66564, QN => n62752);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => 
                           n66563, QN => n62753);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => 
                           n66562, QN => n62754);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => 
                           n66561, QN => n62755);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => 
                           n66560, QN => n62756);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => 
                           n66559, QN => n62757);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => 
                           n66558, QN => n62758);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => 
                           n66557, QN => n62759);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => 
                           n66556, QN => n62760);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => 
                           n66555, QN => n62761);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => n8899
                           , QN => n62632);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => n8900
                           , QN => n62633);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => n8901
                           , QN => n62634);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => n8902
                           , QN => n62635);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => n8903
                           , QN => n62636);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => n8904
                           , QN => n62637);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => n8905
                           , QN => n62638);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => n8906
                           , QN => n62639);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => n8907
                           , QN => n62640);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => n8908
                           , QN => n62641);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => n8909
                           , QN => n62642);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => n8910
                           , QN => n62643);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => n8911
                           , QN => n62644);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => n8912
                           , QN => n62645);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => n8913
                           , QN => n62646);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => n8914
                           , QN => n62647);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => n8915
                           , QN => n62648);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => n8916
                           , QN => n62649);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => n8917
                           , QN => n62650);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => n8918
                           , QN => n62651);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => n8919
                           , QN => n62652);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => n8920
                           , QN => n62653);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => n8921
                           , QN => n62654);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => n8922
                           , QN => n62655);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => n8923
                           , QN => n62656);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => n8924
                           , QN => n62657);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => n8925
                           , QN => n62658);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => n8926
                           , QN => n62659);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => n8927
                           , QN => n62660);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => n8928
                           , QN => n62661);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => n8929
                           , QN => n62662);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => n8930
                           , QN => n62663);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => n8931
                           , QN => n62664);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => n8932
                           , QN => n62665);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => n8933
                           , QN => n62666);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => n8934
                           , QN => n62667);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => n8935
                           , QN => n62668);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => n8936
                           , QN => n62669);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => n8937
                           , QN => n62670);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => n8938
                           , QN => n62671);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => n8939
                           , QN => n62672);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => n8940
                           , QN => n62673);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => n8941
                           , QN => n62674);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => n8942
                           , QN => n62675);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => n8943
                           , QN => n62676);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => n8944
                           , QN => n62677);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => n8945
                           , QN => n62678);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => n8946
                           , QN => n62679);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => n8947
                           , QN => n62680);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => n8948
                           , QN => n62681);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => n8949,
                           QN => n62682);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => n8950,
                           QN => n62683);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => n8951,
                           QN => n62684);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => n8952,
                           QN => n62685);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => n8953,
                           QN => n62686);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => n8954,
                           QN => n62687);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => n8955,
                           QN => n62688);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => n8956,
                           QN => n62689);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => n8957,
                           QN => n62690);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => n8958,
                           QN => n62691);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n58650, QN => n62898);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n58649, QN => n62899);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n58648, QN => n62900);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n58647, QN => n62901);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n58646, QN => n62902);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n58645, QN => n62903);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n58644, QN => n62904);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n58643, QN => n62905);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n56791, QN => n62906);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n56815, QN => n62907);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n56839, QN => n62908);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n56863, QN => n62909);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n56887, QN => n62910);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n56911, QN => n62911);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n56935, QN => n62912);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n56959, QN => n62913);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n56983, QN => n62914);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n57007, QN => n62915);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n57031, QN => n62916);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n57055, QN => n62917);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n57079, QN => n62918);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n57103, QN => n62919);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n57127, QN => n62920);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n57151, QN => n62921);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n57175, QN => n62922);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n57199, QN => n62923);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n57223, QN => n62924);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n57247, QN => n62925);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n57271, QN => n62926);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n57295, QN => n62927);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n57319, QN => n62928);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n57343, QN => n62929);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n57367, QN => n62930);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n57391, QN => n62931);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n57415, QN => n62932);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n57439, QN => n62933);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n57463, QN => n62934);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n57487, QN => n62935);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n57511, QN => n62936);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n57535, QN => n62937);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n57559, QN => n62938);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n57583, QN => n62939);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n57607, QN => n62940);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n57631, QN => n62941);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n58642, QN => n62942);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n58641, QN => n62943);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n58640, QN => n62944);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n58639, QN => n62945);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n58638, QN => n62946);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n58637, QN => n62947);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n58636, QN => n62948);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => 
                           n58635, QN => n62949);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => 
                           n58634, QN => n62950);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => 
                           n58633, QN => n62951);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => 
                           n58632, QN => n62952);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => 
                           n58631, QN => n62953);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => 
                           n58630, QN => n62954);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => 
                           n58629, QN => n62955);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => 
                           n58628, QN => n62956);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => 
                           n58627, QN => n62957);
   OUT1_reg_63_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => OUT1_63_port
                           , QN => n66554);
   OUT1_reg_62_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => OUT1_62_port
                           , QN => n66553);
   OUT1_reg_61_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => OUT1_61_port
                           , QN => n66552);
   OUT1_reg_60_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => OUT1_60_port
                           , QN => n66551);
   U45462 : NOR3_X1 port map( A1 => n67434, A2 => ADD_RD2(1), A3 => n66299, ZN 
                           => n66278);
   U45463 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n67434,
                           ZN => n66281);
   U45464 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n67632,
                           ZN => n65078);
   U45465 : NOR3_X1 port map( A1 => n67632, A2 => ADD_RD1(1), A3 => n65099, ZN 
                           => n65086);
   U45466 : AND3_X1 port map( A1 => ENABLE, A2 => n68057, A3 => RD1, ZN => 
                           n66494);
   U45467 : BUF_X1 port map( A => n67852, Z => n67854);
   U45468 : BUF_X1 port map( A => n68256, Z => n68258);
   U45469 : BUF_X1 port map( A => n67852, Z => n67855);
   U45470 : BUF_X1 port map( A => n67852, Z => n67856);
   U45471 : BUF_X1 port map( A => n67853, Z => n67857);
   U45472 : BUF_X1 port map( A => n67853, Z => n67858);
   U45473 : BUF_X1 port map( A => n68256, Z => n68259);
   U45474 : BUF_X1 port map( A => n68256, Z => n68260);
   U45475 : BUF_X1 port map( A => n68257, Z => n68261);
   U45476 : BUF_X1 port map( A => n68257, Z => n68262);
   U45477 : BUF_X1 port map( A => n61959, Z => n68251);
   U45478 : BUF_X1 port map( A => n61959, Z => n68252);
   U45479 : BUF_X1 port map( A => n61959, Z => n68253);
   U45480 : BUF_X1 port map( A => n61959, Z => n68254);
   U45481 : BUF_X1 port map( A => n65111, Z => n67440);
   U45482 : BUF_X1 port map( A => n65111, Z => n67441);
   U45483 : BUF_X1 port map( A => n65111, Z => n67442);
   U45484 : BUF_X1 port map( A => n65111, Z => n67443);
   U45485 : BUF_X1 port map( A => n65111, Z => n67444);
   U45486 : BUF_X1 port map( A => n67891, Z => n67893);
   U45487 : BUF_X1 port map( A => n67941, Z => n67943);
   U45488 : BUF_X1 port map( A => n67954, Z => n67956);
   U45489 : BUF_X1 port map( A => n68045, Z => n68047);
   U45490 : BUF_X1 port map( A => n68006, Z => n68008);
   U45491 : BUF_X1 port map( A => n67967, Z => n67969);
   U45492 : BUF_X1 port map( A => n67801, Z => n67803);
   U45493 : BUF_X1 port map( A => n67839, Z => n67841);
   U45494 : BUF_X1 port map( A => n67750, Z => n67752);
   U45495 : BUF_X1 port map( A => n67737, Z => n67739);
   U45496 : BUF_X1 port map( A => n67660, Z => n67662);
   U45497 : BUF_X1 port map( A => n67878, Z => n67880);
   U45498 : BUF_X1 port map( A => n68032, Z => n68034);
   U45499 : BUF_X1 port map( A => n68019, Z => n68021);
   U45500 : BUF_X1 port map( A => n67993, Z => n67995);
   U45501 : BUF_X1 port map( A => n67814, Z => n67816);
   U45502 : BUF_X1 port map( A => n67686, Z => n67688);
   U45503 : BUF_X1 port map( A => n67673, Z => n67675);
   U45504 : BUF_X1 port map( A => n67980, Z => n67982);
   U45505 : BUF_X1 port map( A => n67776, Z => n67778);
   U45506 : BUF_X1 port map( A => n67763, Z => n67765);
   U45507 : BUF_X1 port map( A => n67712, Z => n67714);
   U45508 : BUF_X1 port map( A => n67699, Z => n67701);
   U45509 : BUF_X1 port map( A => n67865, Z => n67867);
   U45510 : BUF_X1 port map( A => n67916, Z => n67918);
   U45511 : BUF_X1 port map( A => n67941, Z => n67944);
   U45512 : BUF_X1 port map( A => n67941, Z => n67945);
   U45513 : BUF_X1 port map( A => n67942, Z => n67946);
   U45514 : BUF_X1 port map( A => n67954, Z => n67957);
   U45515 : BUF_X1 port map( A => n67954, Z => n67958);
   U45516 : BUF_X1 port map( A => n67955, Z => n67959);
   U45517 : BUF_X1 port map( A => n68045, Z => n68048);
   U45518 : BUF_X1 port map( A => n68045, Z => n68049);
   U45519 : BUF_X1 port map( A => n68046, Z => n68050);
   U45520 : BUF_X1 port map( A => n68006, Z => n68009);
   U45521 : BUF_X1 port map( A => n68006, Z => n68010);
   U45522 : BUF_X1 port map( A => n68007, Z => n68011);
   U45523 : BUF_X1 port map( A => n67967, Z => n67970);
   U45524 : BUF_X1 port map( A => n67967, Z => n67971);
   U45525 : BUF_X1 port map( A => n67968, Z => n67972);
   U45526 : BUF_X1 port map( A => n67942, Z => n67947);
   U45527 : BUF_X1 port map( A => n67801, Z => n67804);
   U45528 : BUF_X1 port map( A => n67801, Z => n67805);
   U45529 : BUF_X1 port map( A => n67802, Z => n67806);
   U45530 : BUF_X1 port map( A => n67839, Z => n67842);
   U45531 : BUF_X1 port map( A => n67839, Z => n67843);
   U45532 : BUF_X1 port map( A => n67840, Z => n67844);
   U45533 : BUF_X1 port map( A => n67750, Z => n67753);
   U45534 : BUF_X1 port map( A => n67750, Z => n67754);
   U45535 : BUF_X1 port map( A => n67751, Z => n67755);
   U45536 : BUF_X1 port map( A => n67737, Z => n67740);
   U45537 : BUF_X1 port map( A => n67737, Z => n67741);
   U45538 : BUF_X1 port map( A => n67738, Z => n67742);
   U45539 : BUF_X1 port map( A => n67955, Z => n67960);
   U45540 : BUF_X1 port map( A => n68046, Z => n68051);
   U45541 : BUF_X1 port map( A => n68007, Z => n68012);
   U45542 : BUF_X1 port map( A => n67660, Z => n67663);
   U45543 : BUF_X1 port map( A => n67660, Z => n67664);
   U45544 : BUF_X1 port map( A => n67661, Z => n67665);
   U45545 : BUF_X1 port map( A => n67968, Z => n67973);
   U45546 : BUF_X1 port map( A => n67802, Z => n67807);
   U45547 : BUF_X1 port map( A => n67840, Z => n67845);
   U45548 : BUF_X1 port map( A => n67751, Z => n67756);
   U45549 : BUF_X1 port map( A => n67738, Z => n67743);
   U45550 : BUF_X1 port map( A => n67661, Z => n67666);
   U45551 : BUF_X1 port map( A => n67878, Z => n67881);
   U45552 : BUF_X1 port map( A => n67878, Z => n67882);
   U45553 : BUF_X1 port map( A => n67879, Z => n67883);
   U45554 : BUF_X1 port map( A => n68032, Z => n68035);
   U45555 : BUF_X1 port map( A => n68032, Z => n68036);
   U45556 : BUF_X1 port map( A => n68033, Z => n68037);
   U45557 : BUF_X1 port map( A => n68019, Z => n68022);
   U45558 : BUF_X1 port map( A => n68019, Z => n68023);
   U45559 : BUF_X1 port map( A => n68020, Z => n68024);
   U45560 : BUF_X1 port map( A => n67993, Z => n67996);
   U45561 : BUF_X1 port map( A => n67993, Z => n67997);
   U45562 : BUF_X1 port map( A => n67994, Z => n67998);
   U45563 : BUF_X1 port map( A => n67814, Z => n67817);
   U45564 : BUF_X1 port map( A => n67814, Z => n67818);
   U45565 : BUF_X1 port map( A => n67815, Z => n67819);
   U45566 : BUF_X1 port map( A => n67686, Z => n67689);
   U45567 : BUF_X1 port map( A => n67686, Z => n67690);
   U45568 : BUF_X1 port map( A => n67687, Z => n67691);
   U45569 : BUF_X1 port map( A => n67673, Z => n67676);
   U45570 : BUF_X1 port map( A => n67673, Z => n67677);
   U45571 : BUF_X1 port map( A => n67674, Z => n67678);
   U45572 : BUF_X1 port map( A => n67879, Z => n67884);
   U45573 : BUF_X1 port map( A => n68033, Z => n68038);
   U45574 : BUF_X1 port map( A => n68020, Z => n68025);
   U45575 : BUF_X1 port map( A => n67994, Z => n67999);
   U45576 : BUF_X1 port map( A => n67815, Z => n67820);
   U45577 : BUF_X1 port map( A => n67687, Z => n67692);
   U45578 : BUF_X1 port map( A => n67674, Z => n67679);
   U45579 : BUF_X1 port map( A => n67980, Z => n67983);
   U45580 : BUF_X1 port map( A => n67980, Z => n67984);
   U45581 : BUF_X1 port map( A => n67981, Z => n67985);
   U45582 : BUF_X1 port map( A => n67776, Z => n67779);
   U45583 : BUF_X1 port map( A => n67776, Z => n67780);
   U45584 : BUF_X1 port map( A => n67777, Z => n67781);
   U45585 : BUF_X1 port map( A => n67763, Z => n67766);
   U45586 : BUF_X1 port map( A => n67763, Z => n67767);
   U45587 : BUF_X1 port map( A => n67764, Z => n67768);
   U45588 : BUF_X1 port map( A => n67712, Z => n67715);
   U45589 : BUF_X1 port map( A => n67712, Z => n67716);
   U45590 : BUF_X1 port map( A => n67713, Z => n67717);
   U45591 : BUF_X1 port map( A => n67699, Z => n67702);
   U45592 : BUF_X1 port map( A => n67699, Z => n67703);
   U45593 : BUF_X1 port map( A => n67700, Z => n67704);
   U45594 : BUF_X1 port map( A => n67981, Z => n67986);
   U45595 : BUF_X1 port map( A => n67777, Z => n67782);
   U45596 : BUF_X1 port map( A => n67764, Z => n67769);
   U45597 : BUF_X1 port map( A => n67713, Z => n67718);
   U45598 : BUF_X1 port map( A => n67700, Z => n67705);
   U45599 : BUF_X1 port map( A => n67865, Z => n67868);
   U45600 : BUF_X1 port map( A => n67865, Z => n67869);
   U45601 : BUF_X1 port map( A => n67866, Z => n67870);
   U45602 : BUF_X1 port map( A => n67866, Z => n67871);
   U45603 : BUF_X1 port map( A => n67892, Z => n67897);
   U45604 : BUF_X1 port map( A => n67892, Z => n67896);
   U45605 : BUF_X1 port map( A => n67891, Z => n67895);
   U45606 : BUF_X1 port map( A => n67891, Z => n67894);
   U45607 : BUF_X1 port map( A => n67916, Z => n67919);
   U45608 : BUF_X1 port map( A => n67916, Z => n67920);
   U45609 : BUF_X1 port map( A => n67917, Z => n67921);
   U45610 : BUF_X1 port map( A => n67917, Z => n67922);
   U45611 : BUF_X1 port map( A => n62092, Z => n68039);
   U45612 : BUF_X1 port map( A => n62092, Z => n68040);
   U45613 : BUF_X1 port map( A => n62092, Z => n68041);
   U45614 : BUF_X1 port map( A => n62092, Z => n68042);
   U45615 : BUF_X1 port map( A => n62092, Z => n68043);
   U45616 : BUF_X1 port map( A => n63766, Z => n67654);
   U45617 : BUF_X1 port map( A => n63766, Z => n67655);
   U45618 : BUF_X1 port map( A => n63766, Z => n67656);
   U45619 : BUF_X1 port map( A => n63766, Z => n67657);
   U45620 : BUF_X1 port map( A => n63766, Z => n67658);
   U45621 : BUF_X1 port map( A => n62159, Z => n68026);
   U45622 : BUF_X1 port map( A => n62159, Z => n68027);
   U45623 : BUF_X1 port map( A => n62159, Z => n68028);
   U45624 : BUF_X1 port map( A => n62159, Z => n68029);
   U45625 : BUF_X1 port map( A => n62159, Z => n68030);
   U45626 : BUF_X1 port map( A => n62628, Z => n67935);
   U45627 : BUF_X1 port map( A => n62628, Z => n67936);
   U45628 : BUF_X1 port map( A => n62628, Z => n67937);
   U45629 : BUF_X1 port map( A => n62628, Z => n67938);
   U45630 : BUF_X1 port map( A => n62628, Z => n67939);
   U45631 : BUF_X1 port map( A => n62561, Z => n67948);
   U45632 : BUF_X1 port map( A => n62561, Z => n67949);
   U45633 : BUF_X1 port map( A => n62561, Z => n67950);
   U45634 : BUF_X1 port map( A => n62561, Z => n67951);
   U45635 : BUF_X1 port map( A => n62561, Z => n67952);
   U45636 : BUF_X1 port map( A => n62695, Z => n67923);
   U45637 : BUF_X1 port map( A => n62695, Z => n67924);
   U45638 : BUF_X1 port map( A => n62695, Z => n67925);
   U45639 : BUF_X1 port map( A => n62695, Z => n67926);
   U45640 : BUF_X1 port map( A => n62695, Z => n67927);
   U45641 : BUF_X1 port map( A => n62292, Z => n68000);
   U45642 : BUF_X1 port map( A => n62292, Z => n68001);
   U45643 : BUF_X1 port map( A => n62292, Z => n68002);
   U45644 : BUF_X1 port map( A => n62292, Z => n68003);
   U45645 : BUF_X1 port map( A => n62292, Z => n68004);
   U45646 : BUF_X1 port map( A => n62495, Z => n67961);
   U45647 : BUF_X1 port map( A => n62495, Z => n67962);
   U45648 : BUF_X1 port map( A => n62495, Z => n67963);
   U45649 : BUF_X1 port map( A => n62495, Z => n67964);
   U45650 : BUF_X1 port map( A => n62495, Z => n67965);
   U45651 : BUF_X1 port map( A => n63163, Z => n67795);
   U45652 : BUF_X1 port map( A => n63163, Z => n67796);
   U45653 : BUF_X1 port map( A => n63163, Z => n67797);
   U45654 : BUF_X1 port map( A => n63163, Z => n67798);
   U45655 : BUF_X1 port map( A => n63163, Z => n67799);
   U45656 : BUF_X1 port map( A => n62961, Z => n67846);
   U45657 : BUF_X1 port map( A => n62961, Z => n67847);
   U45658 : BUF_X1 port map( A => n62961, Z => n67848);
   U45659 : BUF_X1 port map( A => n62961, Z => n67849);
   U45660 : BUF_X1 port map( A => n62961, Z => n67850);
   U45661 : BUF_X1 port map( A => n63028, Z => n67833);
   U45662 : BUF_X1 port map( A => n63028, Z => n67834);
   U45663 : BUF_X1 port map( A => n63028, Z => n67835);
   U45664 : BUF_X1 port map( A => n63028, Z => n67836);
   U45665 : BUF_X1 port map( A => n63028, Z => n67837);
   U45666 : BUF_X1 port map( A => n63364, Z => n67744);
   U45667 : BUF_X1 port map( A => n63364, Z => n67745);
   U45668 : BUF_X1 port map( A => n63364, Z => n67746);
   U45669 : BUF_X1 port map( A => n63364, Z => n67747);
   U45670 : BUF_X1 port map( A => n63364, Z => n67748);
   U45671 : BUF_X1 port map( A => n63431, Z => n67731);
   U45672 : BUF_X1 port map( A => n63431, Z => n67732);
   U45673 : BUF_X1 port map( A => n63431, Z => n67733);
   U45674 : BUF_X1 port map( A => n63431, Z => n67734);
   U45675 : BUF_X1 port map( A => n63431, Z => n67735);
   U45676 : BUF_X1 port map( A => n63499, Z => n67719);
   U45677 : BUF_X1 port map( A => n63499, Z => n67720);
   U45678 : BUF_X1 port map( A => n63499, Z => n67721);
   U45679 : BUF_X1 port map( A => n63499, Z => n67722);
   U45680 : BUF_X1 port map( A => n63499, Z => n67723);
   U45681 : BUF_X1 port map( A => n62763, Z => n67898);
   U45682 : BUF_X1 port map( A => n62763, Z => n67899);
   U45683 : BUF_X1 port map( A => n62763, Z => n67900);
   U45684 : BUF_X1 port map( A => n62763, Z => n67901);
   U45685 : BUF_X1 port map( A => n62763, Z => n67902);
   U45686 : BUF_X1 port map( A => n62828, Z => n67872);
   U45687 : BUF_X1 port map( A => n62828, Z => n67873);
   U45688 : BUF_X1 port map( A => n62828, Z => n67874);
   U45689 : BUF_X1 port map( A => n62828, Z => n67875);
   U45690 : BUF_X1 port map( A => n62828, Z => n67876);
   U45691 : BUF_X1 port map( A => n62226, Z => n68013);
   U45692 : BUF_X1 port map( A => n62226, Z => n68014);
   U45693 : BUF_X1 port map( A => n62226, Z => n68015);
   U45694 : BUF_X1 port map( A => n62226, Z => n68016);
   U45695 : BUF_X1 port map( A => n62226, Z => n68017);
   U45696 : BUF_X1 port map( A => n62359, Z => n67987);
   U45697 : BUF_X1 port map( A => n62359, Z => n67988);
   U45698 : BUF_X1 port map( A => n62359, Z => n67989);
   U45699 : BUF_X1 port map( A => n62359, Z => n67990);
   U45700 : BUF_X1 port map( A => n62359, Z => n67991);
   U45701 : BUF_X1 port map( A => n63097, Z => n67808);
   U45702 : BUF_X1 port map( A => n63097, Z => n67809);
   U45703 : BUF_X1 port map( A => n63097, Z => n67810);
   U45704 : BUF_X1 port map( A => n63097, Z => n67811);
   U45705 : BUF_X1 port map( A => n63097, Z => n67812);
   U45706 : BUF_X1 port map( A => n63634, Z => n67680);
   U45707 : BUF_X1 port map( A => n63634, Z => n67681);
   U45708 : BUF_X1 port map( A => n63634, Z => n67682);
   U45709 : BUF_X1 port map( A => n63634, Z => n67683);
   U45710 : BUF_X1 port map( A => n63634, Z => n67684);
   U45711 : BUF_X1 port map( A => n63700, Z => n67667);
   U45712 : BUF_X1 port map( A => n63700, Z => n67668);
   U45713 : BUF_X1 port map( A => n63700, Z => n67669);
   U45714 : BUF_X1 port map( A => n63700, Z => n67670);
   U45715 : BUF_X1 port map( A => n63700, Z => n67671);
   U45716 : BUF_X1 port map( A => n62425, Z => n67974);
   U45717 : BUF_X1 port map( A => n62425, Z => n67975);
   U45718 : BUF_X1 port map( A => n62425, Z => n67976);
   U45719 : BUF_X1 port map( A => n62425, Z => n67977);
   U45720 : BUF_X1 port map( A => n62425, Z => n67978);
   U45721 : BUF_X1 port map( A => n63094, Z => n67821);
   U45722 : BUF_X1 port map( A => n63094, Z => n67822);
   U45723 : BUF_X1 port map( A => n63094, Z => n67823);
   U45724 : BUF_X1 port map( A => n63094, Z => n67824);
   U45725 : BUF_X1 port map( A => n63094, Z => n67825);
   U45726 : BUF_X1 port map( A => n63231, Z => n67770);
   U45727 : BUF_X1 port map( A => n63231, Z => n67771);
   U45728 : BUF_X1 port map( A => n63231, Z => n67772);
   U45729 : BUF_X1 port map( A => n63231, Z => n67773);
   U45730 : BUF_X1 port map( A => n63231, Z => n67774);
   U45731 : BUF_X1 port map( A => n63228, Z => n67783);
   U45732 : BUF_X1 port map( A => n63228, Z => n67784);
   U45733 : BUF_X1 port map( A => n63228, Z => n67785);
   U45734 : BUF_X1 port map( A => n63228, Z => n67786);
   U45735 : BUF_X1 port map( A => n63228, Z => n67787);
   U45736 : BUF_X1 port map( A => n63298, Z => n67757);
   U45737 : BUF_X1 port map( A => n63298, Z => n67758);
   U45738 : BUF_X1 port map( A => n63298, Z => n67759);
   U45739 : BUF_X1 port map( A => n63298, Z => n67760);
   U45740 : BUF_X1 port map( A => n63298, Z => n67761);
   U45741 : BUF_X1 port map( A => n63502, Z => n67706);
   U45742 : BUF_X1 port map( A => n63502, Z => n67707);
   U45743 : BUF_X1 port map( A => n63502, Z => n67708);
   U45744 : BUF_X1 port map( A => n63502, Z => n67709);
   U45745 : BUF_X1 port map( A => n63502, Z => n67710);
   U45746 : BUF_X1 port map( A => n63568, Z => n67693);
   U45747 : BUF_X1 port map( A => n63568, Z => n67694);
   U45748 : BUF_X1 port map( A => n63568, Z => n67695);
   U45749 : BUF_X1 port map( A => n63568, Z => n67696);
   U45750 : BUF_X1 port map( A => n63568, Z => n67697);
   U45751 : BUF_X1 port map( A => n62894, Z => n67859);
   U45752 : BUF_X1 port map( A => n62894, Z => n67860);
   U45753 : BUF_X1 port map( A => n62894, Z => n67861);
   U45754 : BUF_X1 port map( A => n62894, Z => n67862);
   U45755 : BUF_X1 port map( A => n62894, Z => n67863);
   U45756 : BUF_X1 port map( A => n62765, Z => n67885);
   U45757 : BUF_X1 port map( A => n62765, Z => n67886);
   U45758 : BUF_X1 port map( A => n62765, Z => n67887);
   U45759 : BUF_X1 port map( A => n62765, Z => n67888);
   U45760 : BUF_X1 port map( A => n62765, Z => n67889);
   U45761 : BUF_X1 port map( A => n62698, Z => n67910);
   U45762 : BUF_X1 port map( A => n62698, Z => n67911);
   U45763 : BUF_X1 port map( A => n62698, Z => n67912);
   U45764 : BUF_X1 port map( A => n62698, Z => n67913);
   U45765 : BUF_X1 port map( A => n62698, Z => n67914);
   U45766 : BUF_X1 port map( A => n61959, Z => n68250);
   U45767 : BUF_X1 port map( A => n61957, Z => n68256);
   U45768 : BUF_X1 port map( A => n62959, Z => n67852);
   U45769 : BUF_X1 port map( A => n61957, Z => n68257);
   U45770 : BUF_X1 port map( A => n62959, Z => n67853);
   U45771 : INV_X1 port map( A => n66494, ZN => n67632);
   U45772 : INV_X1 port map( A => n66494, ZN => n67633);
   U45773 : INV_X1 port map( A => n66494, ZN => n67634);
   U45774 : INV_X1 port map( A => n66494, ZN => n67635);
   U45775 : BUF_X1 port map( A => n63790, Z => n67588);
   U45776 : BUF_X1 port map( A => n65146, Z => n67278);
   U45777 : BUF_X1 port map( A => n65146, Z => n67279);
   U45778 : BUF_X1 port map( A => n65146, Z => n67280);
   U45779 : BUF_X1 port map( A => n65146, Z => n67281);
   U45780 : BUF_X1 port map( A => n65146, Z => n67282);
   U45781 : BUF_X1 port map( A => n65141, Z => n67302);
   U45782 : BUF_X1 port map( A => n65141, Z => n67303);
   U45783 : BUF_X1 port map( A => n65141, Z => n67304);
   U45784 : BUF_X1 port map( A => n65141, Z => n67305);
   U45785 : BUF_X1 port map( A => n65141, Z => n67306);
   U45786 : BUF_X1 port map( A => n63815, Z => n67476);
   U45787 : BUF_X1 port map( A => n63815, Z => n67477);
   U45788 : BUF_X1 port map( A => n63815, Z => n67478);
   U45789 : BUF_X1 port map( A => n63815, Z => n67479);
   U45790 : BUF_X1 port map( A => n63815, Z => n67480);
   U45791 : BUF_X1 port map( A => n63810, Z => n67500);
   U45792 : BUF_X1 port map( A => n63810, Z => n67501);
   U45793 : BUF_X1 port map( A => n63810, Z => n67502);
   U45794 : BUF_X1 port map( A => n63810, Z => n67503);
   U45795 : BUF_X1 port map( A => n63810, Z => n67504);
   U45796 : BUF_X1 port map( A => n65116, Z => n67416);
   U45797 : BUF_X1 port map( A => n65121, Z => n67392);
   U45798 : BUF_X1 port map( A => n65126, Z => n67368);
   U45799 : BUF_X1 port map( A => n65116, Z => n67417);
   U45800 : BUF_X1 port map( A => n65121, Z => n67393);
   U45801 : BUF_X1 port map( A => n65126, Z => n67369);
   U45802 : BUF_X1 port map( A => n65116, Z => n67418);
   U45803 : BUF_X1 port map( A => n65121, Z => n67394);
   U45804 : BUF_X1 port map( A => n65126, Z => n67370);
   U45805 : BUF_X1 port map( A => n65116, Z => n67419);
   U45806 : BUF_X1 port map( A => n65121, Z => n67395);
   U45807 : BUF_X1 port map( A => n65126, Z => n67371);
   U45808 : BUF_X1 port map( A => n65116, Z => n67420);
   U45809 : BUF_X1 port map( A => n65121, Z => n67396);
   U45810 : BUF_X1 port map( A => n65126, Z => n67372);
   U45811 : BUF_X1 port map( A => n63794, Z => n67566);
   U45812 : BUF_X1 port map( A => n63788, Z => n67590);
   U45813 : BUF_X1 port map( A => n63794, Z => n67567);
   U45814 : BUF_X1 port map( A => n63788, Z => n67591);
   U45815 : BUF_X1 port map( A => n63794, Z => n67568);
   U45816 : BUF_X1 port map( A => n63788, Z => n67592);
   U45817 : BUF_X1 port map( A => n63794, Z => n67569);
   U45818 : BUF_X1 port map( A => n63788, Z => n67593);
   U45819 : BUF_X1 port map( A => n63794, Z => n67570);
   U45820 : BUF_X1 port map( A => n63788, Z => n67594);
   U45821 : BUF_X1 port map( A => n63778, Z => n67636);
   U45822 : BUF_X1 port map( A => n63783, Z => n67614);
   U45823 : BUF_X1 port map( A => n63778, Z => n67637);
   U45824 : BUF_X1 port map( A => n63783, Z => n67615);
   U45825 : BUF_X1 port map( A => n63778, Z => n67638);
   U45826 : BUF_X1 port map( A => n63783, Z => n67616);
   U45827 : BUF_X1 port map( A => n63778, Z => n67639);
   U45828 : BUF_X1 port map( A => n63783, Z => n67617);
   U45829 : BUF_X1 port map( A => n63778, Z => n67640);
   U45830 : BUF_X1 port map( A => n63783, Z => n67618);
   U45831 : BUF_X1 port map( A => n65142, Z => n67296);
   U45832 : BUF_X1 port map( A => n65147, Z => n67272);
   U45833 : BUF_X1 port map( A => n65142, Z => n67297);
   U45834 : BUF_X1 port map( A => n65147, Z => n67273);
   U45835 : BUF_X1 port map( A => n65142, Z => n67298);
   U45836 : BUF_X1 port map( A => n65147, Z => n67274);
   U45837 : BUF_X1 port map( A => n65142, Z => n67299);
   U45838 : BUF_X1 port map( A => n65147, Z => n67275);
   U45839 : BUF_X1 port map( A => n65142, Z => n67300);
   U45840 : BUF_X1 port map( A => n65147, Z => n67276);
   U45841 : BUF_X1 port map( A => n63811, Z => n67494);
   U45842 : BUF_X1 port map( A => n63816, Z => n67470);
   U45843 : BUF_X1 port map( A => n63811, Z => n67495);
   U45844 : BUF_X1 port map( A => n63816, Z => n67471);
   U45845 : BUF_X1 port map( A => n63811, Z => n67496);
   U45846 : BUF_X1 port map( A => n63816, Z => n67472);
   U45847 : BUF_X1 port map( A => n63811, Z => n67497);
   U45848 : BUF_X1 port map( A => n63816, Z => n67473);
   U45849 : BUF_X1 port map( A => n63811, Z => n67498);
   U45850 : BUF_X1 port map( A => n63816, Z => n67474);
   U45851 : BUF_X1 port map( A => n65113, Z => n67429);
   U45852 : BUF_X1 port map( A => n65113, Z => n67430);
   U45853 : BUF_X1 port map( A => n65113, Z => n67431);
   U45854 : BUF_X1 port map( A => n65113, Z => n67432);
   U45855 : BUF_X1 port map( A => n65108, Z => n67453);
   U45856 : BUF_X1 port map( A => n65118, Z => n67405);
   U45857 : BUF_X1 port map( A => n65123, Z => n67381);
   U45858 : BUF_X1 port map( A => n65108, Z => n67454);
   U45859 : BUF_X1 port map( A => n65118, Z => n67406);
   U45860 : BUF_X1 port map( A => n65123, Z => n67382);
   U45861 : BUF_X1 port map( A => n65108, Z => n67455);
   U45862 : BUF_X1 port map( A => n65118, Z => n67407);
   U45863 : BUF_X1 port map( A => n65123, Z => n67383);
   U45864 : BUF_X1 port map( A => n65108, Z => n67456);
   U45865 : BUF_X1 port map( A => n65118, Z => n67408);
   U45866 : BUF_X1 port map( A => n65123, Z => n67384);
   U45867 : BUF_X1 port map( A => n63775, Z => n67649);
   U45868 : BUF_X1 port map( A => n63775, Z => n67650);
   U45869 : BUF_X1 port map( A => n63775, Z => n67651);
   U45870 : BUF_X1 port map( A => n63775, Z => n67652);
   U45871 : BUF_X1 port map( A => n63791, Z => n67579);
   U45872 : BUF_X1 port map( A => n63785, Z => n67603);
   U45873 : BUF_X1 port map( A => n63780, Z => n67627);
   U45874 : BUF_X1 port map( A => n63791, Z => n67580);
   U45875 : BUF_X1 port map( A => n63785, Z => n67604);
   U45876 : BUF_X1 port map( A => n63780, Z => n67628);
   U45877 : BUF_X1 port map( A => n63791, Z => n67581);
   U45878 : BUF_X1 port map( A => n63785, Z => n67605);
   U45879 : BUF_X1 port map( A => n63780, Z => n67629);
   U45880 : BUF_X1 port map( A => n63791, Z => n67582);
   U45881 : BUF_X1 port map( A => n63785, Z => n67606);
   U45882 : BUF_X1 port map( A => n63780, Z => n67630);
   U45883 : BUF_X1 port map( A => n65140, Z => n67308);
   U45884 : BUF_X1 port map( A => n65140, Z => n67309);
   U45885 : BUF_X1 port map( A => n65140, Z => n67310);
   U45886 : BUF_X1 port map( A => n65140, Z => n67311);
   U45887 : BUF_X1 port map( A => n65140, Z => n67312);
   U45888 : BUF_X1 port map( A => n63809, Z => n67506);
   U45889 : BUF_X1 port map( A => n63809, Z => n67507);
   U45890 : BUF_X1 port map( A => n63809, Z => n67508);
   U45891 : BUF_X1 port map( A => n63809, Z => n67509);
   U45892 : BUF_X1 port map( A => n63809, Z => n67510);
   U45893 : BUF_X1 port map( A => n63807, Z => n67518);
   U45894 : BUF_X1 port map( A => n63807, Z => n67519);
   U45895 : BUF_X1 port map( A => n63807, Z => n67520);
   U45896 : BUF_X1 port map( A => n63807, Z => n67521);
   U45897 : BUF_X1 port map( A => n63807, Z => n67522);
   U45898 : BUF_X1 port map( A => n65138, Z => n67320);
   U45899 : BUF_X1 port map( A => n65138, Z => n67321);
   U45900 : BUF_X1 port map( A => n65138, Z => n67322);
   U45901 : BUF_X1 port map( A => n65138, Z => n67323);
   U45902 : BUF_X1 port map( A => n65138, Z => n67324);
   U45903 : BUF_X1 port map( A => n65139, Z => n67314);
   U45904 : BUF_X1 port map( A => n65139, Z => n67315);
   U45905 : BUF_X1 port map( A => n65139, Z => n67316);
   U45906 : BUF_X1 port map( A => n65139, Z => n67317);
   U45907 : BUF_X1 port map( A => n65139, Z => n67318);
   U45908 : BUF_X1 port map( A => n63808, Z => n67512);
   U45909 : BUF_X1 port map( A => n63808, Z => n67513);
   U45910 : BUF_X1 port map( A => n63808, Z => n67514);
   U45911 : BUF_X1 port map( A => n63808, Z => n67515);
   U45912 : BUF_X1 port map( A => n63808, Z => n67516);
   U45913 : BUF_X1 port map( A => n65117, Z => n67410);
   U45914 : BUF_X1 port map( A => n65117, Z => n67411);
   U45915 : BUF_X1 port map( A => n65117, Z => n67412);
   U45916 : BUF_X1 port map( A => n65117, Z => n67413);
   U45917 : BUF_X1 port map( A => n65117, Z => n67414);
   U45918 : BUF_X1 port map( A => n65122, Z => n67386);
   U45919 : BUF_X1 port map( A => n65127, Z => n67362);
   U45920 : BUF_X1 port map( A => n65122, Z => n67387);
   U45921 : BUF_X1 port map( A => n65127, Z => n67363);
   U45922 : BUF_X1 port map( A => n65122, Z => n67388);
   U45923 : BUF_X1 port map( A => n65127, Z => n67364);
   U45924 : BUF_X1 port map( A => n65122, Z => n67389);
   U45925 : BUF_X1 port map( A => n65127, Z => n67365);
   U45926 : BUF_X1 port map( A => n65122, Z => n67390);
   U45927 : BUF_X1 port map( A => n65127, Z => n67366);
   U45928 : BUF_X1 port map( A => n63795, Z => n67560);
   U45929 : BUF_X1 port map( A => n63795, Z => n67561);
   U45930 : BUF_X1 port map( A => n63795, Z => n67562);
   U45931 : BUF_X1 port map( A => n63795, Z => n67563);
   U45932 : BUF_X1 port map( A => n63795, Z => n67564);
   U45933 : BUF_X1 port map( A => n63784, Z => n67608);
   U45934 : BUF_X1 port map( A => n63784, Z => n67609);
   U45935 : BUF_X1 port map( A => n63784, Z => n67610);
   U45936 : BUF_X1 port map( A => n63784, Z => n67611);
   U45937 : BUF_X1 port map( A => n63784, Z => n67612);
   U45938 : NAND2_X1 port map( A1 => n68057, A2 => n68047, ZN => n62092);
   U45939 : NAND2_X1 port map( A1 => n68057, A2 => n67662, ZN => n63766);
   U45940 : NAND2_X1 port map( A1 => n68057, A2 => n68034, ZN => n62159);
   U45941 : BUF_X1 port map( A => n63790, Z => n67584);
   U45942 : BUF_X1 port map( A => n63790, Z => n67585);
   U45943 : BUF_X1 port map( A => n63790, Z => n67586);
   U45944 : BUF_X1 port map( A => n63790, Z => n67587);
   U45945 : BUF_X1 port map( A => n62693, Z => n67929);
   U45946 : BUF_X1 port map( A => n63498, Z => n67725);
   U45947 : BUF_X1 port map( A => n62762, Z => n67904);
   U45948 : BUF_X1 port map( A => n63093, Z => n67827);
   U45949 : BUF_X1 port map( A => n63227, Z => n67789);
   U45950 : BUF_X1 port map( A => n62693, Z => n67930);
   U45951 : BUF_X1 port map( A => n62693, Z => n67931);
   U45952 : BUF_X1 port map( A => n62693, Z => n67932);
   U45953 : BUF_X1 port map( A => n62693, Z => n67933);
   U45954 : BUF_X1 port map( A => n63498, Z => n67726);
   U45955 : BUF_X1 port map( A => n63498, Z => n67727);
   U45956 : BUF_X1 port map( A => n63498, Z => n67728);
   U45957 : BUF_X1 port map( A => n63498, Z => n67729);
   U45958 : BUF_X1 port map( A => n62762, Z => n67905);
   U45959 : BUF_X1 port map( A => n62762, Z => n67906);
   U45960 : BUF_X1 port map( A => n62762, Z => n67907);
   U45961 : BUF_X1 port map( A => n62762, Z => n67908);
   U45962 : BUF_X1 port map( A => n63093, Z => n67828);
   U45963 : BUF_X1 port map( A => n63093, Z => n67829);
   U45964 : BUF_X1 port map( A => n63093, Z => n67830);
   U45965 : BUF_X1 port map( A => n63093, Z => n67831);
   U45966 : BUF_X1 port map( A => n63227, Z => n67790);
   U45967 : BUF_X1 port map( A => n63227, Z => n67791);
   U45968 : BUF_X1 port map( A => n63227, Z => n67792);
   U45969 : BUF_X1 port map( A => n63227, Z => n67793);
   U45970 : BUF_X1 port map( A => n65132, Z => n67356);
   U45971 : BUF_X1 port map( A => n65134, Z => n67344);
   U45972 : BUF_X1 port map( A => n65132, Z => n67357);
   U45973 : BUF_X1 port map( A => n65134, Z => n67345);
   U45974 : BUF_X1 port map( A => n65132, Z => n67358);
   U45975 : BUF_X1 port map( A => n65134, Z => n67346);
   U45976 : BUF_X1 port map( A => n65132, Z => n67359);
   U45977 : BUF_X1 port map( A => n65134, Z => n67347);
   U45978 : BUF_X1 port map( A => n65132, Z => n67360);
   U45979 : BUF_X1 port map( A => n65134, Z => n67348);
   U45980 : BUF_X1 port map( A => n65144, Z => n67290);
   U45981 : BUF_X1 port map( A => n65149, Z => n67266);
   U45982 : BUF_X1 port map( A => n65144, Z => n67291);
   U45983 : BUF_X1 port map( A => n65149, Z => n67267);
   U45984 : BUF_X1 port map( A => n65144, Z => n67292);
   U45985 : BUF_X1 port map( A => n65149, Z => n67268);
   U45986 : BUF_X1 port map( A => n65144, Z => n67293);
   U45987 : BUF_X1 port map( A => n65149, Z => n67269);
   U45988 : BUF_X1 port map( A => n65144, Z => n67294);
   U45989 : BUF_X1 port map( A => n65149, Z => n67270);
   U45990 : BUF_X1 port map( A => n63805, Z => n67530);
   U45991 : BUF_X1 port map( A => n63801, Z => n67554);
   U45992 : BUF_X1 port map( A => n63803, Z => n67542);
   U45993 : BUF_X1 port map( A => n63805, Z => n67531);
   U45994 : BUF_X1 port map( A => n63801, Z => n67555);
   U45995 : BUF_X1 port map( A => n63803, Z => n67543);
   U45996 : BUF_X1 port map( A => n63805, Z => n67532);
   U45997 : BUF_X1 port map( A => n63801, Z => n67556);
   U45998 : BUF_X1 port map( A => n63803, Z => n67544);
   U45999 : BUF_X1 port map( A => n63805, Z => n67533);
   U46000 : BUF_X1 port map( A => n63801, Z => n67557);
   U46001 : BUF_X1 port map( A => n63803, Z => n67545);
   U46002 : BUF_X1 port map( A => n63805, Z => n67534);
   U46003 : BUF_X1 port map( A => n63801, Z => n67558);
   U46004 : BUF_X1 port map( A => n63803, Z => n67546);
   U46005 : BUF_X1 port map( A => n63818, Z => n67464);
   U46006 : BUF_X1 port map( A => n63818, Z => n67465);
   U46007 : BUF_X1 port map( A => n63818, Z => n67466);
   U46008 : BUF_X1 port map( A => n63818, Z => n67467);
   U46009 : BUF_X1 port map( A => n63818, Z => n67468);
   U46010 : BUF_X1 port map( A => n65136, Z => n67332);
   U46011 : BUF_X1 port map( A => n65136, Z => n67333);
   U46012 : BUF_X1 port map( A => n65136, Z => n67334);
   U46013 : BUF_X1 port map( A => n65136, Z => n67335);
   U46014 : BUF_X1 port map( A => n65136, Z => n67336);
   U46015 : BUF_X1 port map( A => n63813, Z => n67488);
   U46016 : BUF_X1 port map( A => n63813, Z => n67489);
   U46017 : BUF_X1 port map( A => n63813, Z => n67490);
   U46018 : BUF_X1 port map( A => n63813, Z => n67491);
   U46019 : BUF_X1 port map( A => n63813, Z => n67492);
   U46020 : NAND2_X1 port map( A1 => n68054, A2 => n67803, ZN => n63163);
   U46021 : NAND2_X1 port map( A1 => n68054, A2 => n67827, ZN => n63094);
   U46022 : NAND2_X1 port map( A1 => n68054, A2 => n67778, ZN => n63231);
   U46023 : NAND2_X1 port map( A1 => n68054, A2 => n67789, ZN => n63228);
   U46024 : NAND2_X1 port map( A1 => n68056, A2 => n67943, ZN => n62628);
   U46025 : NAND2_X1 port map( A1 => n68056, A2 => n67956, ZN => n62561);
   U46026 : NAND2_X1 port map( A1 => n68056, A2 => n68008, ZN => n62292);
   U46027 : NAND2_X1 port map( A1 => n68056, A2 => n67969, ZN => n62495);
   U46028 : NAND2_X1 port map( A1 => n68055, A2 => n67854, ZN => n62961);
   U46029 : NAND2_X1 port map( A1 => n68055, A2 => n67841, ZN => n63028);
   U46030 : NAND2_X1 port map( A1 => n68055, A2 => n67752, ZN => n63364);
   U46031 : NAND2_X1 port map( A1 => n68056, A2 => n67739, ZN => n63431);
   U46032 : NAND2_X1 port map( A1 => n68055, A2 => n67725, ZN => n63499);
   U46033 : NAND2_X1 port map( A1 => n68055, A2 => n67904, ZN => n62763);
   U46034 : NAND2_X1 port map( A1 => n68055, A2 => n67880, ZN => n62828);
   U46035 : NAND2_X1 port map( A1 => n68056, A2 => n68021, ZN => n62226);
   U46036 : NAND2_X1 port map( A1 => n68056, A2 => n67995, ZN => n62359);
   U46037 : NAND2_X1 port map( A1 => n68055, A2 => n67816, ZN => n63097);
   U46038 : NAND2_X1 port map( A1 => n68056, A2 => n67688, ZN => n63634);
   U46039 : NAND2_X1 port map( A1 => n68056, A2 => n67675, ZN => n63700);
   U46040 : NAND2_X1 port map( A1 => n68055, A2 => n67929, ZN => n62695);
   U46041 : NAND2_X1 port map( A1 => n68056, A2 => n67982, ZN => n62425);
   U46042 : NAND2_X1 port map( A1 => n68055, A2 => n67765, ZN => n63298);
   U46043 : NAND2_X1 port map( A1 => n68056, A2 => n67714, ZN => n63502);
   U46044 : NAND2_X1 port map( A1 => n68056, A2 => n67701, ZN => n63568);
   U46045 : NAND2_X1 port map( A1 => n68055, A2 => n67867, ZN => n62894);
   U46046 : NAND2_X1 port map( A1 => n68055, A2 => n67893, ZN => n62765);
   U46047 : NAND2_X1 port map( A1 => n68055, A2 => n67918, ZN => n62698);
   U46048 : BUF_X1 port map( A => n65145, Z => n67284);
   U46049 : BUF_X1 port map( A => n65133, Z => n67350);
   U46050 : BUF_X1 port map( A => n65150, Z => n67260);
   U46051 : BUF_X1 port map( A => n65145, Z => n67285);
   U46052 : BUF_X1 port map( A => n65133, Z => n67351);
   U46053 : BUF_X1 port map( A => n65150, Z => n67261);
   U46054 : BUF_X1 port map( A => n65145, Z => n67286);
   U46055 : BUF_X1 port map( A => n65133, Z => n67352);
   U46056 : BUF_X1 port map( A => n65150, Z => n67262);
   U46057 : BUF_X1 port map( A => n65145, Z => n67287);
   U46058 : BUF_X1 port map( A => n65133, Z => n67353);
   U46059 : BUF_X1 port map( A => n65150, Z => n67263);
   U46060 : BUF_X1 port map( A => n65145, Z => n67288);
   U46061 : BUF_X1 port map( A => n65133, Z => n67354);
   U46062 : BUF_X1 port map( A => n65150, Z => n67264);
   U46063 : BUF_X1 port map( A => n65135, Z => n67338);
   U46064 : BUF_X1 port map( A => n65135, Z => n67339);
   U46065 : BUF_X1 port map( A => n65135, Z => n67340);
   U46066 : BUF_X1 port map( A => n65135, Z => n67341);
   U46067 : BUF_X1 port map( A => n65135, Z => n67342);
   U46068 : BUF_X1 port map( A => n63806, Z => n67524);
   U46069 : BUF_X1 port map( A => n63814, Z => n67482);
   U46070 : BUF_X1 port map( A => n63806, Z => n67525);
   U46071 : BUF_X1 port map( A => n63814, Z => n67483);
   U46072 : BUF_X1 port map( A => n63806, Z => n67526);
   U46073 : BUF_X1 port map( A => n63814, Z => n67484);
   U46074 : BUF_X1 port map( A => n63806, Z => n67527);
   U46075 : BUF_X1 port map( A => n63814, Z => n67485);
   U46076 : BUF_X1 port map( A => n63806, Z => n67528);
   U46077 : BUF_X1 port map( A => n63814, Z => n67486);
   U46078 : BUF_X1 port map( A => n63819, Z => n67458);
   U46079 : BUF_X1 port map( A => n63819, Z => n67459);
   U46080 : BUF_X1 port map( A => n63819, Z => n67460);
   U46081 : BUF_X1 port map( A => n63819, Z => n67461);
   U46082 : BUF_X1 port map( A => n63819, Z => n67462);
   U46083 : BUF_X1 port map( A => n65137, Z => n67326);
   U46084 : BUF_X1 port map( A => n65137, Z => n67327);
   U46085 : BUF_X1 port map( A => n65137, Z => n67328);
   U46086 : BUF_X1 port map( A => n65137, Z => n67329);
   U46087 : BUF_X1 port map( A => n65137, Z => n67330);
   U46088 : BUF_X1 port map( A => n63802, Z => n67548);
   U46089 : BUF_X1 port map( A => n63804, Z => n67536);
   U46090 : BUF_X1 port map( A => n63802, Z => n67549);
   U46091 : BUF_X1 port map( A => n63804, Z => n67537);
   U46092 : BUF_X1 port map( A => n63802, Z => n67550);
   U46093 : BUF_X1 port map( A => n63804, Z => n67538);
   U46094 : BUF_X1 port map( A => n63802, Z => n67551);
   U46095 : BUF_X1 port map( A => n63804, Z => n67539);
   U46096 : BUF_X1 port map( A => n63802, Z => n67552);
   U46097 : BUF_X1 port map( A => n63804, Z => n67540);
   U46098 : BUF_X1 port map( A => n65114, Z => n67422);
   U46099 : BUF_X1 port map( A => n65114, Z => n67423);
   U46100 : BUF_X1 port map( A => n65114, Z => n67424);
   U46101 : BUF_X1 port map( A => n65114, Z => n67425);
   U46102 : BUF_X1 port map( A => n65114, Z => n67426);
   U46103 : BUF_X1 port map( A => n65119, Z => n67398);
   U46104 : BUF_X1 port map( A => n65119, Z => n67399);
   U46105 : BUF_X1 port map( A => n65119, Z => n67400);
   U46106 : BUF_X1 port map( A => n65119, Z => n67401);
   U46107 : BUF_X1 port map( A => n65119, Z => n67402);
   U46108 : BUF_X1 port map( A => n63792, Z => n67572);
   U46109 : BUF_X1 port map( A => n63792, Z => n67573);
   U46110 : BUF_X1 port map( A => n63792, Z => n67574);
   U46111 : BUF_X1 port map( A => n63792, Z => n67575);
   U46112 : BUF_X1 port map( A => n63792, Z => n67576);
   U46113 : BUF_X1 port map( A => n63786, Z => n67596);
   U46114 : BUF_X1 port map( A => n63786, Z => n67597);
   U46115 : BUF_X1 port map( A => n63786, Z => n67598);
   U46116 : BUF_X1 port map( A => n63786, Z => n67599);
   U46117 : BUF_X1 port map( A => n63786, Z => n67600);
   U46118 : BUF_X1 port map( A => n65109, Z => n67446);
   U46119 : BUF_X1 port map( A => n65124, Z => n67374);
   U46120 : BUF_X1 port map( A => n65109, Z => n67447);
   U46121 : BUF_X1 port map( A => n65124, Z => n67375);
   U46122 : BUF_X1 port map( A => n65109, Z => n67448);
   U46123 : BUF_X1 port map( A => n65124, Z => n67376);
   U46124 : BUF_X1 port map( A => n65109, Z => n67449);
   U46125 : BUF_X1 port map( A => n65124, Z => n67377);
   U46126 : BUF_X1 port map( A => n65109, Z => n67450);
   U46127 : BUF_X1 port map( A => n65124, Z => n67378);
   U46128 : BUF_X1 port map( A => n63776, Z => n67642);
   U46129 : BUF_X1 port map( A => n63781, Z => n67620);
   U46130 : BUF_X1 port map( A => n63776, Z => n67643);
   U46131 : BUF_X1 port map( A => n63781, Z => n67621);
   U46132 : BUF_X1 port map( A => n63776, Z => n67644);
   U46133 : BUF_X1 port map( A => n63781, Z => n67622);
   U46134 : BUF_X1 port map( A => n63776, Z => n67645);
   U46135 : BUF_X1 port map( A => n63781, Z => n67623);
   U46136 : BUF_X1 port map( A => n63776, Z => n67646);
   U46137 : BUF_X1 port map( A => n63781, Z => n67624);
   U46138 : BUF_X1 port map( A => n65113, Z => n67428);
   U46139 : BUF_X1 port map( A => n65108, Z => n67452);
   U46140 : BUF_X1 port map( A => n63775, Z => n67648);
   U46141 : BUF_X1 port map( A => n65118, Z => n67404);
   U46142 : BUF_X1 port map( A => n65123, Z => n67380);
   U46143 : BUF_X1 port map( A => n63791, Z => n67578);
   U46144 : BUF_X1 port map( A => n63785, Z => n67602);
   U46145 : BUF_X1 port map( A => n63780, Z => n67626);
   U46146 : NAND2_X1 port map( A1 => n68057, A2 => n68258, ZN => n61959);
   U46147 : OAI21_X1 port map( B1 => n62088, B2 => n62089, A => n68052, ZN => 
                           n61957);
   U46148 : OAI21_X1 port map( B1 => n62089, B2 => n63025, A => n68053, ZN => 
                           n62959);
   U46149 : AND2_X1 port map( A1 => n66276, A2 => n66277, ZN => n65111);
   U46150 : BUF_X1 port map( A => n62493, Z => n67967);
   U46151 : BUF_X1 port map( A => n62224, Z => n68019);
   U46152 : BUF_X1 port map( A => n62357, Z => n67993);
   U46153 : BUF_X1 port map( A => n62290, Z => n68006);
   U46154 : BUF_X1 port map( A => n62157, Z => n68032);
   U46155 : BUF_X1 port map( A => n62423, Z => n67980);
   U46156 : BUF_X1 port map( A => n62626, Z => n67941);
   U46157 : BUF_X1 port map( A => n62559, Z => n67954);
   U46158 : BUF_X1 port map( A => n63161, Z => n67801);
   U46159 : BUF_X1 port map( A => n63026, Z => n67839);
   U46160 : BUF_X1 port map( A => n63362, Z => n67750);
   U46161 : BUF_X1 port map( A => n63429, Z => n67737);
   U46162 : BUF_X1 port map( A => n63764, Z => n67660);
   U46163 : BUF_X1 port map( A => n62826, Z => n67878);
   U46164 : BUF_X1 port map( A => n63095, Z => n67814);
   U46165 : BUF_X1 port map( A => n63632, Z => n67686);
   U46166 : BUF_X1 port map( A => n63698, Z => n67673);
   U46167 : BUF_X1 port map( A => n63229, Z => n67776);
   U46168 : BUF_X1 port map( A => n63296, Z => n67763);
   U46169 : BUF_X1 port map( A => n63500, Z => n67712);
   U46170 : BUF_X1 port map( A => n63566, Z => n67699);
   U46171 : BUF_X1 port map( A => n62892, Z => n67865);
   U46172 : BUF_X1 port map( A => n62764, Z => n67891);
   U46173 : BUF_X1 port map( A => n62696, Z => n67916);
   U46174 : BUF_X1 port map( A => n62090, Z => n68045);
   U46175 : BUF_X1 port map( A => n62493, Z => n67968);
   U46176 : BUF_X1 port map( A => n62224, Z => n68020);
   U46177 : BUF_X1 port map( A => n62357, Z => n67994);
   U46178 : BUF_X1 port map( A => n62290, Z => n68007);
   U46179 : BUF_X1 port map( A => n62157, Z => n68033);
   U46180 : BUF_X1 port map( A => n62423, Z => n67981);
   U46181 : BUF_X1 port map( A => n62626, Z => n67942);
   U46182 : BUF_X1 port map( A => n62559, Z => n67955);
   U46183 : BUF_X1 port map( A => n63161, Z => n67802);
   U46184 : BUF_X1 port map( A => n63026, Z => n67840);
   U46185 : BUF_X1 port map( A => n63362, Z => n67751);
   U46186 : BUF_X1 port map( A => n63429, Z => n67738);
   U46187 : BUF_X1 port map( A => n63764, Z => n67661);
   U46188 : BUF_X1 port map( A => n62826, Z => n67879);
   U46189 : BUF_X1 port map( A => n63095, Z => n67815);
   U46190 : BUF_X1 port map( A => n63632, Z => n67687);
   U46191 : BUF_X1 port map( A => n63698, Z => n67674);
   U46192 : BUF_X1 port map( A => n63229, Z => n67777);
   U46193 : BUF_X1 port map( A => n63296, Z => n67764);
   U46194 : BUF_X1 port map( A => n63500, Z => n67713);
   U46195 : BUF_X1 port map( A => n63566, Z => n67700);
   U46196 : BUF_X1 port map( A => n62892, Z => n67866);
   U46197 : BUF_X1 port map( A => n62764, Z => n67892);
   U46198 : BUF_X1 port map( A => n62696, Z => n67917);
   U46199 : BUF_X1 port map( A => n62090, Z => n68046);
   U46200 : NOR3_X1 port map( A1 => n66301, A2 => n67434, A3 => n66299, ZN => 
                           n66277);
   U46201 : NOR3_X1 port map( A1 => n66291, A2 => n66297, A3 => n66292, ZN => 
                           n66276);
   U46202 : OAI21_X1 port map( B1 => n62223, B2 => n63428, A => n68054, ZN => 
                           n63498);
   U46203 : OAI21_X1 port map( B1 => n62356, B2 => n62625, A => n68053, ZN => 
                           n62762);
   U46204 : OAI21_X1 port map( B1 => n62223, B2 => n62625, A => n68052, ZN => 
                           n62693);
   U46205 : OAI21_X1 port map( B1 => n62223, B2 => n63025, A => n68053, ZN => 
                           n63093);
   U46206 : OAI21_X1 port map( B1 => n62356, B2 => n63092, A => n68053, ZN => 
                           n63227);
   U46207 : BUF_X1 port map( A => n65112, Z => n67434);
   U46208 : BUF_X1 port map( A => n65112, Z => n67435);
   U46209 : BUF_X1 port map( A => n65112, Z => n67436);
   U46210 : BUF_X1 port map( A => n65112, Z => n67437);
   U46211 : NOR3_X1 port map( A1 => n65095, A2 => n65094, A3 => n65093, ZN => 
                           n65085);
   U46212 : OAI222_X1 port map( A1 => n62891, A2 => n67320, B1 => n63160, B2 =>
                           n67314, C1 => n62355, C2 => n67308, ZN => n66293);
   U46213 : OAI222_X1 port map( A1 => n62890, A2 => n67320, B1 => n63159, B2 =>
                           n67314, C1 => n62354, C2 => n67308, ZN => n66261);
   U46214 : OAI222_X1 port map( A1 => n62889, A2 => n67320, B1 => n63158, B2 =>
                           n67314, C1 => n62353, C2 => n67308, ZN => n66243);
   U46215 : OAI222_X1 port map( A1 => n62888, A2 => n67320, B1 => n63157, B2 =>
                           n67314, C1 => n62352, C2 => n67308, ZN => n66225);
   U46216 : OAI222_X1 port map( A1 => n62887, A2 => n67320, B1 => n63156, B2 =>
                           n67314, C1 => n62351, C2 => n67308, ZN => n66207);
   U46217 : OAI222_X1 port map( A1 => n62886, A2 => n67320, B1 => n63155, B2 =>
                           n67314, C1 => n62350, C2 => n67308, ZN => n66189);
   U46218 : OAI222_X1 port map( A1 => n62885, A2 => n67320, B1 => n63154, B2 =>
                           n67314, C1 => n62349, C2 => n67308, ZN => n66171);
   U46219 : OAI222_X1 port map( A1 => n62884, A2 => n67320, B1 => n63153, B2 =>
                           n67314, C1 => n62348, C2 => n67308, ZN => n66153);
   U46220 : OAI222_X1 port map( A1 => n62883, A2 => n67320, B1 => n63152, B2 =>
                           n67314, C1 => n62347, C2 => n67308, ZN => n66135);
   U46221 : OAI222_X1 port map( A1 => n62882, A2 => n67320, B1 => n63151, B2 =>
                           n67314, C1 => n62346, C2 => n67308, ZN => n66117);
   U46222 : OAI222_X1 port map( A1 => n62881, A2 => n67320, B1 => n63150, B2 =>
                           n67314, C1 => n62345, C2 => n67308, ZN => n66099);
   U46223 : OAI222_X1 port map( A1 => n62880, A2 => n67320, B1 => n63149, B2 =>
                           n67314, C1 => n62344, C2 => n67308, ZN => n66081);
   U46224 : OAI222_X1 port map( A1 => n62879, A2 => n67321, B1 => n63148, B2 =>
                           n67315, C1 => n62343, C2 => n67309, ZN => n66063);
   U46225 : OAI222_X1 port map( A1 => n62878, A2 => n67321, B1 => n63147, B2 =>
                           n67315, C1 => n62342, C2 => n67309, ZN => n66045);
   U46226 : OAI222_X1 port map( A1 => n62877, A2 => n67321, B1 => n63146, B2 =>
                           n67315, C1 => n62341, C2 => n67309, ZN => n66027);
   U46227 : OAI222_X1 port map( A1 => n62876, A2 => n67321, B1 => n63145, B2 =>
                           n67315, C1 => n62340, C2 => n67309, ZN => n66009);
   U46228 : OAI222_X1 port map( A1 => n62875, A2 => n67321, B1 => n63144, B2 =>
                           n67315, C1 => n62339, C2 => n67309, ZN => n65991);
   U46229 : OAI222_X1 port map( A1 => n62874, A2 => n67321, B1 => n63143, B2 =>
                           n67315, C1 => n62338, C2 => n67309, ZN => n65973);
   U46230 : OAI222_X1 port map( A1 => n62873, A2 => n67321, B1 => n63142, B2 =>
                           n67315, C1 => n62337, C2 => n67309, ZN => n65955);
   U46231 : OAI222_X1 port map( A1 => n62872, A2 => n67321, B1 => n63141, B2 =>
                           n67315, C1 => n62336, C2 => n67309, ZN => n65937);
   U46232 : OAI222_X1 port map( A1 => n62871, A2 => n67321, B1 => n63140, B2 =>
                           n67315, C1 => n62335, C2 => n67309, ZN => n65919);
   U46233 : OAI222_X1 port map( A1 => n62870, A2 => n67321, B1 => n63139, B2 =>
                           n67315, C1 => n62334, C2 => n67309, ZN => n65901);
   U46234 : OAI222_X1 port map( A1 => n62869, A2 => n67321, B1 => n63138, B2 =>
                           n67315, C1 => n62333, C2 => n67309, ZN => n65883);
   U46235 : OAI222_X1 port map( A1 => n62868, A2 => n67321, B1 => n63137, B2 =>
                           n67315, C1 => n62332, C2 => n67309, ZN => n65865);
   U46236 : OAI222_X1 port map( A1 => n62867, A2 => n67322, B1 => n63136, B2 =>
                           n67316, C1 => n62331, C2 => n67310, ZN => n65847);
   U46237 : OAI222_X1 port map( A1 => n62866, A2 => n67322, B1 => n63135, B2 =>
                           n67316, C1 => n62330, C2 => n67310, ZN => n65829);
   U46238 : OAI222_X1 port map( A1 => n62865, A2 => n67322, B1 => n63134, B2 =>
                           n67316, C1 => n62329, C2 => n67310, ZN => n65811);
   U46239 : OAI222_X1 port map( A1 => n62864, A2 => n67322, B1 => n63133, B2 =>
                           n67316, C1 => n62328, C2 => n67310, ZN => n65793);
   U46240 : OAI222_X1 port map( A1 => n62863, A2 => n67322, B1 => n63132, B2 =>
                           n67316, C1 => n62327, C2 => n67310, ZN => n65775);
   U46241 : OAI222_X1 port map( A1 => n62862, A2 => n67322, B1 => n63131, B2 =>
                           n67316, C1 => n62326, C2 => n67310, ZN => n65757);
   U46242 : OAI222_X1 port map( A1 => n62861, A2 => n67322, B1 => n63130, B2 =>
                           n67316, C1 => n62325, C2 => n67310, ZN => n65739);
   U46243 : OAI222_X1 port map( A1 => n62860, A2 => n67322, B1 => n63129, B2 =>
                           n67316, C1 => n62324, C2 => n67310, ZN => n65721);
   U46244 : OAI222_X1 port map( A1 => n62859, A2 => n67322, B1 => n63128, B2 =>
                           n67316, C1 => n62323, C2 => n67310, ZN => n65703);
   U46245 : OAI222_X1 port map( A1 => n62858, A2 => n67322, B1 => n63127, B2 =>
                           n67316, C1 => n62322, C2 => n67310, ZN => n65685);
   U46246 : OAI222_X1 port map( A1 => n62857, A2 => n67322, B1 => n63126, B2 =>
                           n67316, C1 => n62321, C2 => n67310, ZN => n65667);
   U46247 : OAI222_X1 port map( A1 => n62856, A2 => n67322, B1 => n63125, B2 =>
                           n67316, C1 => n62320, C2 => n67310, ZN => n65649);
   U46248 : OAI222_X1 port map( A1 => n62855, A2 => n67323, B1 => n63124, B2 =>
                           n67317, C1 => n62319, C2 => n67311, ZN => n65631);
   U46249 : OAI222_X1 port map( A1 => n62854, A2 => n67323, B1 => n63123, B2 =>
                           n67317, C1 => n62318, C2 => n67311, ZN => n65613);
   U46250 : OAI222_X1 port map( A1 => n62853, A2 => n67323, B1 => n63122, B2 =>
                           n67317, C1 => n62317, C2 => n67311, ZN => n65595);
   U46251 : OAI222_X1 port map( A1 => n62852, A2 => n67323, B1 => n63121, B2 =>
                           n67317, C1 => n62316, C2 => n67311, ZN => n65577);
   U46252 : OAI222_X1 port map( A1 => n62851, A2 => n67323, B1 => n63120, B2 =>
                           n67317, C1 => n62315, C2 => n67311, ZN => n65559);
   U46253 : OAI222_X1 port map( A1 => n62850, A2 => n67323, B1 => n63119, B2 =>
                           n67317, C1 => n62314, C2 => n67311, ZN => n65541);
   U46254 : OAI222_X1 port map( A1 => n62849, A2 => n67323, B1 => n63118, B2 =>
                           n67317, C1 => n62313, C2 => n67311, ZN => n65523);
   U46255 : OAI222_X1 port map( A1 => n62848, A2 => n67323, B1 => n63117, B2 =>
                           n67317, C1 => n62312, C2 => n67311, ZN => n65505);
   U46256 : OAI222_X1 port map( A1 => n62847, A2 => n67323, B1 => n63116, B2 =>
                           n67317, C1 => n62311, C2 => n67311, ZN => n65487);
   U46257 : OAI222_X1 port map( A1 => n62846, A2 => n67323, B1 => n63115, B2 =>
                           n67317, C1 => n62310, C2 => n67311, ZN => n65469);
   U46258 : OAI222_X1 port map( A1 => n62845, A2 => n67323, B1 => n63114, B2 =>
                           n67317, C1 => n62309, C2 => n67311, ZN => n65451);
   U46259 : OAI222_X1 port map( A1 => n62844, A2 => n67323, B1 => n63113, B2 =>
                           n67317, C1 => n62308, C2 => n67311, ZN => n65433);
   U46260 : OAI222_X1 port map( A1 => n62843, A2 => n67324, B1 => n63112, B2 =>
                           n67318, C1 => n62307, C2 => n67312, ZN => n65415);
   U46261 : OAI222_X1 port map( A1 => n62842, A2 => n67324, B1 => n63111, B2 =>
                           n67318, C1 => n62306, C2 => n67312, ZN => n65397);
   U46262 : OAI222_X1 port map( A1 => n62841, A2 => n67324, B1 => n63110, B2 =>
                           n67318, C1 => n62305, C2 => n67312, ZN => n65379);
   U46263 : OAI222_X1 port map( A1 => n62840, A2 => n67324, B1 => n63109, B2 =>
                           n67318, C1 => n62304, C2 => n67312, ZN => n65361);
   U46264 : OAI222_X1 port map( A1 => n62839, A2 => n67324, B1 => n63108, B2 =>
                           n67318, C1 => n62303, C2 => n67312, ZN => n65343);
   U46265 : OAI222_X1 port map( A1 => n62838, A2 => n67324, B1 => n63107, B2 =>
                           n67318, C1 => n62302, C2 => n67312, ZN => n65325);
   U46266 : OAI222_X1 port map( A1 => n62837, A2 => n67324, B1 => n63106, B2 =>
                           n67318, C1 => n62301, C2 => n67312, ZN => n65307);
   U46267 : OAI222_X1 port map( A1 => n62836, A2 => n67324, B1 => n63105, B2 =>
                           n67318, C1 => n62300, C2 => n67312, ZN => n65289);
   U46268 : OAI222_X1 port map( A1 => n62835, A2 => n67324, B1 => n63104, B2 =>
                           n67318, C1 => n62299, C2 => n67312, ZN => n65271);
   U46269 : OAI222_X1 port map( A1 => n62834, A2 => n67324, B1 => n63103, B2 =>
                           n67318, C1 => n62298, C2 => n67312, ZN => n65253);
   U46270 : OAI222_X1 port map( A1 => n62833, A2 => n67324, B1 => n63102, B2 =>
                           n67318, C1 => n62297, C2 => n67312, ZN => n65235);
   U46271 : OAI222_X1 port map( A1 => n62832, A2 => n67324, B1 => n63101, B2 =>
                           n67318, C1 => n62296, C2 => n67312, ZN => n65217);
   U46272 : OAI222_X1 port map( A1 => n63226, A2 => n67518, B1 => n62155, B2 =>
                           n67512, C1 => n62558, C2 => n67506, ZN => n65089);
   U46273 : OAI222_X1 port map( A1 => n63225, A2 => n67518, B1 => n62154, B2 =>
                           n67512, C1 => n62557, C2 => n67506, ZN => n65057);
   U46274 : OAI222_X1 port map( A1 => n63224, A2 => n67518, B1 => n62153, B2 =>
                           n67512, C1 => n62556, C2 => n67506, ZN => n65037);
   U46275 : OAI222_X1 port map( A1 => n63223, A2 => n67518, B1 => n62152, B2 =>
                           n67512, C1 => n62555, C2 => n67506, ZN => n65017);
   U46276 : OAI222_X1 port map( A1 => n63222, A2 => n67518, B1 => n62151, B2 =>
                           n67512, C1 => n62554, C2 => n67506, ZN => n64997);
   U46277 : OAI222_X1 port map( A1 => n63221, A2 => n67518, B1 => n62150, B2 =>
                           n67512, C1 => n62553, C2 => n67506, ZN => n64977);
   U46278 : OAI222_X1 port map( A1 => n63220, A2 => n67518, B1 => n62149, B2 =>
                           n67512, C1 => n62552, C2 => n67506, ZN => n64957);
   U46279 : OAI222_X1 port map( A1 => n63219, A2 => n67518, B1 => n62148, B2 =>
                           n67512, C1 => n62551, C2 => n67506, ZN => n64937);
   U46280 : OAI222_X1 port map( A1 => n63218, A2 => n67518, B1 => n62147, B2 =>
                           n67512, C1 => n62550, C2 => n67506, ZN => n64917);
   U46281 : OAI222_X1 port map( A1 => n63217, A2 => n67518, B1 => n62146, B2 =>
                           n67512, C1 => n62549, C2 => n67506, ZN => n64897);
   U46282 : OAI222_X1 port map( A1 => n63216, A2 => n67518, B1 => n62145, B2 =>
                           n67512, C1 => n62548, C2 => n67506, ZN => n64877);
   U46283 : OAI222_X1 port map( A1 => n63215, A2 => n67518, B1 => n62144, B2 =>
                           n67512, C1 => n62547, C2 => n67506, ZN => n64857);
   U46284 : OAI222_X1 port map( A1 => n63214, A2 => n67519, B1 => n62143, B2 =>
                           n67513, C1 => n62546, C2 => n67507, ZN => n64837);
   U46285 : OAI222_X1 port map( A1 => n63213, A2 => n67519, B1 => n62142, B2 =>
                           n67513, C1 => n62545, C2 => n67507, ZN => n64817);
   U46286 : OAI222_X1 port map( A1 => n63212, A2 => n67519, B1 => n62141, B2 =>
                           n67513, C1 => n62544, C2 => n67507, ZN => n64797);
   U46287 : OAI222_X1 port map( A1 => n63211, A2 => n67519, B1 => n62140, B2 =>
                           n67513, C1 => n62543, C2 => n67507, ZN => n64777);
   U46288 : OAI222_X1 port map( A1 => n63210, A2 => n67519, B1 => n62139, B2 =>
                           n67513, C1 => n62542, C2 => n67507, ZN => n64757);
   U46289 : OAI222_X1 port map( A1 => n63209, A2 => n67519, B1 => n62138, B2 =>
                           n67513, C1 => n62541, C2 => n67507, ZN => n64737);
   U46290 : OAI222_X1 port map( A1 => n63208, A2 => n67519, B1 => n62137, B2 =>
                           n67513, C1 => n62540, C2 => n67507, ZN => n64717);
   U46291 : OAI222_X1 port map( A1 => n63207, A2 => n67519, B1 => n62136, B2 =>
                           n67513, C1 => n62539, C2 => n67507, ZN => n64697);
   U46292 : OAI222_X1 port map( A1 => n63206, A2 => n67519, B1 => n62135, B2 =>
                           n67513, C1 => n62538, C2 => n67507, ZN => n64677);
   U46293 : OAI222_X1 port map( A1 => n63205, A2 => n67519, B1 => n62134, B2 =>
                           n67513, C1 => n62537, C2 => n67507, ZN => n64657);
   U46294 : OAI222_X1 port map( A1 => n63204, A2 => n67519, B1 => n62133, B2 =>
                           n67513, C1 => n62536, C2 => n67507, ZN => n64637);
   U46295 : OAI222_X1 port map( A1 => n63203, A2 => n67519, B1 => n62132, B2 =>
                           n67513, C1 => n62535, C2 => n67507, ZN => n64617);
   U46296 : OAI222_X1 port map( A1 => n63202, A2 => n67520, B1 => n62131, B2 =>
                           n67514, C1 => n62534, C2 => n67508, ZN => n64597);
   U46297 : OAI222_X1 port map( A1 => n63201, A2 => n67520, B1 => n62130, B2 =>
                           n67514, C1 => n62533, C2 => n67508, ZN => n64577);
   U46298 : OAI222_X1 port map( A1 => n63200, A2 => n67520, B1 => n62129, B2 =>
                           n67514, C1 => n62532, C2 => n67508, ZN => n64557);
   U46299 : OAI222_X1 port map( A1 => n63199, A2 => n67520, B1 => n62128, B2 =>
                           n67514, C1 => n62531, C2 => n67508, ZN => n64537);
   U46300 : OAI222_X1 port map( A1 => n63198, A2 => n67520, B1 => n62127, B2 =>
                           n67514, C1 => n62530, C2 => n67508, ZN => n64517);
   U46301 : OAI222_X1 port map( A1 => n63197, A2 => n67520, B1 => n62126, B2 =>
                           n67514, C1 => n62529, C2 => n67508, ZN => n64497);
   U46302 : OAI222_X1 port map( A1 => n63196, A2 => n67520, B1 => n62125, B2 =>
                           n67514, C1 => n62528, C2 => n67508, ZN => n64477);
   U46303 : OAI222_X1 port map( A1 => n63195, A2 => n67520, B1 => n62124, B2 =>
                           n67514, C1 => n62527, C2 => n67508, ZN => n64457);
   U46304 : OAI222_X1 port map( A1 => n63194, A2 => n67520, B1 => n62123, B2 =>
                           n67514, C1 => n62526, C2 => n67508, ZN => n64437);
   U46305 : OAI222_X1 port map( A1 => n63193, A2 => n67520, B1 => n62122, B2 =>
                           n67514, C1 => n62525, C2 => n67508, ZN => n64417);
   U46306 : OAI222_X1 port map( A1 => n63192, A2 => n67520, B1 => n62121, B2 =>
                           n67514, C1 => n62524, C2 => n67508, ZN => n64397);
   U46307 : OAI222_X1 port map( A1 => n63191, A2 => n67520, B1 => n62120, B2 =>
                           n67514, C1 => n62523, C2 => n67508, ZN => n64377);
   U46308 : OAI222_X1 port map( A1 => n63190, A2 => n67521, B1 => n62119, B2 =>
                           n67515, C1 => n62522, C2 => n67509, ZN => n64357);
   U46309 : OAI222_X1 port map( A1 => n63189, A2 => n67521, B1 => n62118, B2 =>
                           n67515, C1 => n62521, C2 => n67509, ZN => n64337);
   U46310 : OAI222_X1 port map( A1 => n63188, A2 => n67521, B1 => n62117, B2 =>
                           n67515, C1 => n62520, C2 => n67509, ZN => n64317);
   U46311 : OAI222_X1 port map( A1 => n63187, A2 => n67521, B1 => n62116, B2 =>
                           n67515, C1 => n62519, C2 => n67509, ZN => n64297);
   U46312 : OAI222_X1 port map( A1 => n63186, A2 => n67521, B1 => n62115, B2 =>
                           n67515, C1 => n62518, C2 => n67509, ZN => n64277);
   U46313 : OAI222_X1 port map( A1 => n63185, A2 => n67521, B1 => n62114, B2 =>
                           n67515, C1 => n62517, C2 => n67509, ZN => n64257);
   U46314 : OAI222_X1 port map( A1 => n63184, A2 => n67521, B1 => n62113, B2 =>
                           n67515, C1 => n62516, C2 => n67509, ZN => n64237);
   U46315 : OAI222_X1 port map( A1 => n63183, A2 => n67521, B1 => n62112, B2 =>
                           n67515, C1 => n62515, C2 => n67509, ZN => n64217);
   U46316 : OAI222_X1 port map( A1 => n63182, A2 => n67521, B1 => n62111, B2 =>
                           n67515, C1 => n62514, C2 => n67509, ZN => n64197);
   U46317 : OAI222_X1 port map( A1 => n63181, A2 => n67521, B1 => n62110, B2 =>
                           n67515, C1 => n62513, C2 => n67509, ZN => n64177);
   U46318 : OAI222_X1 port map( A1 => n63180, A2 => n67521, B1 => n62109, B2 =>
                           n67515, C1 => n62512, C2 => n67509, ZN => n64157);
   U46319 : OAI222_X1 port map( A1 => n63179, A2 => n67521, B1 => n62108, B2 =>
                           n67515, C1 => n62511, C2 => n67509, ZN => n64137);
   U46320 : OAI222_X1 port map( A1 => n63178, A2 => n67522, B1 => n62107, B2 =>
                           n67516, C1 => n62510, C2 => n67510, ZN => n64117);
   U46321 : OAI222_X1 port map( A1 => n63177, A2 => n67522, B1 => n62106, B2 =>
                           n67516, C1 => n62509, C2 => n67510, ZN => n64097);
   U46322 : OAI222_X1 port map( A1 => n63176, A2 => n67522, B1 => n62105, B2 =>
                           n67516, C1 => n62508, C2 => n67510, ZN => n64077);
   U46323 : OAI222_X1 port map( A1 => n63175, A2 => n67522, B1 => n62104, B2 =>
                           n67516, C1 => n62507, C2 => n67510, ZN => n64057);
   U46324 : OAI222_X1 port map( A1 => n63174, A2 => n67522, B1 => n62103, B2 =>
                           n67516, C1 => n62506, C2 => n67510, ZN => n64037);
   U46325 : OAI222_X1 port map( A1 => n63173, A2 => n67522, B1 => n62102, B2 =>
                           n67516, C1 => n62505, C2 => n67510, ZN => n64017);
   U46326 : OAI222_X1 port map( A1 => n63172, A2 => n67522, B1 => n62101, B2 =>
                           n67516, C1 => n62504, C2 => n67510, ZN => n63997);
   U46327 : OAI222_X1 port map( A1 => n63171, A2 => n67522, B1 => n62100, B2 =>
                           n67516, C1 => n62503, C2 => n67510, ZN => n63977);
   U46328 : OAI222_X1 port map( A1 => n63170, A2 => n67522, B1 => n62099, B2 =>
                           n67516, C1 => n62502, C2 => n67510, ZN => n63957);
   U46329 : OAI222_X1 port map( A1 => n63169, A2 => n67522, B1 => n62098, B2 =>
                           n67516, C1 => n62501, C2 => n67510, ZN => n63937);
   U46330 : OAI222_X1 port map( A1 => n63168, A2 => n67522, B1 => n62097, B2 =>
                           n67516, C1 => n62500, C2 => n67510, ZN => n63917);
   U46331 : OAI222_X1 port map( A1 => n63167, A2 => n67522, B1 => n62096, B2 =>
                           n67516, C1 => n62499, C2 => n67510, ZN => n63897);
   U46332 : OAI222_X1 port map( A1 => n62829, A2 => n67325, B1 => n63098, B2 =>
                           n67319, C1 => n62293, C2 => n67313, ZN => n65163);
   U46333 : OAI222_X1 port map( A1 => n62827, A2 => n67325, B1 => n63096, B2 =>
                           n67319, C1 => n62291, C2 => n67313, ZN => n65128);
   U46334 : OAI222_X1 port map( A1 => n62831, A2 => n67325, B1 => n63100, B2 =>
                           n67319, C1 => n62295, C2 => n67313, ZN => n65199);
   U46335 : OAI222_X1 port map( A1 => n62830, A2 => n67325, B1 => n63099, B2 =>
                           n67319, C1 => n62294, C2 => n67313, ZN => n65181);
   U46336 : NAND2_X1 port map( A1 => n65086, A2 => n65081, ZN => n63804);
   U46337 : NAND2_X1 port map( A1 => n66278, A2 => n66279, ZN => n65109);
   U46338 : NAND2_X1 port map( A1 => n66278, A2 => n66290, ZN => n65124);
   U46339 : NAND2_X1 port map( A1 => n66281, A2 => n66290, ZN => n65137);
   U46340 : NAND2_X1 port map( A1 => n66277, A2 => n66290, ZN => n65136);
   U46341 : NAND2_X1 port map( A1 => n63496, A2 => n63497, ZN => n62089);
   U46342 : BUF_X1 port map( A => n62087, Z => n68053);
   U46343 : BUF_X1 port map( A => n62087, Z => n68052);
   U46344 : BUF_X1 port map( A => n62087, Z => n68054);
   U46345 : BUF_X1 port map( A => n62087, Z => n68056);
   U46346 : BUF_X1 port map( A => n62087, Z => n68055);
   U46347 : NAND2_X1 port map( A1 => n66283, A2 => n66290, ZN => n65139);
   U46348 : NAND2_X1 port map( A1 => n66287, A2 => n66283, ZN => n65145);
   U46349 : NAND2_X1 port map( A1 => n66285, A2 => n66283, ZN => n65133);
   U46350 : NAND2_X1 port map( A1 => n66279, A2 => n66283, ZN => n65132);
   U46351 : NAND2_X1 port map( A1 => n66289, A2 => n66283, ZN => n65134);
   U46352 : NAND2_X1 port map( A1 => n66286, A2 => n66283, ZN => n65150);
   U46353 : NAND2_X1 port map( A1 => n66276, A2 => n66283, ZN => n65114);
   U46354 : NAND2_X1 port map( A1 => n65073, A2 => n65078, ZN => n63806);
   U46355 : NAND2_X1 port map( A1 => n65076, A2 => n65078, ZN => n63805);
   U46356 : NAND2_X1 port map( A1 => n65080, A2 => n65078, ZN => n63801);
   U46357 : NAND2_X1 port map( A1 => n65082, A2 => n65086, ZN => n63803);
   U46358 : NAND2_X1 port map( A1 => n65077, A2 => n65086, ZN => n63792);
   U46359 : NAND2_X1 port map( A1 => n65085, A2 => n65086, ZN => n63814);
   U46360 : NAND2_X1 port map( A1 => n66276, A2 => n66278, ZN => n65119);
   U46361 : NAND2_X1 port map( A1 => n65078, A2 => n65081, ZN => n63808);
   U46362 : OAI22_X1 port map( A1 => n62699, A2 => n67349, B1 => n62895, B2 => 
                           n67343, ZN => n65165);
   U46363 : OAI22_X1 port map( A1 => n62697, A2 => n67349, B1 => n62893, B2 => 
                           n67343, ZN => n65130);
   U46364 : OAI22_X1 port map( A1 => n62701, A2 => n67349, B1 => n62897, B2 => 
                           n67343, ZN => n65201);
   U46365 : OAI22_X1 port map( A1 => n62700, A2 => n67349, B1 => n62896, B2 => 
                           n67343, ZN => n65183);
   U46366 : OAI22_X1 port map( A1 => n63432, A2 => n67271, B1 => n62227, B2 => 
                           n67265, ZN => n65168);
   U46367 : OAI22_X1 port map( A1 => n63430, A2 => n67271, B1 => n62225, B2 => 
                           n67265, ZN => n65148);
   U46368 : OAI22_X1 port map( A1 => n63434, A2 => n67271, B1 => n62229, B2 => 
                           n67265, ZN => n65204);
   U46369 : OAI22_X1 port map( A1 => n63433, A2 => n67271, B1 => n62228, B2 => 
                           n67265, ZN => n65186);
   U46370 : OAI22_X1 port map( A1 => n63301, A2 => n67493, B1 => n63637, B2 => 
                           n67487, ZN => n63881);
   U46371 : OAI22_X1 port map( A1 => n62701, A2 => n67469, B1 => n62162, B2 => 
                           n67463, ZN => n63882);
   U46372 : OAI22_X1 port map( A1 => n63300, A2 => n67493, B1 => n63636, B2 => 
                           n67487, ZN => n63860);
   U46373 : OAI22_X1 port map( A1 => n62700, A2 => n67469, B1 => n62161, B2 => 
                           n67463, ZN => n63861);
   U46374 : OAI22_X1 port map( A1 => n63299, A2 => n67493, B1 => n63635, B2 => 
                           n67487, ZN => n63839);
   U46375 : OAI22_X1 port map( A1 => n62699, A2 => n67469, B1 => n62160, B2 => 
                           n67463, ZN => n63840);
   U46376 : OAI22_X1 port map( A1 => n63297, A2 => n67493, B1 => n63633, B2 => 
                           n67487, ZN => n63812);
   U46377 : OAI22_X1 port map( A1 => n62697, A2 => n67469, B1 => n62158, B2 => 
                           n67463, ZN => n63817);
   U46378 : OAI22_X1 port map( A1 => n63299, A2 => n67337, B1 => n63029, B2 => 
                           n67331, ZN => n65164);
   U46379 : OAI22_X1 port map( A1 => n63297, A2 => n67337, B1 => n63027, B2 => 
                           n67331, ZN => n65129);
   U46380 : OAI22_X1 port map( A1 => n63301, A2 => n67337, B1 => n63031, B2 => 
                           n67331, ZN => n65200);
   U46381 : OAI22_X1 port map( A1 => n63300, A2 => n67337, B1 => n63030, B2 => 
                           n67331, ZN => n65182);
   U46382 : OAI22_X1 port map( A1 => n62964, A2 => n67535, B1 => n62564, B2 => 
                           n67529, ZN => n63878);
   U46383 : OAI22_X1 port map( A1 => n62963, A2 => n67535, B1 => n62563, B2 => 
                           n67529, ZN => n63857);
   U46384 : OAI22_X1 port map( A1 => n62962, A2 => n67535, B1 => n62562, B2 => 
                           n67529, ZN => n63836);
   U46385 : OAI22_X1 port map( A1 => n62960, A2 => n67535, B1 => n62560, B2 => 
                           n67529, ZN => n63798);
   U46386 : NAND2_X1 port map( A1 => n66286, A2 => n66281, ZN => n65144);
   U46387 : NAND2_X1 port map( A1 => n66276, A2 => n66281, ZN => n65149);
   U46388 : NAND2_X1 port map( A1 => n66278, A2 => n66287, ZN => n65140);
   U46389 : NAND2_X1 port map( A1 => n66289, A2 => n66277, ZN => n65135);
   U46390 : OAI22_X1 port map( A1 => n62761, A2 => n67344, B1 => n62957, B2 => 
                           n67338, ZN => n66295);
   U46391 : OAI22_X1 port map( A1 => n62760, A2 => n67344, B1 => n62956, B2 => 
                           n67338, ZN => n66263);
   U46392 : OAI22_X1 port map( A1 => n62759, A2 => n67344, B1 => n62955, B2 => 
                           n67338, ZN => n66245);
   U46393 : OAI22_X1 port map( A1 => n62758, A2 => n67344, B1 => n62954, B2 => 
                           n67338, ZN => n66227);
   U46394 : OAI22_X1 port map( A1 => n62757, A2 => n67344, B1 => n62953, B2 => 
                           n67338, ZN => n66209);
   U46395 : OAI22_X1 port map( A1 => n62756, A2 => n67344, B1 => n62952, B2 => 
                           n67338, ZN => n66191);
   U46396 : OAI22_X1 port map( A1 => n62755, A2 => n67344, B1 => n62951, B2 => 
                           n67338, ZN => n66173);
   U46397 : OAI22_X1 port map( A1 => n62754, A2 => n67344, B1 => n62950, B2 => 
                           n67338, ZN => n66155);
   U46398 : OAI22_X1 port map( A1 => n62753, A2 => n67344, B1 => n62949, B2 => 
                           n67338, ZN => n66137);
   U46399 : OAI22_X1 port map( A1 => n62752, A2 => n67344, B1 => n62948, B2 => 
                           n67338, ZN => n66119);
   U46400 : OAI22_X1 port map( A1 => n62751, A2 => n67344, B1 => n62947, B2 => 
                           n67338, ZN => n66101);
   U46401 : OAI22_X1 port map( A1 => n62750, A2 => n67344, B1 => n62946, B2 => 
                           n67338, ZN => n66083);
   U46402 : OAI22_X1 port map( A1 => n62749, A2 => n67345, B1 => n62945, B2 => 
                           n67339, ZN => n66065);
   U46403 : OAI22_X1 port map( A1 => n62748, A2 => n67345, B1 => n62944, B2 => 
                           n67339, ZN => n66047);
   U46404 : OAI22_X1 port map( A1 => n62747, A2 => n67345, B1 => n62943, B2 => 
                           n67339, ZN => n66029);
   U46405 : OAI22_X1 port map( A1 => n62746, A2 => n67345, B1 => n62942, B2 => 
                           n67339, ZN => n66011);
   U46406 : OAI22_X1 port map( A1 => n62745, A2 => n67345, B1 => n62941, B2 => 
                           n67339, ZN => n65993);
   U46407 : OAI22_X1 port map( A1 => n62744, A2 => n67345, B1 => n62940, B2 => 
                           n67339, ZN => n65975);
   U46408 : OAI22_X1 port map( A1 => n62743, A2 => n67345, B1 => n62939, B2 => 
                           n67339, ZN => n65957);
   U46409 : OAI22_X1 port map( A1 => n62742, A2 => n67345, B1 => n62938, B2 => 
                           n67339, ZN => n65939);
   U46410 : OAI22_X1 port map( A1 => n62741, A2 => n67345, B1 => n62937, B2 => 
                           n67339, ZN => n65921);
   U46411 : OAI22_X1 port map( A1 => n62740, A2 => n67345, B1 => n62936, B2 => 
                           n67339, ZN => n65903);
   U46412 : OAI22_X1 port map( A1 => n62739, A2 => n67345, B1 => n62935, B2 => 
                           n67339, ZN => n65885);
   U46413 : OAI22_X1 port map( A1 => n62738, A2 => n67345, B1 => n62934, B2 => 
                           n67339, ZN => n65867);
   U46414 : OAI22_X1 port map( A1 => n62737, A2 => n67346, B1 => n62933, B2 => 
                           n67340, ZN => n65849);
   U46415 : OAI22_X1 port map( A1 => n62736, A2 => n67346, B1 => n62932, B2 => 
                           n67340, ZN => n65831);
   U46416 : OAI22_X1 port map( A1 => n62735, A2 => n67346, B1 => n62931, B2 => 
                           n67340, ZN => n65813);
   U46417 : OAI22_X1 port map( A1 => n62734, A2 => n67346, B1 => n62930, B2 => 
                           n67340, ZN => n65795);
   U46418 : OAI22_X1 port map( A1 => n62733, A2 => n67346, B1 => n62929, B2 => 
                           n67340, ZN => n65777);
   U46419 : OAI22_X1 port map( A1 => n62732, A2 => n67346, B1 => n62928, B2 => 
                           n67340, ZN => n65759);
   U46420 : OAI22_X1 port map( A1 => n62731, A2 => n67346, B1 => n62927, B2 => 
                           n67340, ZN => n65741);
   U46421 : OAI22_X1 port map( A1 => n62730, A2 => n67346, B1 => n62926, B2 => 
                           n67340, ZN => n65723);
   U46422 : OAI22_X1 port map( A1 => n62729, A2 => n67346, B1 => n62925, B2 => 
                           n67340, ZN => n65705);
   U46423 : OAI22_X1 port map( A1 => n62728, A2 => n67346, B1 => n62924, B2 => 
                           n67340, ZN => n65687);
   U46424 : OAI22_X1 port map( A1 => n62727, A2 => n67346, B1 => n62923, B2 => 
                           n67340, ZN => n65669);
   U46425 : OAI22_X1 port map( A1 => n62726, A2 => n67346, B1 => n62922, B2 => 
                           n67340, ZN => n65651);
   U46426 : OAI22_X1 port map( A1 => n62725, A2 => n67347, B1 => n62921, B2 => 
                           n67341, ZN => n65633);
   U46427 : OAI22_X1 port map( A1 => n62724, A2 => n67347, B1 => n62920, B2 => 
                           n67341, ZN => n65615);
   U46428 : OAI22_X1 port map( A1 => n62723, A2 => n67347, B1 => n62919, B2 => 
                           n67341, ZN => n65597);
   U46429 : OAI22_X1 port map( A1 => n62722, A2 => n67347, B1 => n62918, B2 => 
                           n67341, ZN => n65579);
   U46430 : OAI22_X1 port map( A1 => n62721, A2 => n67347, B1 => n62917, B2 => 
                           n67341, ZN => n65561);
   U46431 : OAI22_X1 port map( A1 => n62720, A2 => n67347, B1 => n62916, B2 => 
                           n67341, ZN => n65543);
   U46432 : OAI22_X1 port map( A1 => n62719, A2 => n67347, B1 => n62915, B2 => 
                           n67341, ZN => n65525);
   U46433 : OAI22_X1 port map( A1 => n62718, A2 => n67347, B1 => n62914, B2 => 
                           n67341, ZN => n65507);
   U46434 : OAI22_X1 port map( A1 => n62717, A2 => n67347, B1 => n62913, B2 => 
                           n67341, ZN => n65489);
   U46435 : OAI22_X1 port map( A1 => n62716, A2 => n67347, B1 => n62912, B2 => 
                           n67341, ZN => n65471);
   U46436 : OAI22_X1 port map( A1 => n62715, A2 => n67347, B1 => n62911, B2 => 
                           n67341, ZN => n65453);
   U46437 : OAI22_X1 port map( A1 => n62714, A2 => n67347, B1 => n62910, B2 => 
                           n67341, ZN => n65435);
   U46438 : OAI22_X1 port map( A1 => n62713, A2 => n67348, B1 => n62909, B2 => 
                           n67342, ZN => n65417);
   U46439 : OAI22_X1 port map( A1 => n62712, A2 => n67348, B1 => n62908, B2 => 
                           n67342, ZN => n65399);
   U46440 : OAI22_X1 port map( A1 => n62711, A2 => n67348, B1 => n62907, B2 => 
                           n67342, ZN => n65381);
   U46441 : OAI22_X1 port map( A1 => n62710, A2 => n67348, B1 => n62906, B2 => 
                           n67342, ZN => n65363);
   U46442 : OAI22_X1 port map( A1 => n62709, A2 => n67348, B1 => n62905, B2 => 
                           n67342, ZN => n65345);
   U46443 : OAI22_X1 port map( A1 => n62708, A2 => n67348, B1 => n62904, B2 => 
                           n67342, ZN => n65327);
   U46444 : OAI22_X1 port map( A1 => n62707, A2 => n67348, B1 => n62903, B2 => 
                           n67342, ZN => n65309);
   U46445 : OAI22_X1 port map( A1 => n62706, A2 => n67348, B1 => n62902, B2 => 
                           n67342, ZN => n65291);
   U46446 : OAI22_X1 port map( A1 => n62705, A2 => n67348, B1 => n62901, B2 => 
                           n67342, ZN => n65273);
   U46447 : OAI22_X1 port map( A1 => n62704, A2 => n67348, B1 => n62900, B2 => 
                           n67342, ZN => n65255);
   U46448 : OAI22_X1 port map( A1 => n62703, A2 => n67348, B1 => n62899, B2 => 
                           n67342, ZN => n65237);
   U46449 : OAI22_X1 port map( A1 => n62702, A2 => n67348, B1 => n62898, B2 => 
                           n67342, ZN => n65219);
   U46450 : OAI22_X1 port map( A1 => n62155, A2 => n67290, B1 => n62222, B2 => 
                           n67284, ZN => n66298);
   U46451 : OAI22_X1 port map( A1 => n63494, A2 => n67266, B1 => n62289, B2 => 
                           n67260, ZN => n66300);
   U46452 : OAI22_X1 port map( A1 => n62154, A2 => n67290, B1 => n62221, B2 => 
                           n67284, ZN => n66265);
   U46453 : OAI22_X1 port map( A1 => n63493, A2 => n67266, B1 => n62288, B2 => 
                           n67260, ZN => n66266);
   U46454 : OAI22_X1 port map( A1 => n62153, A2 => n67290, B1 => n62220, B2 => 
                           n67284, ZN => n66247);
   U46455 : OAI22_X1 port map( A1 => n63492, A2 => n67266, B1 => n62287, B2 => 
                           n67260, ZN => n66248);
   U46456 : OAI22_X1 port map( A1 => n62152, A2 => n67290, B1 => n62219, B2 => 
                           n67284, ZN => n66229);
   U46457 : OAI22_X1 port map( A1 => n63491, A2 => n67266, B1 => n62286, B2 => 
                           n67260, ZN => n66230);
   U46458 : OAI22_X1 port map( A1 => n62151, A2 => n67290, B1 => n62218, B2 => 
                           n67284, ZN => n66211);
   U46459 : OAI22_X1 port map( A1 => n63490, A2 => n67266, B1 => n62285, B2 => 
                           n67260, ZN => n66212);
   U46460 : OAI22_X1 port map( A1 => n62150, A2 => n67290, B1 => n62217, B2 => 
                           n67284, ZN => n66193);
   U46461 : OAI22_X1 port map( A1 => n63489, A2 => n67266, B1 => n62284, B2 => 
                           n67260, ZN => n66194);
   U46462 : OAI22_X1 port map( A1 => n62149, A2 => n67290, B1 => n62216, B2 => 
                           n67284, ZN => n66175);
   U46463 : OAI22_X1 port map( A1 => n63488, A2 => n67266, B1 => n62283, B2 => 
                           n67260, ZN => n66176);
   U46464 : OAI22_X1 port map( A1 => n62148, A2 => n67290, B1 => n62215, B2 => 
                           n67284, ZN => n66157);
   U46465 : OAI22_X1 port map( A1 => n63487, A2 => n67266, B1 => n62282, B2 => 
                           n67260, ZN => n66158);
   U46466 : OAI22_X1 port map( A1 => n62147, A2 => n67290, B1 => n62214, B2 => 
                           n67284, ZN => n66139);
   U46467 : OAI22_X1 port map( A1 => n63486, A2 => n67266, B1 => n62281, B2 => 
                           n67260, ZN => n66140);
   U46468 : OAI22_X1 port map( A1 => n62146, A2 => n67290, B1 => n62213, B2 => 
                           n67284, ZN => n66121);
   U46469 : OAI22_X1 port map( A1 => n63485, A2 => n67266, B1 => n62280, B2 => 
                           n67260, ZN => n66122);
   U46470 : OAI22_X1 port map( A1 => n62145, A2 => n67290, B1 => n62212, B2 => 
                           n67284, ZN => n66103);
   U46471 : OAI22_X1 port map( A1 => n63484, A2 => n67266, B1 => n62279, B2 => 
                           n67260, ZN => n66104);
   U46472 : OAI22_X1 port map( A1 => n62144, A2 => n67290, B1 => n62211, B2 => 
                           n67284, ZN => n66085);
   U46473 : OAI22_X1 port map( A1 => n63483, A2 => n67266, B1 => n62278, B2 => 
                           n67260, ZN => n66086);
   U46474 : OAI22_X1 port map( A1 => n62143, A2 => n67291, B1 => n62210, B2 => 
                           n67285, ZN => n66067);
   U46475 : OAI22_X1 port map( A1 => n63482, A2 => n67267, B1 => n62277, B2 => 
                           n67261, ZN => n66068);
   U46476 : OAI22_X1 port map( A1 => n62142, A2 => n67291, B1 => n62209, B2 => 
                           n67285, ZN => n66049);
   U46477 : OAI22_X1 port map( A1 => n63481, A2 => n67267, B1 => n62276, B2 => 
                           n67261, ZN => n66050);
   U46478 : OAI22_X1 port map( A1 => n62141, A2 => n67291, B1 => n62208, B2 => 
                           n67285, ZN => n66031);
   U46479 : OAI22_X1 port map( A1 => n63480, A2 => n67267, B1 => n62275, B2 => 
                           n67261, ZN => n66032);
   U46480 : OAI22_X1 port map( A1 => n62140, A2 => n67291, B1 => n62207, B2 => 
                           n67285, ZN => n66013);
   U46481 : OAI22_X1 port map( A1 => n63479, A2 => n67267, B1 => n62274, B2 => 
                           n67261, ZN => n66014);
   U46482 : OAI22_X1 port map( A1 => n62139, A2 => n67291, B1 => n62206, B2 => 
                           n67285, ZN => n65995);
   U46483 : OAI22_X1 port map( A1 => n63478, A2 => n67267, B1 => n62273, B2 => 
                           n67261, ZN => n65996);
   U46484 : OAI22_X1 port map( A1 => n62138, A2 => n67291, B1 => n62205, B2 => 
                           n67285, ZN => n65977);
   U46485 : OAI22_X1 port map( A1 => n63477, A2 => n67267, B1 => n62272, B2 => 
                           n67261, ZN => n65978);
   U46486 : OAI22_X1 port map( A1 => n62137, A2 => n67291, B1 => n62204, B2 => 
                           n67285, ZN => n65959);
   U46487 : OAI22_X1 port map( A1 => n63476, A2 => n67267, B1 => n62271, B2 => 
                           n67261, ZN => n65960);
   U46488 : OAI22_X1 port map( A1 => n62136, A2 => n67291, B1 => n62203, B2 => 
                           n67285, ZN => n65941);
   U46489 : OAI22_X1 port map( A1 => n63475, A2 => n67267, B1 => n62270, B2 => 
                           n67261, ZN => n65942);
   U46490 : OAI22_X1 port map( A1 => n62135, A2 => n67291, B1 => n62202, B2 => 
                           n67285, ZN => n65923);
   U46491 : OAI22_X1 port map( A1 => n63474, A2 => n67267, B1 => n62269, B2 => 
                           n67261, ZN => n65924);
   U46492 : OAI22_X1 port map( A1 => n62134, A2 => n67291, B1 => n62201, B2 => 
                           n67285, ZN => n65905);
   U46493 : OAI22_X1 port map( A1 => n63473, A2 => n67267, B1 => n62268, B2 => 
                           n67261, ZN => n65906);
   U46494 : OAI22_X1 port map( A1 => n62133, A2 => n67291, B1 => n62200, B2 => 
                           n67285, ZN => n65887);
   U46495 : OAI22_X1 port map( A1 => n63472, A2 => n67267, B1 => n62267, B2 => 
                           n67261, ZN => n65888);
   U46496 : OAI22_X1 port map( A1 => n62132, A2 => n67291, B1 => n62199, B2 => 
                           n67285, ZN => n65869);
   U46497 : OAI22_X1 port map( A1 => n63471, A2 => n67267, B1 => n62266, B2 => 
                           n67261, ZN => n65870);
   U46498 : OAI22_X1 port map( A1 => n62131, A2 => n67292, B1 => n62198, B2 => 
                           n67286, ZN => n65851);
   U46499 : OAI22_X1 port map( A1 => n63470, A2 => n67268, B1 => n62265, B2 => 
                           n67262, ZN => n65852);
   U46500 : OAI22_X1 port map( A1 => n62130, A2 => n67292, B1 => n62197, B2 => 
                           n67286, ZN => n65833);
   U46501 : OAI22_X1 port map( A1 => n63469, A2 => n67268, B1 => n62264, B2 => 
                           n67262, ZN => n65834);
   U46502 : OAI22_X1 port map( A1 => n62129, A2 => n67292, B1 => n62196, B2 => 
                           n67286, ZN => n65815);
   U46503 : OAI22_X1 port map( A1 => n63468, A2 => n67268, B1 => n62263, B2 => 
                           n67262, ZN => n65816);
   U46504 : OAI22_X1 port map( A1 => n62128, A2 => n67292, B1 => n62195, B2 => 
                           n67286, ZN => n65797);
   U46505 : OAI22_X1 port map( A1 => n63467, A2 => n67268, B1 => n62262, B2 => 
                           n67262, ZN => n65798);
   U46506 : OAI22_X1 port map( A1 => n62127, A2 => n67292, B1 => n62194, B2 => 
                           n67286, ZN => n65779);
   U46507 : OAI22_X1 port map( A1 => n63466, A2 => n67268, B1 => n62261, B2 => 
                           n67262, ZN => n65780);
   U46508 : OAI22_X1 port map( A1 => n62126, A2 => n67292, B1 => n62193, B2 => 
                           n67286, ZN => n65761);
   U46509 : OAI22_X1 port map( A1 => n63465, A2 => n67268, B1 => n62260, B2 => 
                           n67262, ZN => n65762);
   U46510 : OAI22_X1 port map( A1 => n62125, A2 => n67292, B1 => n62192, B2 => 
                           n67286, ZN => n65743);
   U46511 : OAI22_X1 port map( A1 => n63464, A2 => n67268, B1 => n62259, B2 => 
                           n67262, ZN => n65744);
   U46512 : OAI22_X1 port map( A1 => n62124, A2 => n67292, B1 => n62191, B2 => 
                           n67286, ZN => n65725);
   U46513 : OAI22_X1 port map( A1 => n63463, A2 => n67268, B1 => n62258, B2 => 
                           n67262, ZN => n65726);
   U46514 : OAI22_X1 port map( A1 => n62123, A2 => n67292, B1 => n62190, B2 => 
                           n67286, ZN => n65707);
   U46515 : OAI22_X1 port map( A1 => n63462, A2 => n67268, B1 => n62257, B2 => 
                           n67262, ZN => n65708);
   U46516 : OAI22_X1 port map( A1 => n62122, A2 => n67292, B1 => n62189, B2 => 
                           n67286, ZN => n65689);
   U46517 : OAI22_X1 port map( A1 => n63461, A2 => n67268, B1 => n62256, B2 => 
                           n67262, ZN => n65690);
   U46518 : OAI22_X1 port map( A1 => n62121, A2 => n67292, B1 => n62188, B2 => 
                           n67286, ZN => n65671);
   U46519 : OAI22_X1 port map( A1 => n63460, A2 => n67268, B1 => n62255, B2 => 
                           n67262, ZN => n65672);
   U46520 : OAI22_X1 port map( A1 => n62120, A2 => n67292, B1 => n62187, B2 => 
                           n67286, ZN => n65653);
   U46521 : OAI22_X1 port map( A1 => n63459, A2 => n67268, B1 => n62254, B2 => 
                           n67262, ZN => n65654);
   U46522 : OAI22_X1 port map( A1 => n62119, A2 => n67293, B1 => n62186, B2 => 
                           n67287, ZN => n65635);
   U46523 : OAI22_X1 port map( A1 => n63458, A2 => n67269, B1 => n62253, B2 => 
                           n67263, ZN => n65636);
   U46524 : OAI22_X1 port map( A1 => n62118, A2 => n67293, B1 => n62185, B2 => 
                           n67287, ZN => n65617);
   U46525 : OAI22_X1 port map( A1 => n63457, A2 => n67269, B1 => n62252, B2 => 
                           n67263, ZN => n65618);
   U46526 : OAI22_X1 port map( A1 => n62117, A2 => n67293, B1 => n62184, B2 => 
                           n67287, ZN => n65599);
   U46527 : OAI22_X1 port map( A1 => n63456, A2 => n67269, B1 => n62251, B2 => 
                           n67263, ZN => n65600);
   U46528 : OAI22_X1 port map( A1 => n62116, A2 => n67293, B1 => n62183, B2 => 
                           n67287, ZN => n65581);
   U46529 : OAI22_X1 port map( A1 => n63455, A2 => n67269, B1 => n62250, B2 => 
                           n67263, ZN => n65582);
   U46530 : OAI22_X1 port map( A1 => n62115, A2 => n67293, B1 => n62182, B2 => 
                           n67287, ZN => n65563);
   U46531 : OAI22_X1 port map( A1 => n63454, A2 => n67269, B1 => n62249, B2 => 
                           n67263, ZN => n65564);
   U46532 : OAI22_X1 port map( A1 => n62114, A2 => n67293, B1 => n62181, B2 => 
                           n67287, ZN => n65545);
   U46533 : OAI22_X1 port map( A1 => n63453, A2 => n67269, B1 => n62248, B2 => 
                           n67263, ZN => n65546);
   U46534 : OAI22_X1 port map( A1 => n62113, A2 => n67293, B1 => n62180, B2 => 
                           n67287, ZN => n65527);
   U46535 : OAI22_X1 port map( A1 => n63452, A2 => n67269, B1 => n62247, B2 => 
                           n67263, ZN => n65528);
   U46536 : OAI22_X1 port map( A1 => n62112, A2 => n67293, B1 => n62179, B2 => 
                           n67287, ZN => n65509);
   U46537 : OAI22_X1 port map( A1 => n63451, A2 => n67269, B1 => n62246, B2 => 
                           n67263, ZN => n65510);
   U46538 : OAI22_X1 port map( A1 => n62111, A2 => n67293, B1 => n62178, B2 => 
                           n67287, ZN => n65491);
   U46539 : OAI22_X1 port map( A1 => n63450, A2 => n67269, B1 => n62245, B2 => 
                           n67263, ZN => n65492);
   U46540 : OAI22_X1 port map( A1 => n62110, A2 => n67293, B1 => n62177, B2 => 
                           n67287, ZN => n65473);
   U46541 : OAI22_X1 port map( A1 => n63449, A2 => n67269, B1 => n62244, B2 => 
                           n67263, ZN => n65474);
   U46542 : OAI22_X1 port map( A1 => n62109, A2 => n67293, B1 => n62176, B2 => 
                           n67287, ZN => n65455);
   U46543 : OAI22_X1 port map( A1 => n63448, A2 => n67269, B1 => n62243, B2 => 
                           n67263, ZN => n65456);
   U46544 : OAI22_X1 port map( A1 => n62108, A2 => n67293, B1 => n62175, B2 => 
                           n67287, ZN => n65437);
   U46545 : OAI22_X1 port map( A1 => n63447, A2 => n67269, B1 => n62242, B2 => 
                           n67263, ZN => n65438);
   U46546 : OAI22_X1 port map( A1 => n62107, A2 => n67294, B1 => n62174, B2 => 
                           n67288, ZN => n65419);
   U46547 : OAI22_X1 port map( A1 => n63446, A2 => n67270, B1 => n62241, B2 => 
                           n67264, ZN => n65420);
   U46548 : OAI22_X1 port map( A1 => n62106, A2 => n67294, B1 => n62173, B2 => 
                           n67288, ZN => n65401);
   U46549 : OAI22_X1 port map( A1 => n63445, A2 => n67270, B1 => n62240, B2 => 
                           n67264, ZN => n65402);
   U46550 : OAI22_X1 port map( A1 => n62105, A2 => n67294, B1 => n62172, B2 => 
                           n67288, ZN => n65383);
   U46551 : OAI22_X1 port map( A1 => n63444, A2 => n67270, B1 => n62239, B2 => 
                           n67264, ZN => n65384);
   U46552 : OAI22_X1 port map( A1 => n62104, A2 => n67294, B1 => n62171, B2 => 
                           n67288, ZN => n65365);
   U46553 : OAI22_X1 port map( A1 => n63443, A2 => n67270, B1 => n62238, B2 => 
                           n67264, ZN => n65366);
   U46554 : OAI22_X1 port map( A1 => n62103, A2 => n67294, B1 => n62170, B2 => 
                           n67288, ZN => n65347);
   U46555 : OAI22_X1 port map( A1 => n63442, A2 => n67270, B1 => n62237, B2 => 
                           n67264, ZN => n65348);
   U46556 : OAI22_X1 port map( A1 => n62102, A2 => n67294, B1 => n62169, B2 => 
                           n67288, ZN => n65329);
   U46557 : OAI22_X1 port map( A1 => n63441, A2 => n67270, B1 => n62236, B2 => 
                           n67264, ZN => n65330);
   U46558 : OAI22_X1 port map( A1 => n62101, A2 => n67294, B1 => n62168, B2 => 
                           n67288, ZN => n65311);
   U46559 : OAI22_X1 port map( A1 => n63440, A2 => n67270, B1 => n62235, B2 => 
                           n67264, ZN => n65312);
   U46560 : OAI22_X1 port map( A1 => n62100, A2 => n67294, B1 => n62167, B2 => 
                           n67288, ZN => n65293);
   U46561 : OAI22_X1 port map( A1 => n63439, A2 => n67270, B1 => n62234, B2 => 
                           n67264, ZN => n65294);
   U46562 : OAI22_X1 port map( A1 => n62099, A2 => n67294, B1 => n62166, B2 => 
                           n67288, ZN => n65275);
   U46563 : OAI22_X1 port map( A1 => n63438, A2 => n67270, B1 => n62233, B2 => 
                           n67264, ZN => n65276);
   U46564 : OAI22_X1 port map( A1 => n62098, A2 => n67294, B1 => n62165, B2 => 
                           n67288, ZN => n65257);
   U46565 : OAI22_X1 port map( A1 => n63437, A2 => n67270, B1 => n62232, B2 => 
                           n67264, ZN => n65258);
   U46566 : OAI22_X1 port map( A1 => n62097, A2 => n67294, B1 => n62164, B2 => 
                           n67288, ZN => n65239);
   U46567 : OAI22_X1 port map( A1 => n63436, A2 => n67270, B1 => n62231, B2 => 
                           n67264, ZN => n65240);
   U46568 : OAI22_X1 port map( A1 => n62096, A2 => n67294, B1 => n62163, B2 => 
                           n67288, ZN => n65221);
   U46569 : OAI22_X1 port map( A1 => n63435, A2 => n67270, B1 => n62230, B2 => 
                           n67264, ZN => n65222);
   U46570 : OAI22_X1 port map( A1 => n63361, A2 => n67488, B1 => n63697, B2 => 
                           n67482, ZN => n65096);
   U46571 : OAI22_X1 port map( A1 => n62761, A2 => n67464, B1 => n62222, B2 => 
                           n67458, ZN => n65098);
   U46572 : OAI22_X1 port map( A1 => n63360, A2 => n67488, B1 => n63696, B2 => 
                           n67482, ZN => n65061);
   U46573 : OAI22_X1 port map( A1 => n62760, A2 => n67464, B1 => n62221, B2 => 
                           n67458, ZN => n65062);
   U46574 : OAI22_X1 port map( A1 => n63359, A2 => n67488, B1 => n63695, B2 => 
                           n67482, ZN => n65041);
   U46575 : OAI22_X1 port map( A1 => n62759, A2 => n67464, B1 => n62220, B2 => 
                           n67458, ZN => n65042);
   U46576 : OAI22_X1 port map( A1 => n63358, A2 => n67488, B1 => n63694, B2 => 
                           n67482, ZN => n65021);
   U46577 : OAI22_X1 port map( A1 => n62758, A2 => n67464, B1 => n62219, B2 => 
                           n67458, ZN => n65022);
   U46578 : OAI22_X1 port map( A1 => n63357, A2 => n67488, B1 => n63693, B2 => 
                           n67482, ZN => n65001);
   U46579 : OAI22_X1 port map( A1 => n62757, A2 => n67464, B1 => n62218, B2 => 
                           n67458, ZN => n65002);
   U46580 : OAI22_X1 port map( A1 => n63356, A2 => n67488, B1 => n63692, B2 => 
                           n67482, ZN => n64981);
   U46581 : OAI22_X1 port map( A1 => n62756, A2 => n67464, B1 => n62217, B2 => 
                           n67458, ZN => n64982);
   U46582 : OAI22_X1 port map( A1 => n63355, A2 => n67488, B1 => n63691, B2 => 
                           n67482, ZN => n64961);
   U46583 : OAI22_X1 port map( A1 => n62755, A2 => n67464, B1 => n62216, B2 => 
                           n67458, ZN => n64962);
   U46584 : OAI22_X1 port map( A1 => n63354, A2 => n67488, B1 => n63690, B2 => 
                           n67482, ZN => n64941);
   U46585 : OAI22_X1 port map( A1 => n62754, A2 => n67464, B1 => n62215, B2 => 
                           n67458, ZN => n64942);
   U46586 : OAI22_X1 port map( A1 => n63353, A2 => n67488, B1 => n63689, B2 => 
                           n67482, ZN => n64921);
   U46587 : OAI22_X1 port map( A1 => n62753, A2 => n67464, B1 => n62214, B2 => 
                           n67458, ZN => n64922);
   U46588 : OAI22_X1 port map( A1 => n63352, A2 => n67488, B1 => n63688, B2 => 
                           n67482, ZN => n64901);
   U46589 : OAI22_X1 port map( A1 => n62752, A2 => n67464, B1 => n62213, B2 => 
                           n67458, ZN => n64902);
   U46590 : OAI22_X1 port map( A1 => n63351, A2 => n67488, B1 => n63687, B2 => 
                           n67482, ZN => n64881);
   U46591 : OAI22_X1 port map( A1 => n62751, A2 => n67464, B1 => n62212, B2 => 
                           n67458, ZN => n64882);
   U46592 : OAI22_X1 port map( A1 => n63350, A2 => n67488, B1 => n63686, B2 => 
                           n67482, ZN => n64861);
   U46593 : OAI22_X1 port map( A1 => n62750, A2 => n67464, B1 => n62211, B2 => 
                           n67458, ZN => n64862);
   U46594 : OAI22_X1 port map( A1 => n63349, A2 => n67489, B1 => n63685, B2 => 
                           n67483, ZN => n64841);
   U46595 : OAI22_X1 port map( A1 => n62749, A2 => n67465, B1 => n62210, B2 => 
                           n67459, ZN => n64842);
   U46596 : OAI22_X1 port map( A1 => n63348, A2 => n67489, B1 => n63684, B2 => 
                           n67483, ZN => n64821);
   U46597 : OAI22_X1 port map( A1 => n62748, A2 => n67465, B1 => n62209, B2 => 
                           n67459, ZN => n64822);
   U46598 : OAI22_X1 port map( A1 => n63347, A2 => n67489, B1 => n63683, B2 => 
                           n67483, ZN => n64801);
   U46599 : OAI22_X1 port map( A1 => n62747, A2 => n67465, B1 => n62208, B2 => 
                           n67459, ZN => n64802);
   U46600 : OAI22_X1 port map( A1 => n63346, A2 => n67489, B1 => n63682, B2 => 
                           n67483, ZN => n64781);
   U46601 : OAI22_X1 port map( A1 => n62746, A2 => n67465, B1 => n62207, B2 => 
                           n67459, ZN => n64782);
   U46602 : OAI22_X1 port map( A1 => n63345, A2 => n67489, B1 => n63681, B2 => 
                           n67483, ZN => n64761);
   U46603 : OAI22_X1 port map( A1 => n62745, A2 => n67465, B1 => n62206, B2 => 
                           n67459, ZN => n64762);
   U46604 : OAI22_X1 port map( A1 => n63344, A2 => n67489, B1 => n63680, B2 => 
                           n67483, ZN => n64741);
   U46605 : OAI22_X1 port map( A1 => n62744, A2 => n67465, B1 => n62205, B2 => 
                           n67459, ZN => n64742);
   U46606 : OAI22_X1 port map( A1 => n63343, A2 => n67489, B1 => n63679, B2 => 
                           n67483, ZN => n64721);
   U46607 : OAI22_X1 port map( A1 => n62743, A2 => n67465, B1 => n62204, B2 => 
                           n67459, ZN => n64722);
   U46608 : OAI22_X1 port map( A1 => n63342, A2 => n67489, B1 => n63678, B2 => 
                           n67483, ZN => n64701);
   U46609 : OAI22_X1 port map( A1 => n62742, A2 => n67465, B1 => n62203, B2 => 
                           n67459, ZN => n64702);
   U46610 : OAI22_X1 port map( A1 => n63341, A2 => n67489, B1 => n63677, B2 => 
                           n67483, ZN => n64681);
   U46611 : OAI22_X1 port map( A1 => n62741, A2 => n67465, B1 => n62202, B2 => 
                           n67459, ZN => n64682);
   U46612 : OAI22_X1 port map( A1 => n63340, A2 => n67489, B1 => n63676, B2 => 
                           n67483, ZN => n64661);
   U46613 : OAI22_X1 port map( A1 => n62740, A2 => n67465, B1 => n62201, B2 => 
                           n67459, ZN => n64662);
   U46614 : OAI22_X1 port map( A1 => n63339, A2 => n67489, B1 => n63675, B2 => 
                           n67483, ZN => n64641);
   U46615 : OAI22_X1 port map( A1 => n62739, A2 => n67465, B1 => n62200, B2 => 
                           n67459, ZN => n64642);
   U46616 : OAI22_X1 port map( A1 => n63338, A2 => n67489, B1 => n63674, B2 => 
                           n67483, ZN => n64621);
   U46617 : OAI22_X1 port map( A1 => n62738, A2 => n67465, B1 => n62199, B2 => 
                           n67459, ZN => n64622);
   U46618 : OAI22_X1 port map( A1 => n63337, A2 => n67490, B1 => n63673, B2 => 
                           n67484, ZN => n64601);
   U46619 : OAI22_X1 port map( A1 => n62737, A2 => n67466, B1 => n62198, B2 => 
                           n67460, ZN => n64602);
   U46620 : OAI22_X1 port map( A1 => n63336, A2 => n67490, B1 => n63672, B2 => 
                           n67484, ZN => n64581);
   U46621 : OAI22_X1 port map( A1 => n62736, A2 => n67466, B1 => n62197, B2 => 
                           n67460, ZN => n64582);
   U46622 : OAI22_X1 port map( A1 => n63335, A2 => n67490, B1 => n63671, B2 => 
                           n67484, ZN => n64561);
   U46623 : OAI22_X1 port map( A1 => n62735, A2 => n67466, B1 => n62196, B2 => 
                           n67460, ZN => n64562);
   U46624 : OAI22_X1 port map( A1 => n63334, A2 => n67490, B1 => n63670, B2 => 
                           n67484, ZN => n64541);
   U46625 : OAI22_X1 port map( A1 => n62734, A2 => n67466, B1 => n62195, B2 => 
                           n67460, ZN => n64542);
   U46626 : OAI22_X1 port map( A1 => n63333, A2 => n67490, B1 => n63669, B2 => 
                           n67484, ZN => n64521);
   U46627 : OAI22_X1 port map( A1 => n62733, A2 => n67466, B1 => n62194, B2 => 
                           n67460, ZN => n64522);
   U46628 : OAI22_X1 port map( A1 => n63332, A2 => n67490, B1 => n63668, B2 => 
                           n67484, ZN => n64501);
   U46629 : OAI22_X1 port map( A1 => n62732, A2 => n67466, B1 => n62193, B2 => 
                           n67460, ZN => n64502);
   U46630 : OAI22_X1 port map( A1 => n63331, A2 => n67490, B1 => n63667, B2 => 
                           n67484, ZN => n64481);
   U46631 : OAI22_X1 port map( A1 => n62731, A2 => n67466, B1 => n62192, B2 => 
                           n67460, ZN => n64482);
   U46632 : OAI22_X1 port map( A1 => n63330, A2 => n67490, B1 => n63666, B2 => 
                           n67484, ZN => n64461);
   U46633 : OAI22_X1 port map( A1 => n62730, A2 => n67466, B1 => n62191, B2 => 
                           n67460, ZN => n64462);
   U46634 : OAI22_X1 port map( A1 => n63329, A2 => n67490, B1 => n63665, B2 => 
                           n67484, ZN => n64441);
   U46635 : OAI22_X1 port map( A1 => n62729, A2 => n67466, B1 => n62190, B2 => 
                           n67460, ZN => n64442);
   U46636 : OAI22_X1 port map( A1 => n63328, A2 => n67490, B1 => n63664, B2 => 
                           n67484, ZN => n64421);
   U46637 : OAI22_X1 port map( A1 => n62728, A2 => n67466, B1 => n62189, B2 => 
                           n67460, ZN => n64422);
   U46638 : OAI22_X1 port map( A1 => n63327, A2 => n67490, B1 => n63663, B2 => 
                           n67484, ZN => n64401);
   U46639 : OAI22_X1 port map( A1 => n62727, A2 => n67466, B1 => n62188, B2 => 
                           n67460, ZN => n64402);
   U46640 : OAI22_X1 port map( A1 => n63326, A2 => n67490, B1 => n63662, B2 => 
                           n67484, ZN => n64381);
   U46641 : OAI22_X1 port map( A1 => n62726, A2 => n67466, B1 => n62187, B2 => 
                           n67460, ZN => n64382);
   U46642 : OAI22_X1 port map( A1 => n63325, A2 => n67491, B1 => n63661, B2 => 
                           n67485, ZN => n64361);
   U46643 : OAI22_X1 port map( A1 => n62725, A2 => n67467, B1 => n62186, B2 => 
                           n67461, ZN => n64362);
   U46644 : OAI22_X1 port map( A1 => n63324, A2 => n67491, B1 => n63660, B2 => 
                           n67485, ZN => n64341);
   U46645 : OAI22_X1 port map( A1 => n62724, A2 => n67467, B1 => n62185, B2 => 
                           n67461, ZN => n64342);
   U46646 : OAI22_X1 port map( A1 => n63323, A2 => n67491, B1 => n63659, B2 => 
                           n67485, ZN => n64321);
   U46647 : OAI22_X1 port map( A1 => n62723, A2 => n67467, B1 => n62184, B2 => 
                           n67461, ZN => n64322);
   U46648 : OAI22_X1 port map( A1 => n63322, A2 => n67491, B1 => n63658, B2 => 
                           n67485, ZN => n64301);
   U46649 : OAI22_X1 port map( A1 => n62722, A2 => n67467, B1 => n62183, B2 => 
                           n67461, ZN => n64302);
   U46650 : OAI22_X1 port map( A1 => n63321, A2 => n67491, B1 => n63657, B2 => 
                           n67485, ZN => n64281);
   U46651 : OAI22_X1 port map( A1 => n62721, A2 => n67467, B1 => n62182, B2 => 
                           n67461, ZN => n64282);
   U46652 : OAI22_X1 port map( A1 => n63320, A2 => n67491, B1 => n63656, B2 => 
                           n67485, ZN => n64261);
   U46653 : OAI22_X1 port map( A1 => n62720, A2 => n67467, B1 => n62181, B2 => 
                           n67461, ZN => n64262);
   U46654 : OAI22_X1 port map( A1 => n63319, A2 => n67491, B1 => n63655, B2 => 
                           n67485, ZN => n64241);
   U46655 : OAI22_X1 port map( A1 => n62719, A2 => n67467, B1 => n62180, B2 => 
                           n67461, ZN => n64242);
   U46656 : OAI22_X1 port map( A1 => n63318, A2 => n67491, B1 => n63654, B2 => 
                           n67485, ZN => n64221);
   U46657 : OAI22_X1 port map( A1 => n62718, A2 => n67467, B1 => n62179, B2 => 
                           n67461, ZN => n64222);
   U46658 : OAI22_X1 port map( A1 => n63317, A2 => n67491, B1 => n63653, B2 => 
                           n67485, ZN => n64201);
   U46659 : OAI22_X1 port map( A1 => n62717, A2 => n67467, B1 => n62178, B2 => 
                           n67461, ZN => n64202);
   U46660 : OAI22_X1 port map( A1 => n63316, A2 => n67491, B1 => n63652, B2 => 
                           n67485, ZN => n64181);
   U46661 : OAI22_X1 port map( A1 => n62716, A2 => n67467, B1 => n62177, B2 => 
                           n67461, ZN => n64182);
   U46662 : OAI22_X1 port map( A1 => n63315, A2 => n67491, B1 => n63651, B2 => 
                           n67485, ZN => n64161);
   U46663 : OAI22_X1 port map( A1 => n62715, A2 => n67467, B1 => n62176, B2 => 
                           n67461, ZN => n64162);
   U46664 : OAI22_X1 port map( A1 => n63314, A2 => n67491, B1 => n63650, B2 => 
                           n67485, ZN => n64141);
   U46665 : OAI22_X1 port map( A1 => n62714, A2 => n67467, B1 => n62175, B2 => 
                           n67461, ZN => n64142);
   U46666 : OAI22_X1 port map( A1 => n63313, A2 => n67492, B1 => n63649, B2 => 
                           n67486, ZN => n64121);
   U46667 : OAI22_X1 port map( A1 => n62713, A2 => n67468, B1 => n62174, B2 => 
                           n67462, ZN => n64122);
   U46668 : OAI22_X1 port map( A1 => n63312, A2 => n67492, B1 => n63648, B2 => 
                           n67486, ZN => n64101);
   U46669 : OAI22_X1 port map( A1 => n62712, A2 => n67468, B1 => n62173, B2 => 
                           n67462, ZN => n64102);
   U46670 : OAI22_X1 port map( A1 => n63311, A2 => n67492, B1 => n63647, B2 => 
                           n67486, ZN => n64081);
   U46671 : OAI22_X1 port map( A1 => n62711, A2 => n67468, B1 => n62172, B2 => 
                           n67462, ZN => n64082);
   U46672 : OAI22_X1 port map( A1 => n63310, A2 => n67492, B1 => n63646, B2 => 
                           n67486, ZN => n64061);
   U46673 : OAI22_X1 port map( A1 => n62710, A2 => n67468, B1 => n62171, B2 => 
                           n67462, ZN => n64062);
   U46674 : OAI22_X1 port map( A1 => n63309, A2 => n67492, B1 => n63645, B2 => 
                           n67486, ZN => n64041);
   U46675 : OAI22_X1 port map( A1 => n62709, A2 => n67468, B1 => n62170, B2 => 
                           n67462, ZN => n64042);
   U46676 : OAI22_X1 port map( A1 => n63308, A2 => n67492, B1 => n63644, B2 => 
                           n67486, ZN => n64021);
   U46677 : OAI22_X1 port map( A1 => n62708, A2 => n67468, B1 => n62169, B2 => 
                           n67462, ZN => n64022);
   U46678 : OAI22_X1 port map( A1 => n63307, A2 => n67492, B1 => n63643, B2 => 
                           n67486, ZN => n64001);
   U46679 : OAI22_X1 port map( A1 => n62707, A2 => n67468, B1 => n62168, B2 => 
                           n67462, ZN => n64002);
   U46680 : OAI22_X1 port map( A1 => n63306, A2 => n67492, B1 => n63642, B2 => 
                           n67486, ZN => n63981);
   U46681 : OAI22_X1 port map( A1 => n62706, A2 => n67468, B1 => n62167, B2 => 
                           n67462, ZN => n63982);
   U46682 : OAI22_X1 port map( A1 => n63305, A2 => n67492, B1 => n63641, B2 => 
                           n67486, ZN => n63961);
   U46683 : OAI22_X1 port map( A1 => n62705, A2 => n67468, B1 => n62166, B2 => 
                           n67462, ZN => n63962);
   U46684 : OAI22_X1 port map( A1 => n63304, A2 => n67492, B1 => n63640, B2 => 
                           n67486, ZN => n63941);
   U46685 : OAI22_X1 port map( A1 => n62704, A2 => n67468, B1 => n62165, B2 => 
                           n67462, ZN => n63942);
   U46686 : OAI22_X1 port map( A1 => n63303, A2 => n67492, B1 => n63639, B2 => 
                           n67486, ZN => n63921);
   U46687 : OAI22_X1 port map( A1 => n62703, A2 => n67468, B1 => n62164, B2 => 
                           n67462, ZN => n63922);
   U46688 : OAI22_X1 port map( A1 => n63302, A2 => n67492, B1 => n63638, B2 => 
                           n67486, ZN => n63901);
   U46689 : OAI22_X1 port map( A1 => n62702, A2 => n67468, B1 => n62163, B2 => 
                           n67462, ZN => n63902);
   U46690 : OAI22_X1 port map( A1 => n63361, A2 => n67332, B1 => n63091, B2 => 
                           n67326, ZN => n66294);
   U46691 : OAI22_X1 port map( A1 => n63360, A2 => n67332, B1 => n63090, B2 => 
                           n67326, ZN => n66262);
   U46692 : OAI22_X1 port map( A1 => n63359, A2 => n67332, B1 => n63089, B2 => 
                           n67326, ZN => n66244);
   U46693 : OAI22_X1 port map( A1 => n63358, A2 => n67332, B1 => n63088, B2 => 
                           n67326, ZN => n66226);
   U46694 : OAI22_X1 port map( A1 => n63357, A2 => n67332, B1 => n63087, B2 => 
                           n67326, ZN => n66208);
   U46695 : OAI22_X1 port map( A1 => n63356, A2 => n67332, B1 => n63086, B2 => 
                           n67326, ZN => n66190);
   U46696 : OAI22_X1 port map( A1 => n63355, A2 => n67332, B1 => n63085, B2 => 
                           n67326, ZN => n66172);
   U46697 : OAI22_X1 port map( A1 => n63354, A2 => n67332, B1 => n63084, B2 => 
                           n67326, ZN => n66154);
   U46698 : OAI22_X1 port map( A1 => n63353, A2 => n67332, B1 => n63083, B2 => 
                           n67326, ZN => n66136);
   U46699 : OAI22_X1 port map( A1 => n63352, A2 => n67332, B1 => n63082, B2 => 
                           n67326, ZN => n66118);
   U46700 : OAI22_X1 port map( A1 => n63351, A2 => n67332, B1 => n63081, B2 => 
                           n67326, ZN => n66100);
   U46701 : OAI22_X1 port map( A1 => n63350, A2 => n67332, B1 => n63080, B2 => 
                           n67326, ZN => n66082);
   U46702 : OAI22_X1 port map( A1 => n63349, A2 => n67333, B1 => n63079, B2 => 
                           n67327, ZN => n66064);
   U46703 : OAI22_X1 port map( A1 => n63348, A2 => n67333, B1 => n63078, B2 => 
                           n67327, ZN => n66046);
   U46704 : OAI22_X1 port map( A1 => n63347, A2 => n67333, B1 => n63077, B2 => 
                           n67327, ZN => n66028);
   U46705 : OAI22_X1 port map( A1 => n63346, A2 => n67333, B1 => n63076, B2 => 
                           n67327, ZN => n66010);
   U46706 : OAI22_X1 port map( A1 => n63345, A2 => n67333, B1 => n63075, B2 => 
                           n67327, ZN => n65992);
   U46707 : OAI22_X1 port map( A1 => n63344, A2 => n67333, B1 => n63074, B2 => 
                           n67327, ZN => n65974);
   U46708 : OAI22_X1 port map( A1 => n63343, A2 => n67333, B1 => n63073, B2 => 
                           n67327, ZN => n65956);
   U46709 : OAI22_X1 port map( A1 => n63342, A2 => n67333, B1 => n63072, B2 => 
                           n67327, ZN => n65938);
   U46710 : OAI22_X1 port map( A1 => n63341, A2 => n67333, B1 => n63071, B2 => 
                           n67327, ZN => n65920);
   U46711 : OAI22_X1 port map( A1 => n63340, A2 => n67333, B1 => n63070, B2 => 
                           n67327, ZN => n65902);
   U46712 : OAI22_X1 port map( A1 => n63339, A2 => n67333, B1 => n63069, B2 => 
                           n67327, ZN => n65884);
   U46713 : OAI22_X1 port map( A1 => n63338, A2 => n67333, B1 => n63068, B2 => 
                           n67327, ZN => n65866);
   U46714 : OAI22_X1 port map( A1 => n63337, A2 => n67334, B1 => n63067, B2 => 
                           n67328, ZN => n65848);
   U46715 : OAI22_X1 port map( A1 => n63336, A2 => n67334, B1 => n63066, B2 => 
                           n67328, ZN => n65830);
   U46716 : OAI22_X1 port map( A1 => n63335, A2 => n67334, B1 => n63065, B2 => 
                           n67328, ZN => n65812);
   U46717 : OAI22_X1 port map( A1 => n63334, A2 => n67334, B1 => n63064, B2 => 
                           n67328, ZN => n65794);
   U46718 : OAI22_X1 port map( A1 => n63333, A2 => n67334, B1 => n63063, B2 => 
                           n67328, ZN => n65776);
   U46719 : OAI22_X1 port map( A1 => n63332, A2 => n67334, B1 => n63062, B2 => 
                           n67328, ZN => n65758);
   U46720 : OAI22_X1 port map( A1 => n63331, A2 => n67334, B1 => n63061, B2 => 
                           n67328, ZN => n65740);
   U46721 : OAI22_X1 port map( A1 => n63330, A2 => n67334, B1 => n63060, B2 => 
                           n67328, ZN => n65722);
   U46722 : OAI22_X1 port map( A1 => n63329, A2 => n67334, B1 => n63059, B2 => 
                           n67328, ZN => n65704);
   U46723 : OAI22_X1 port map( A1 => n63328, A2 => n67334, B1 => n63058, B2 => 
                           n67328, ZN => n65686);
   U46724 : OAI22_X1 port map( A1 => n63327, A2 => n67334, B1 => n63057, B2 => 
                           n67328, ZN => n65668);
   U46725 : OAI22_X1 port map( A1 => n63326, A2 => n67334, B1 => n63056, B2 => 
                           n67328, ZN => n65650);
   U46726 : OAI22_X1 port map( A1 => n63325, A2 => n67335, B1 => n63055, B2 => 
                           n67329, ZN => n65632);
   U46727 : OAI22_X1 port map( A1 => n63324, A2 => n67335, B1 => n63054, B2 => 
                           n67329, ZN => n65614);
   U46728 : OAI22_X1 port map( A1 => n63323, A2 => n67335, B1 => n63053, B2 => 
                           n67329, ZN => n65596);
   U46729 : OAI22_X1 port map( A1 => n63322, A2 => n67335, B1 => n63052, B2 => 
                           n67329, ZN => n65578);
   U46730 : OAI22_X1 port map( A1 => n63321, A2 => n67335, B1 => n63051, B2 => 
                           n67329, ZN => n65560);
   U46731 : OAI22_X1 port map( A1 => n63320, A2 => n67335, B1 => n63050, B2 => 
                           n67329, ZN => n65542);
   U46732 : OAI22_X1 port map( A1 => n63319, A2 => n67335, B1 => n63049, B2 => 
                           n67329, ZN => n65524);
   U46733 : OAI22_X1 port map( A1 => n63318, A2 => n67335, B1 => n63048, B2 => 
                           n67329, ZN => n65506);
   U46734 : OAI22_X1 port map( A1 => n63317, A2 => n67335, B1 => n63047, B2 => 
                           n67329, ZN => n65488);
   U46735 : OAI22_X1 port map( A1 => n63316, A2 => n67335, B1 => n63046, B2 => 
                           n67329, ZN => n65470);
   U46736 : OAI22_X1 port map( A1 => n63315, A2 => n67335, B1 => n63045, B2 => 
                           n67329, ZN => n65452);
   U46737 : OAI22_X1 port map( A1 => n63314, A2 => n67335, B1 => n63044, B2 => 
                           n67329, ZN => n65434);
   U46738 : OAI22_X1 port map( A1 => n63313, A2 => n67336, B1 => n63043, B2 => 
                           n67330, ZN => n65416);
   U46739 : OAI22_X1 port map( A1 => n63312, A2 => n67336, B1 => n63042, B2 => 
                           n67330, ZN => n65398);
   U46740 : OAI22_X1 port map( A1 => n63311, A2 => n67336, B1 => n63041, B2 => 
                           n67330, ZN => n65380);
   U46741 : OAI22_X1 port map( A1 => n63310, A2 => n67336, B1 => n63040, B2 => 
                           n67330, ZN => n65362);
   U46742 : OAI22_X1 port map( A1 => n63309, A2 => n67336, B1 => n63039, B2 => 
                           n67330, ZN => n65344);
   U46743 : OAI22_X1 port map( A1 => n63308, A2 => n67336, B1 => n63038, B2 => 
                           n67330, ZN => n65326);
   U46744 : OAI22_X1 port map( A1 => n63307, A2 => n67336, B1 => n63037, B2 => 
                           n67330, ZN => n65308);
   U46745 : OAI22_X1 port map( A1 => n63306, A2 => n67336, B1 => n63036, B2 => 
                           n67330, ZN => n65290);
   U46746 : OAI22_X1 port map( A1 => n63305, A2 => n67336, B1 => n63035, B2 => 
                           n67330, ZN => n65272);
   U46747 : OAI22_X1 port map( A1 => n63304, A2 => n67336, B1 => n63034, B2 => 
                           n67330, ZN => n65254);
   U46748 : OAI22_X1 port map( A1 => n63303, A2 => n67336, B1 => n63033, B2 => 
                           n67330, ZN => n65236);
   U46749 : OAI22_X1 port map( A1 => n63302, A2 => n67336, B1 => n63032, B2 => 
                           n67330, ZN => n65218);
   U46750 : OAI22_X1 port map( A1 => n63024, A2 => n67530, B1 => n62624, B2 => 
                           n67524, ZN => n65090);
   U46751 : OAI22_X1 port map( A1 => n63023, A2 => n67530, B1 => n62623, B2 => 
                           n67524, ZN => n65058);
   U46752 : OAI22_X1 port map( A1 => n63022, A2 => n67530, B1 => n62622, B2 => 
                           n67524, ZN => n65038);
   U46753 : OAI22_X1 port map( A1 => n63021, A2 => n67530, B1 => n62621, B2 => 
                           n67524, ZN => n65018);
   U46754 : OAI22_X1 port map( A1 => n63020, A2 => n67530, B1 => n62620, B2 => 
                           n67524, ZN => n64998);
   U46755 : OAI22_X1 port map( A1 => n63019, A2 => n67530, B1 => n62619, B2 => 
                           n67524, ZN => n64978);
   U46756 : OAI22_X1 port map( A1 => n63018, A2 => n67530, B1 => n62618, B2 => 
                           n67524, ZN => n64958);
   U46757 : OAI22_X1 port map( A1 => n63017, A2 => n67530, B1 => n62617, B2 => 
                           n67524, ZN => n64938);
   U46758 : OAI22_X1 port map( A1 => n63016, A2 => n67530, B1 => n62616, B2 => 
                           n67524, ZN => n64918);
   U46759 : OAI22_X1 port map( A1 => n63015, A2 => n67530, B1 => n62615, B2 => 
                           n67524, ZN => n64898);
   U46760 : OAI22_X1 port map( A1 => n63014, A2 => n67530, B1 => n62614, B2 => 
                           n67524, ZN => n64878);
   U46761 : OAI22_X1 port map( A1 => n63013, A2 => n67530, B1 => n62613, B2 => 
                           n67524, ZN => n64858);
   U46762 : OAI22_X1 port map( A1 => n63012, A2 => n67531, B1 => n62612, B2 => 
                           n67525, ZN => n64838);
   U46763 : OAI22_X1 port map( A1 => n63011, A2 => n67531, B1 => n62611, B2 => 
                           n67525, ZN => n64818);
   U46764 : OAI22_X1 port map( A1 => n63010, A2 => n67531, B1 => n62610, B2 => 
                           n67525, ZN => n64798);
   U46765 : OAI22_X1 port map( A1 => n63009, A2 => n67531, B1 => n62609, B2 => 
                           n67525, ZN => n64778);
   U46766 : OAI22_X1 port map( A1 => n63008, A2 => n67531, B1 => n62608, B2 => 
                           n67525, ZN => n64758);
   U46767 : OAI22_X1 port map( A1 => n63007, A2 => n67531, B1 => n62607, B2 => 
                           n67525, ZN => n64738);
   U46768 : OAI22_X1 port map( A1 => n63006, A2 => n67531, B1 => n62606, B2 => 
                           n67525, ZN => n64718);
   U46769 : OAI22_X1 port map( A1 => n63005, A2 => n67531, B1 => n62605, B2 => 
                           n67525, ZN => n64698);
   U46770 : OAI22_X1 port map( A1 => n63004, A2 => n67531, B1 => n62604, B2 => 
                           n67525, ZN => n64678);
   U46771 : OAI22_X1 port map( A1 => n63003, A2 => n67531, B1 => n62603, B2 => 
                           n67525, ZN => n64658);
   U46772 : OAI22_X1 port map( A1 => n63002, A2 => n67531, B1 => n62602, B2 => 
                           n67525, ZN => n64638);
   U46773 : OAI22_X1 port map( A1 => n63001, A2 => n67531, B1 => n62601, B2 => 
                           n67525, ZN => n64618);
   U46774 : OAI22_X1 port map( A1 => n63000, A2 => n67532, B1 => n62600, B2 => 
                           n67526, ZN => n64598);
   U46775 : OAI22_X1 port map( A1 => n62999, A2 => n67532, B1 => n62599, B2 => 
                           n67526, ZN => n64578);
   U46776 : OAI22_X1 port map( A1 => n62998, A2 => n67532, B1 => n62598, B2 => 
                           n67526, ZN => n64558);
   U46777 : OAI22_X1 port map( A1 => n62997, A2 => n67532, B1 => n62597, B2 => 
                           n67526, ZN => n64538);
   U46778 : OAI22_X1 port map( A1 => n62996, A2 => n67532, B1 => n62596, B2 => 
                           n67526, ZN => n64518);
   U46779 : OAI22_X1 port map( A1 => n62995, A2 => n67532, B1 => n62595, B2 => 
                           n67526, ZN => n64498);
   U46780 : OAI22_X1 port map( A1 => n62994, A2 => n67532, B1 => n62594, B2 => 
                           n67526, ZN => n64478);
   U46781 : OAI22_X1 port map( A1 => n62993, A2 => n67532, B1 => n62593, B2 => 
                           n67526, ZN => n64458);
   U46782 : OAI22_X1 port map( A1 => n62992, A2 => n67532, B1 => n62592, B2 => 
                           n67526, ZN => n64438);
   U46783 : OAI22_X1 port map( A1 => n62991, A2 => n67532, B1 => n62591, B2 => 
                           n67526, ZN => n64418);
   U46784 : OAI22_X1 port map( A1 => n62990, A2 => n67532, B1 => n62590, B2 => 
                           n67526, ZN => n64398);
   U46785 : OAI22_X1 port map( A1 => n62989, A2 => n67532, B1 => n62589, B2 => 
                           n67526, ZN => n64378);
   U46786 : OAI22_X1 port map( A1 => n62988, A2 => n67533, B1 => n62588, B2 => 
                           n67527, ZN => n64358);
   U46787 : OAI22_X1 port map( A1 => n62987, A2 => n67533, B1 => n62587, B2 => 
                           n67527, ZN => n64338);
   U46788 : OAI22_X1 port map( A1 => n62986, A2 => n67533, B1 => n62586, B2 => 
                           n67527, ZN => n64318);
   U46789 : OAI22_X1 port map( A1 => n62985, A2 => n67533, B1 => n62585, B2 => 
                           n67527, ZN => n64298);
   U46790 : OAI22_X1 port map( A1 => n62984, A2 => n67533, B1 => n62584, B2 => 
                           n67527, ZN => n64278);
   U46791 : OAI22_X1 port map( A1 => n62983, A2 => n67533, B1 => n62583, B2 => 
                           n67527, ZN => n64258);
   U46792 : OAI22_X1 port map( A1 => n62982, A2 => n67533, B1 => n62582, B2 => 
                           n67527, ZN => n64238);
   U46793 : OAI22_X1 port map( A1 => n62981, A2 => n67533, B1 => n62581, B2 => 
                           n67527, ZN => n64218);
   U46794 : OAI22_X1 port map( A1 => n62980, A2 => n67533, B1 => n62580, B2 => 
                           n67527, ZN => n64198);
   U46795 : OAI22_X1 port map( A1 => n62979, A2 => n67533, B1 => n62579, B2 => 
                           n67527, ZN => n64178);
   U46796 : OAI22_X1 port map( A1 => n62978, A2 => n67533, B1 => n62578, B2 => 
                           n67527, ZN => n64158);
   U46797 : OAI22_X1 port map( A1 => n62977, A2 => n67533, B1 => n62577, B2 => 
                           n67527, ZN => n64138);
   U46798 : OAI22_X1 port map( A1 => n62976, A2 => n67534, B1 => n62576, B2 => 
                           n67528, ZN => n64118);
   U46799 : OAI22_X1 port map( A1 => n62975, A2 => n67534, B1 => n62575, B2 => 
                           n67528, ZN => n64098);
   U46800 : OAI22_X1 port map( A1 => n62974, A2 => n67534, B1 => n62574, B2 => 
                           n67528, ZN => n64078);
   U46801 : OAI22_X1 port map( A1 => n62973, A2 => n67534, B1 => n62573, B2 => 
                           n67528, ZN => n64058);
   U46802 : OAI22_X1 port map( A1 => n62972, A2 => n67534, B1 => n62572, B2 => 
                           n67528, ZN => n64038);
   U46803 : OAI22_X1 port map( A1 => n62971, A2 => n67534, B1 => n62571, B2 => 
                           n67528, ZN => n64018);
   U46804 : OAI22_X1 port map( A1 => n62970, A2 => n67534, B1 => n62570, B2 => 
                           n67528, ZN => n63998);
   U46805 : OAI22_X1 port map( A1 => n62969, A2 => n67534, B1 => n62569, B2 => 
                           n67528, ZN => n63978);
   U46806 : OAI22_X1 port map( A1 => n62968, A2 => n67534, B1 => n62568, B2 => 
                           n67528, ZN => n63958);
   U46807 : OAI22_X1 port map( A1 => n62967, A2 => n67534, B1 => n62567, B2 => 
                           n67528, ZN => n63938);
   U46808 : OAI22_X1 port map( A1 => n62966, A2 => n67534, B1 => n62566, B2 => 
                           n67528, ZN => n63918);
   U46809 : OAI22_X1 port map( A1 => n62965, A2 => n67534, B1 => n62565, B2 => 
                           n67528, ZN => n63898);
   U46810 : NAND2_X1 port map( A1 => n66277, A2 => n66279, ZN => n65138);
   U46811 : NAND2_X1 port map( A1 => n65082, A2 => n65074, ZN => n63813);
   U46812 : BUF_X1 port map( A => n61966, Z => n68239);
   U46813 : BUF_X1 port map( A => n61964, Z => n68242);
   U46814 : BUF_X1 port map( A => n61962, Z => n68245);
   U46815 : BUF_X1 port map( A => n61960, Z => n68248);
   U46816 : BUF_X1 port map( A => n62086, Z => n68059);
   U46817 : BUF_X1 port map( A => n62084, Z => n68062);
   U46818 : BUF_X1 port map( A => n62082, Z => n68065);
   U46819 : BUF_X1 port map( A => n62080, Z => n68068);
   U46820 : BUF_X1 port map( A => n62078, Z => n68071);
   U46821 : BUF_X1 port map( A => n62076, Z => n68074);
   U46822 : BUF_X1 port map( A => n62074, Z => n68077);
   U46823 : BUF_X1 port map( A => n62072, Z => n68080);
   U46824 : BUF_X1 port map( A => n62070, Z => n68083);
   U46825 : BUF_X1 port map( A => n62068, Z => n68086);
   U46826 : BUF_X1 port map( A => n62066, Z => n68089);
   U46827 : BUF_X1 port map( A => n62064, Z => n68092);
   U46828 : BUF_X1 port map( A => n62062, Z => n68095);
   U46829 : BUF_X1 port map( A => n62060, Z => n68098);
   U46830 : BUF_X1 port map( A => n62058, Z => n68101);
   U46831 : BUF_X1 port map( A => n62056, Z => n68104);
   U46832 : BUF_X1 port map( A => n62054, Z => n68107);
   U46833 : BUF_X1 port map( A => n62052, Z => n68110);
   U46834 : BUF_X1 port map( A => n62050, Z => n68113);
   U46835 : BUF_X1 port map( A => n62048, Z => n68116);
   U46836 : BUF_X1 port map( A => n62046, Z => n68119);
   U46837 : BUF_X1 port map( A => n62044, Z => n68122);
   U46838 : BUF_X1 port map( A => n62042, Z => n68125);
   U46839 : BUF_X1 port map( A => n62040, Z => n68128);
   U46840 : BUF_X1 port map( A => n62038, Z => n68131);
   U46841 : BUF_X1 port map( A => n62036, Z => n68134);
   U46842 : BUF_X1 port map( A => n62034, Z => n68137);
   U46843 : BUF_X1 port map( A => n62032, Z => n68140);
   U46844 : BUF_X1 port map( A => n62030, Z => n68143);
   U46845 : BUF_X1 port map( A => n62028, Z => n68146);
   U46846 : BUF_X1 port map( A => n62026, Z => n68149);
   U46847 : BUF_X1 port map( A => n62024, Z => n68152);
   U46848 : BUF_X1 port map( A => n62022, Z => n68155);
   U46849 : BUF_X1 port map( A => n62020, Z => n68158);
   U46850 : BUF_X1 port map( A => n62018, Z => n68161);
   U46851 : BUF_X1 port map( A => n62016, Z => n68164);
   U46852 : BUF_X1 port map( A => n62014, Z => n68167);
   U46853 : BUF_X1 port map( A => n62012, Z => n68170);
   U46854 : BUF_X1 port map( A => n62010, Z => n68173);
   U46855 : BUF_X1 port map( A => n62008, Z => n68176);
   U46856 : BUF_X1 port map( A => n62006, Z => n68179);
   U46857 : BUF_X1 port map( A => n62004, Z => n68182);
   U46858 : BUF_X1 port map( A => n62002, Z => n68185);
   U46859 : BUF_X1 port map( A => n62000, Z => n68188);
   U46860 : BUF_X1 port map( A => n61998, Z => n68191);
   U46861 : BUF_X1 port map( A => n61996, Z => n68194);
   U46862 : BUF_X1 port map( A => n61994, Z => n68197);
   U46863 : BUF_X1 port map( A => n61992, Z => n68200);
   U46864 : BUF_X1 port map( A => n61990, Z => n68203);
   U46865 : BUF_X1 port map( A => n61988, Z => n68206);
   U46866 : BUF_X1 port map( A => n61986, Z => n68209);
   U46867 : BUF_X1 port map( A => n61984, Z => n68212);
   U46868 : BUF_X1 port map( A => n61982, Z => n68215);
   U46869 : BUF_X1 port map( A => n61980, Z => n68218);
   U46870 : BUF_X1 port map( A => n61978, Z => n68221);
   U46871 : BUF_X1 port map( A => n61976, Z => n68224);
   U46872 : BUF_X1 port map( A => n61974, Z => n68227);
   U46873 : BUF_X1 port map( A => n61972, Z => n68230);
   U46874 : BUF_X1 port map( A => n61970, Z => n68233);
   U46875 : BUF_X1 port map( A => n61968, Z => n68236);
   U46876 : BUF_X1 port map( A => n65112, Z => n67438);
   U46877 : NAND2_X1 port map( A1 => n65085, A2 => n65075, ZN => n63786);
   U46878 : NAND2_X1 port map( A1 => n65080, A2 => n65075, ZN => n63818);
   U46879 : NAND2_X1 port map( A1 => n65087, A2 => n65075, ZN => n63819);
   U46880 : NAND2_X1 port map( A1 => n66280, A2 => n66283, ZN => n65113);
   U46881 : NAND2_X1 port map( A1 => n65075, A2 => n65077, ZN => n63802);
   U46882 : NAND2_X1 port map( A1 => n65075, A2 => n65076, ZN => n63776);
   U46883 : NAND2_X1 port map( A1 => n65075, A2 => n65081, ZN => n63781);
   U46884 : BUF_X1 port map( A => n61966, Z => n68238);
   U46885 : BUF_X1 port map( A => n61964, Z => n68241);
   U46886 : BUF_X1 port map( A => n61962, Z => n68244);
   U46887 : BUF_X1 port map( A => n61960, Z => n68247);
   U46888 : BUF_X1 port map( A => n62086, Z => n68058);
   U46889 : BUF_X1 port map( A => n62084, Z => n68061);
   U46890 : BUF_X1 port map( A => n62082, Z => n68064);
   U46891 : BUF_X1 port map( A => n62080, Z => n68067);
   U46892 : BUF_X1 port map( A => n62078, Z => n68070);
   U46893 : BUF_X1 port map( A => n62076, Z => n68073);
   U46894 : BUF_X1 port map( A => n62074, Z => n68076);
   U46895 : BUF_X1 port map( A => n62072, Z => n68079);
   U46896 : BUF_X1 port map( A => n62070, Z => n68082);
   U46897 : BUF_X1 port map( A => n62068, Z => n68085);
   U46898 : BUF_X1 port map( A => n62066, Z => n68088);
   U46899 : BUF_X1 port map( A => n62064, Z => n68091);
   U46900 : BUF_X1 port map( A => n62062, Z => n68094);
   U46901 : BUF_X1 port map( A => n62060, Z => n68097);
   U46902 : BUF_X1 port map( A => n62058, Z => n68100);
   U46903 : BUF_X1 port map( A => n62056, Z => n68103);
   U46904 : BUF_X1 port map( A => n62054, Z => n68106);
   U46905 : BUF_X1 port map( A => n62052, Z => n68109);
   U46906 : BUF_X1 port map( A => n62050, Z => n68112);
   U46907 : BUF_X1 port map( A => n62048, Z => n68115);
   U46908 : BUF_X1 port map( A => n62046, Z => n68118);
   U46909 : BUF_X1 port map( A => n62044, Z => n68121);
   U46910 : BUF_X1 port map( A => n62042, Z => n68124);
   U46911 : BUF_X1 port map( A => n62040, Z => n68127);
   U46912 : BUF_X1 port map( A => n62038, Z => n68130);
   U46913 : BUF_X1 port map( A => n62036, Z => n68133);
   U46914 : BUF_X1 port map( A => n62034, Z => n68136);
   U46915 : BUF_X1 port map( A => n62032, Z => n68139);
   U46916 : BUF_X1 port map( A => n62030, Z => n68142);
   U46917 : BUF_X1 port map( A => n62028, Z => n68145);
   U46918 : BUF_X1 port map( A => n62026, Z => n68148);
   U46919 : BUF_X1 port map( A => n62024, Z => n68151);
   U46920 : BUF_X1 port map( A => n62022, Z => n68154);
   U46921 : BUF_X1 port map( A => n62020, Z => n68157);
   U46922 : BUF_X1 port map( A => n62018, Z => n68160);
   U46923 : BUF_X1 port map( A => n62016, Z => n68163);
   U46924 : BUF_X1 port map( A => n62014, Z => n68166);
   U46925 : BUF_X1 port map( A => n62012, Z => n68169);
   U46926 : BUF_X1 port map( A => n62010, Z => n68172);
   U46927 : BUF_X1 port map( A => n62008, Z => n68175);
   U46928 : BUF_X1 port map( A => n62006, Z => n68178);
   U46929 : BUF_X1 port map( A => n62004, Z => n68181);
   U46930 : BUF_X1 port map( A => n62002, Z => n68184);
   U46931 : BUF_X1 port map( A => n62000, Z => n68187);
   U46932 : BUF_X1 port map( A => n61998, Z => n68190);
   U46933 : BUF_X1 port map( A => n61996, Z => n68193);
   U46934 : BUF_X1 port map( A => n61994, Z => n68196);
   U46935 : BUF_X1 port map( A => n61992, Z => n68199);
   U46936 : BUF_X1 port map( A => n61990, Z => n68202);
   U46937 : BUF_X1 port map( A => n61988, Z => n68205);
   U46938 : BUF_X1 port map( A => n61986, Z => n68208);
   U46939 : BUF_X1 port map( A => n61984, Z => n68211);
   U46940 : BUF_X1 port map( A => n61982, Z => n68214);
   U46941 : BUF_X1 port map( A => n61980, Z => n68217);
   U46942 : BUF_X1 port map( A => n61978, Z => n68220);
   U46943 : BUF_X1 port map( A => n61976, Z => n68223);
   U46944 : BUF_X1 port map( A => n61974, Z => n68226);
   U46945 : BUF_X1 port map( A => n61972, Z => n68229);
   U46946 : BUF_X1 port map( A => n61970, Z => n68232);
   U46947 : BUF_X1 port map( A => n61968, Z => n68235);
   U46948 : OAI22_X1 port map( A1 => n67934, A2 => n62694, B1 => n68247, B2 => 
                           n67928, ZN => n6846);
   U46949 : NAND2_X1 port map( A1 => n65077, A2 => n65078, ZN => n63775);
   U46950 : OAI22_X1 port map( A1 => n67947, A2 => n62631, B1 => n68238, B2 => 
                           n67940, ZN => n6907);
   U46951 : OAI22_X1 port map( A1 => n67947, A2 => n62630, B1 => n68241, B2 => 
                           n67940, ZN => n6908);
   U46952 : OAI22_X1 port map( A1 => n67947, A2 => n62629, B1 => n68244, B2 => 
                           n67940, ZN => n6909);
   U46953 : OAI22_X1 port map( A1 => n67947, A2 => n62627, B1 => n68247, B2 => 
                           n67940, ZN => n6910);
   U46954 : OAI22_X1 port map( A1 => n67960, A2 => n62564, B1 => n68238, B2 => 
                           n67953, ZN => n6971);
   U46955 : OAI22_X1 port map( A1 => n67960, A2 => n62563, B1 => n68241, B2 => 
                           n67953, ZN => n6972);
   U46956 : OAI22_X1 port map( A1 => n67960, A2 => n62562, B1 => n68244, B2 => 
                           n67953, ZN => n6973);
   U46957 : OAI22_X1 port map( A1 => n67960, A2 => n62560, B1 => n68247, B2 => 
                           n67953, ZN => n6974);
   U46958 : OAI22_X1 port map( A1 => n68051, A2 => n62095, B1 => n68238, B2 => 
                           n68044, ZN => n7419);
   U46959 : OAI22_X1 port map( A1 => n68051, A2 => n62094, B1 => n68241, B2 => 
                           n68044, ZN => n7420);
   U46960 : OAI22_X1 port map( A1 => n68051, A2 => n62093, B1 => n68244, B2 => 
                           n68044, ZN => n7421);
   U46961 : OAI22_X1 port map( A1 => n68051, A2 => n62091, B1 => n68247, B2 => 
                           n68044, ZN => n7422);
   U46962 : OAI22_X1 port map( A1 => n68012, A2 => n62295, B1 => n68238, B2 => 
                           n68005, ZN => n7227);
   U46963 : OAI22_X1 port map( A1 => n68012, A2 => n62294, B1 => n68241, B2 => 
                           n68005, ZN => n7228);
   U46964 : OAI22_X1 port map( A1 => n68012, A2 => n62293, B1 => n68244, B2 => 
                           n68005, ZN => n7229);
   U46965 : OAI22_X1 port map( A1 => n68012, A2 => n62291, B1 => n68247, B2 => 
                           n68005, ZN => n7230);
   U46966 : OAI22_X1 port map( A1 => n67973, A2 => n62498, B1 => n68238, B2 => 
                           n67966, ZN => n7035);
   U46967 : OAI22_X1 port map( A1 => n67973, A2 => n62497, B1 => n68241, B2 => 
                           n67966, ZN => n7036);
   U46968 : OAI22_X1 port map( A1 => n67973, A2 => n62496, B1 => n68244, B2 => 
                           n67966, ZN => n7037);
   U46969 : OAI22_X1 port map( A1 => n67973, A2 => n62494, B1 => n68247, B2 => 
                           n67966, ZN => n7038);
   U46970 : OAI22_X1 port map( A1 => n67807, A2 => n63166, B1 => n68239, B2 => 
                           n67800, ZN => n6203);
   U46971 : OAI22_X1 port map( A1 => n67807, A2 => n63165, B1 => n68242, B2 => 
                           n67800, ZN => n6204);
   U46972 : OAI22_X1 port map( A1 => n67807, A2 => n63164, B1 => n68245, B2 => 
                           n67800, ZN => n6205);
   U46973 : OAI22_X1 port map( A1 => n67807, A2 => n63162, B1 => n68248, B2 => 
                           n67800, ZN => n6206);
   U46974 : OAI22_X1 port map( A1 => n67858, A2 => n62964, B1 => n68239, B2 => 
                           n67851, ZN => n6459);
   U46975 : OAI22_X1 port map( A1 => n67858, A2 => n62963, B1 => n68242, B2 => 
                           n67851, ZN => n6460);
   U46976 : OAI22_X1 port map( A1 => n67858, A2 => n62962, B1 => n68245, B2 => 
                           n67851, ZN => n6461);
   U46977 : OAI22_X1 port map( A1 => n67858, A2 => n62960, B1 => n68248, B2 => 
                           n67851, ZN => n6462);
   U46978 : OAI22_X1 port map( A1 => n67845, A2 => n63031, B1 => n68239, B2 => 
                           n67838, ZN => n6395);
   U46979 : OAI22_X1 port map( A1 => n67845, A2 => n63030, B1 => n68242, B2 => 
                           n67838, ZN => n6396);
   U46980 : OAI22_X1 port map( A1 => n67845, A2 => n63029, B1 => n68245, B2 => 
                           n67838, ZN => n6397);
   U46981 : OAI22_X1 port map( A1 => n67845, A2 => n63027, B1 => n68248, B2 => 
                           n67838, ZN => n6398);
   U46982 : OAI22_X1 port map( A1 => n67756, A2 => n63367, B1 => n68239, B2 => 
                           n67749, ZN => n5947);
   U46983 : OAI22_X1 port map( A1 => n67756, A2 => n63366, B1 => n68242, B2 => 
                           n67749, ZN => n5948);
   U46984 : OAI22_X1 port map( A1 => n67756, A2 => n63365, B1 => n68245, B2 => 
                           n67749, ZN => n5949);
   U46985 : OAI22_X1 port map( A1 => n67756, A2 => n63363, B1 => n68248, B2 => 
                           n67749, ZN => n5950);
   U46986 : OAI22_X1 port map( A1 => n67743, A2 => n63434, B1 => n68240, B2 => 
                           n67736, ZN => n5883);
   U46987 : OAI22_X1 port map( A1 => n67743, A2 => n63433, B1 => n68243, B2 => 
                           n67736, ZN => n5884);
   U46988 : OAI22_X1 port map( A1 => n67743, A2 => n63432, B1 => n68246, B2 => 
                           n67736, ZN => n5885);
   U46989 : OAI22_X1 port map( A1 => n67743, A2 => n63430, B1 => n68249, B2 => 
                           n67736, ZN => n5886);
   U46990 : OAI22_X1 port map( A1 => n67884, A2 => n62831, B1 => n68239, B2 => 
                           n67877, ZN => n6587);
   U46991 : OAI22_X1 port map( A1 => n67884, A2 => n62830, B1 => n68242, B2 => 
                           n67877, ZN => n6588);
   U46992 : OAI22_X1 port map( A1 => n67884, A2 => n62829, B1 => n68245, B2 => 
                           n67877, ZN => n6589);
   U46993 : OAI22_X1 port map( A1 => n67884, A2 => n62827, B1 => n68248, B2 => 
                           n67877, ZN => n6590);
   U46994 : OAI22_X1 port map( A1 => n68038, A2 => n62162, B1 => n68238, B2 => 
                           n68031, ZN => n7355);
   U46995 : OAI22_X1 port map( A1 => n68038, A2 => n62161, B1 => n68241, B2 => 
                           n68031, ZN => n7356);
   U46996 : OAI22_X1 port map( A1 => n68038, A2 => n62160, B1 => n68244, B2 => 
                           n68031, ZN => n7357);
   U46997 : OAI22_X1 port map( A1 => n68038, A2 => n62158, B1 => n68247, B2 => 
                           n68031, ZN => n7358);
   U46998 : OAI22_X1 port map( A1 => n68025, A2 => n62229, B1 => n68238, B2 => 
                           n68018, ZN => n7291);
   U46999 : OAI22_X1 port map( A1 => n68025, A2 => n62228, B1 => n68241, B2 => 
                           n68018, ZN => n7292);
   U47000 : OAI22_X1 port map( A1 => n68025, A2 => n62227, B1 => n68244, B2 => 
                           n68018, ZN => n7293);
   U47001 : OAI22_X1 port map( A1 => n68025, A2 => n62225, B1 => n68247, B2 => 
                           n68018, ZN => n7294);
   U47002 : OAI22_X1 port map( A1 => n67999, A2 => n62362, B1 => n68238, B2 => 
                           n67992, ZN => n7163);
   U47003 : OAI22_X1 port map( A1 => n67999, A2 => n62361, B1 => n68241, B2 => 
                           n67992, ZN => n7164);
   U47004 : OAI22_X1 port map( A1 => n67999, A2 => n62360, B1 => n68244, B2 => 
                           n67992, ZN => n7165);
   U47005 : OAI22_X1 port map( A1 => n67999, A2 => n62358, B1 => n68247, B2 => 
                           n67992, ZN => n7166);
   U47006 : OAI22_X1 port map( A1 => n67820, A2 => n63100, B1 => n68239, B2 => 
                           n67813, ZN => n6267);
   U47007 : OAI22_X1 port map( A1 => n67820, A2 => n63099, B1 => n68242, B2 => 
                           n67813, ZN => n6268);
   U47008 : OAI22_X1 port map( A1 => n67820, A2 => n63098, B1 => n68245, B2 => 
                           n67813, ZN => n6269);
   U47009 : OAI22_X1 port map( A1 => n67820, A2 => n63096, B1 => n68248, B2 => 
                           n67813, ZN => n6270);
   U47010 : OAI22_X1 port map( A1 => n67692, A2 => n63637, B1 => n68240, B2 => 
                           n67685, ZN => n5627);
   U47011 : OAI22_X1 port map( A1 => n67692, A2 => n63636, B1 => n68243, B2 => 
                           n67685, ZN => n5628);
   U47012 : OAI22_X1 port map( A1 => n67692, A2 => n63635, B1 => n68246, B2 => 
                           n67685, ZN => n5629);
   U47013 : OAI22_X1 port map( A1 => n67692, A2 => n63633, B1 => n68249, B2 => 
                           n67685, ZN => n5630);
   U47014 : OAI22_X1 port map( A1 => n67871, A2 => n62897, B1 => n68239, B2 => 
                           n67864, ZN => n6523);
   U47015 : OAI22_X1 port map( A1 => n67871, A2 => n62896, B1 => n68242, B2 => 
                           n67864, ZN => n6524);
   U47016 : OAI22_X1 port map( A1 => n67871, A2 => n62895, B1 => n68245, B2 => 
                           n67864, ZN => n6525);
   U47017 : OAI22_X1 port map( A1 => n67871, A2 => n62893, B1 => n68248, B2 => 
                           n67864, ZN => n6526);
   U47018 : OAI22_X1 port map( A1 => n67922, A2 => n62701, B1 => n68238, B2 => 
                           n67915, ZN => n6779);
   U47019 : OAI22_X1 port map( A1 => n67922, A2 => n62700, B1 => n68241, B2 => 
                           n67915, ZN => n6780);
   U47020 : OAI22_X1 port map( A1 => n67922, A2 => n62699, B1 => n68244, B2 => 
                           n67915, ZN => n6781);
   U47021 : OAI22_X1 port map( A1 => n67922, A2 => n62697, B1 => n68247, B2 => 
                           n67915, ZN => n6782);
   U47022 : OAI22_X1 port map( A1 => n67986, A2 => n62428, B1 => n68238, B2 => 
                           n67979, ZN => n7099);
   U47023 : OAI22_X1 port map( A1 => n67986, A2 => n62427, B1 => n68241, B2 => 
                           n67979, ZN => n7100);
   U47024 : OAI22_X1 port map( A1 => n67986, A2 => n62426, B1 => n68244, B2 => 
                           n67979, ZN => n7101);
   U47025 : OAI22_X1 port map( A1 => n67986, A2 => n62424, B1 => n68247, B2 => 
                           n67979, ZN => n7102);
   U47026 : OAI22_X1 port map( A1 => n67769, A2 => n63301, B1 => n68239, B2 => 
                           n67762, ZN => n6011);
   U47027 : OAI22_X1 port map( A1 => n67769, A2 => n63300, B1 => n68242, B2 => 
                           n67762, ZN => n6012);
   U47028 : OAI22_X1 port map( A1 => n67769, A2 => n63299, B1 => n68245, B2 => 
                           n67762, ZN => n6013);
   U47029 : OAI22_X1 port map( A1 => n67769, A2 => n63297, B1 => n68248, B2 => 
                           n67762, ZN => n6014);
   U47030 : OAI22_X1 port map( A1 => n67718, A2 => n63505, B1 => n68240, B2 => 
                           n67711, ZN => n5755);
   U47031 : OAI22_X1 port map( A1 => n67718, A2 => n63504, B1 => n68243, B2 => 
                           n67711, ZN => n5756);
   U47032 : OAI22_X1 port map( A1 => n67718, A2 => n63503, B1 => n68246, B2 => 
                           n67711, ZN => n5757);
   U47033 : OAI22_X1 port map( A1 => n67718, A2 => n63501, B1 => n68249, B2 => 
                           n67711, ZN => n5758);
   U47034 : OAI22_X1 port map( A1 => n67705, A2 => n63571, B1 => n68240, B2 => 
                           n67698, ZN => n5691);
   U47035 : OAI22_X1 port map( A1 => n67705, A2 => n63570, B1 => n68243, B2 => 
                           n67698, ZN => n5692);
   U47036 : OAI22_X1 port map( A1 => n67705, A2 => n63569, B1 => n68246, B2 => 
                           n67698, ZN => n5693);
   U47037 : OAI22_X1 port map( A1 => n67705, A2 => n63567, B1 => n68249, B2 => 
                           n67698, ZN => n5694);
   U47038 : NAND2_X1 port map( A1 => n66280, A2 => n66278, ZN => n65123);
   U47039 : OAI22_X1 port map( A1 => n67739, A2 => n63494, B1 => n68060, B2 => 
                           n67731, ZN => n5823);
   U47040 : OAI22_X1 port map( A1 => n67739, A2 => n63493, B1 => n68063, B2 => 
                           n67731, ZN => n5824);
   U47041 : OAI22_X1 port map( A1 => n67739, A2 => n63492, B1 => n68066, B2 => 
                           n67731, ZN => n5825);
   U47042 : OAI22_X1 port map( A1 => n67739, A2 => n63491, B1 => n68069, B2 => 
                           n67731, ZN => n5826);
   U47043 : OAI22_X1 port map( A1 => n67739, A2 => n63490, B1 => n68072, B2 => 
                           n67731, ZN => n5827);
   U47044 : OAI22_X1 port map( A1 => n67739, A2 => n63489, B1 => n68075, B2 => 
                           n67731, ZN => n5828);
   U47045 : OAI22_X1 port map( A1 => n67739, A2 => n63488, B1 => n68078, B2 => 
                           n67731, ZN => n5829);
   U47046 : OAI22_X1 port map( A1 => n67739, A2 => n63487, B1 => n68081, B2 => 
                           n67731, ZN => n5830);
   U47047 : OAI22_X1 port map( A1 => n67739, A2 => n63486, B1 => n68084, B2 => 
                           n67731, ZN => n5831);
   U47048 : OAI22_X1 port map( A1 => n67739, A2 => n63485, B1 => n68087, B2 => 
                           n67731, ZN => n5832);
   U47049 : OAI22_X1 port map( A1 => n67739, A2 => n63484, B1 => n68090, B2 => 
                           n67731, ZN => n5833);
   U47050 : OAI22_X1 port map( A1 => n67739, A2 => n63483, B1 => n68093, B2 => 
                           n67731, ZN => n5834);
   U47051 : OAI22_X1 port map( A1 => n67740, A2 => n63482, B1 => n68096, B2 => 
                           n67732, ZN => n5835);
   U47052 : OAI22_X1 port map( A1 => n67740, A2 => n63481, B1 => n68099, B2 => 
                           n67732, ZN => n5836);
   U47053 : OAI22_X1 port map( A1 => n67740, A2 => n63480, B1 => n68102, B2 => 
                           n67732, ZN => n5837);
   U47054 : OAI22_X1 port map( A1 => n67740, A2 => n63479, B1 => n68105, B2 => 
                           n67732, ZN => n5838);
   U47055 : OAI22_X1 port map( A1 => n67740, A2 => n63478, B1 => n68108, B2 => 
                           n67732, ZN => n5839);
   U47056 : OAI22_X1 port map( A1 => n67740, A2 => n63477, B1 => n68111, B2 => 
                           n67732, ZN => n5840);
   U47057 : OAI22_X1 port map( A1 => n67740, A2 => n63476, B1 => n68114, B2 => 
                           n67732, ZN => n5841);
   U47058 : OAI22_X1 port map( A1 => n67740, A2 => n63475, B1 => n68117, B2 => 
                           n67732, ZN => n5842);
   U47059 : OAI22_X1 port map( A1 => n67740, A2 => n63474, B1 => n68120, B2 => 
                           n67732, ZN => n5843);
   U47060 : OAI22_X1 port map( A1 => n67740, A2 => n63473, B1 => n68123, B2 => 
                           n67732, ZN => n5844);
   U47061 : OAI22_X1 port map( A1 => n67740, A2 => n63472, B1 => n68126, B2 => 
                           n67732, ZN => n5845);
   U47062 : OAI22_X1 port map( A1 => n67740, A2 => n63471, B1 => n68129, B2 => 
                           n67732, ZN => n5846);
   U47063 : OAI22_X1 port map( A1 => n67740, A2 => n63470, B1 => n68132, B2 => 
                           n67733, ZN => n5847);
   U47064 : OAI22_X1 port map( A1 => n67741, A2 => n63469, B1 => n68135, B2 => 
                           n67733, ZN => n5848);
   U47065 : OAI22_X1 port map( A1 => n67741, A2 => n63468, B1 => n68138, B2 => 
                           n67733, ZN => n5849);
   U47066 : OAI22_X1 port map( A1 => n67741, A2 => n63467, B1 => n68141, B2 => 
                           n67733, ZN => n5850);
   U47067 : OAI22_X1 port map( A1 => n67741, A2 => n63466, B1 => n68144, B2 => 
                           n67733, ZN => n5851);
   U47068 : OAI22_X1 port map( A1 => n67741, A2 => n63465, B1 => n68147, B2 => 
                           n67733, ZN => n5852);
   U47069 : OAI22_X1 port map( A1 => n67741, A2 => n63464, B1 => n68150, B2 => 
                           n67733, ZN => n5853);
   U47070 : OAI22_X1 port map( A1 => n67741, A2 => n63463, B1 => n68153, B2 => 
                           n67733, ZN => n5854);
   U47071 : OAI22_X1 port map( A1 => n67741, A2 => n63462, B1 => n68156, B2 => 
                           n67733, ZN => n5855);
   U47072 : OAI22_X1 port map( A1 => n67741, A2 => n63461, B1 => n68159, B2 => 
                           n67733, ZN => n5856);
   U47073 : OAI22_X1 port map( A1 => n67741, A2 => n63460, B1 => n68162, B2 => 
                           n67733, ZN => n5857);
   U47074 : OAI22_X1 port map( A1 => n67741, A2 => n63459, B1 => n68165, B2 => 
                           n67733, ZN => n5858);
   U47075 : OAI22_X1 port map( A1 => n67741, A2 => n63458, B1 => n68168, B2 => 
                           n67734, ZN => n5859);
   U47076 : OAI22_X1 port map( A1 => n67741, A2 => n63457, B1 => n68171, B2 => 
                           n67734, ZN => n5860);
   U47077 : OAI22_X1 port map( A1 => n67742, A2 => n63456, B1 => n68174, B2 => 
                           n67734, ZN => n5861);
   U47078 : OAI22_X1 port map( A1 => n67742, A2 => n63455, B1 => n68177, B2 => 
                           n67734, ZN => n5862);
   U47079 : OAI22_X1 port map( A1 => n67742, A2 => n63454, B1 => n68180, B2 => 
                           n67734, ZN => n5863);
   U47080 : OAI22_X1 port map( A1 => n67742, A2 => n63453, B1 => n68183, B2 => 
                           n67734, ZN => n5864);
   U47081 : OAI22_X1 port map( A1 => n67742, A2 => n63452, B1 => n68186, B2 => 
                           n67734, ZN => n5865);
   U47082 : OAI22_X1 port map( A1 => n67742, A2 => n63451, B1 => n68189, B2 => 
                           n67734, ZN => n5866);
   U47083 : OAI22_X1 port map( A1 => n67742, A2 => n63450, B1 => n68192, B2 => 
                           n67734, ZN => n5867);
   U47084 : OAI22_X1 port map( A1 => n67742, A2 => n63449, B1 => n68195, B2 => 
                           n67734, ZN => n5868);
   U47085 : OAI22_X1 port map( A1 => n67742, A2 => n63448, B1 => n68198, B2 => 
                           n67734, ZN => n5869);
   U47086 : OAI22_X1 port map( A1 => n67742, A2 => n63447, B1 => n68201, B2 => 
                           n67734, ZN => n5870);
   U47087 : OAI22_X1 port map( A1 => n67742, A2 => n63446, B1 => n68204, B2 => 
                           n67735, ZN => n5871);
   U47088 : OAI22_X1 port map( A1 => n67742, A2 => n63445, B1 => n68207, B2 => 
                           n67735, ZN => n5872);
   U47089 : OAI22_X1 port map( A1 => n67742, A2 => n63444, B1 => n68210, B2 => 
                           n67735, ZN => n5873);
   U47090 : OAI22_X1 port map( A1 => n67743, A2 => n63443, B1 => n68213, B2 => 
                           n67735, ZN => n5874);
   U47091 : OAI22_X1 port map( A1 => n67743, A2 => n63442, B1 => n68216, B2 => 
                           n67735, ZN => n5875);
   U47092 : OAI22_X1 port map( A1 => n67743, A2 => n63441, B1 => n68219, B2 => 
                           n67735, ZN => n5876);
   U47093 : OAI22_X1 port map( A1 => n67743, A2 => n63440, B1 => n68222, B2 => 
                           n67735, ZN => n5877);
   U47094 : OAI22_X1 port map( A1 => n67743, A2 => n63439, B1 => n68225, B2 => 
                           n67735, ZN => n5878);
   U47095 : OAI22_X1 port map( A1 => n67743, A2 => n63438, B1 => n68228, B2 => 
                           n67735, ZN => n5879);
   U47096 : OAI22_X1 port map( A1 => n67743, A2 => n63437, B1 => n68231, B2 => 
                           n67735, ZN => n5880);
   U47097 : OAI22_X1 port map( A1 => n67743, A2 => n63436, B1 => n68234, B2 => 
                           n67735, ZN => n5881);
   U47098 : OAI22_X1 port map( A1 => n67743, A2 => n63435, B1 => n68237, B2 => 
                           n67735, ZN => n5882);
   U47099 : OAI22_X1 port map( A1 => n67688, A2 => n63697, B1 => n68060, B2 => 
                           n67680, ZN => n5567);
   U47100 : OAI22_X1 port map( A1 => n67688, A2 => n63696, B1 => n68063, B2 => 
                           n67680, ZN => n5568);
   U47101 : OAI22_X1 port map( A1 => n67688, A2 => n63695, B1 => n68066, B2 => 
                           n67680, ZN => n5569);
   U47102 : OAI22_X1 port map( A1 => n67688, A2 => n63694, B1 => n68069, B2 => 
                           n67680, ZN => n5570);
   U47103 : OAI22_X1 port map( A1 => n67688, A2 => n63693, B1 => n68072, B2 => 
                           n67680, ZN => n5571);
   U47104 : OAI22_X1 port map( A1 => n67688, A2 => n63692, B1 => n68075, B2 => 
                           n67680, ZN => n5572);
   U47105 : OAI22_X1 port map( A1 => n67688, A2 => n63691, B1 => n68078, B2 => 
                           n67680, ZN => n5573);
   U47106 : OAI22_X1 port map( A1 => n67688, A2 => n63690, B1 => n68081, B2 => 
                           n67680, ZN => n5574);
   U47107 : OAI22_X1 port map( A1 => n67688, A2 => n63689, B1 => n68084, B2 => 
                           n67680, ZN => n5575);
   U47108 : OAI22_X1 port map( A1 => n67688, A2 => n63688, B1 => n68087, B2 => 
                           n67680, ZN => n5576);
   U47109 : OAI22_X1 port map( A1 => n67688, A2 => n63687, B1 => n68090, B2 => 
                           n67680, ZN => n5577);
   U47110 : OAI22_X1 port map( A1 => n67688, A2 => n63686, B1 => n68093, B2 => 
                           n67680, ZN => n5578);
   U47111 : OAI22_X1 port map( A1 => n67689, A2 => n63685, B1 => n68096, B2 => 
                           n67681, ZN => n5579);
   U47112 : OAI22_X1 port map( A1 => n67689, A2 => n63684, B1 => n68099, B2 => 
                           n67681, ZN => n5580);
   U47113 : OAI22_X1 port map( A1 => n67689, A2 => n63683, B1 => n68102, B2 => 
                           n67681, ZN => n5581);
   U47114 : OAI22_X1 port map( A1 => n67689, A2 => n63682, B1 => n68105, B2 => 
                           n67681, ZN => n5582);
   U47115 : OAI22_X1 port map( A1 => n67689, A2 => n63681, B1 => n68108, B2 => 
                           n67681, ZN => n5583);
   U47116 : OAI22_X1 port map( A1 => n67689, A2 => n63680, B1 => n68111, B2 => 
                           n67681, ZN => n5584);
   U47117 : OAI22_X1 port map( A1 => n67689, A2 => n63679, B1 => n68114, B2 => 
                           n67681, ZN => n5585);
   U47118 : OAI22_X1 port map( A1 => n67689, A2 => n63678, B1 => n68117, B2 => 
                           n67681, ZN => n5586);
   U47119 : OAI22_X1 port map( A1 => n67689, A2 => n63677, B1 => n68120, B2 => 
                           n67681, ZN => n5587);
   U47120 : OAI22_X1 port map( A1 => n67689, A2 => n63676, B1 => n68123, B2 => 
                           n67681, ZN => n5588);
   U47121 : OAI22_X1 port map( A1 => n67689, A2 => n63675, B1 => n68126, B2 => 
                           n67681, ZN => n5589);
   U47122 : OAI22_X1 port map( A1 => n67689, A2 => n63674, B1 => n68129, B2 => 
                           n67681, ZN => n5590);
   U47123 : OAI22_X1 port map( A1 => n67689, A2 => n63673, B1 => n68132, B2 => 
                           n67682, ZN => n5591);
   U47124 : OAI22_X1 port map( A1 => n67690, A2 => n63672, B1 => n68135, B2 => 
                           n67682, ZN => n5592);
   U47125 : OAI22_X1 port map( A1 => n67690, A2 => n63671, B1 => n68138, B2 => 
                           n67682, ZN => n5593);
   U47126 : OAI22_X1 port map( A1 => n67690, A2 => n63670, B1 => n68141, B2 => 
                           n67682, ZN => n5594);
   U47127 : OAI22_X1 port map( A1 => n67690, A2 => n63669, B1 => n68144, B2 => 
                           n67682, ZN => n5595);
   U47128 : OAI22_X1 port map( A1 => n67690, A2 => n63668, B1 => n68147, B2 => 
                           n67682, ZN => n5596);
   U47129 : OAI22_X1 port map( A1 => n67690, A2 => n63667, B1 => n68150, B2 => 
                           n67682, ZN => n5597);
   U47130 : OAI22_X1 port map( A1 => n67690, A2 => n63666, B1 => n68153, B2 => 
                           n67682, ZN => n5598);
   U47131 : OAI22_X1 port map( A1 => n67690, A2 => n63665, B1 => n68156, B2 => 
                           n67682, ZN => n5599);
   U47132 : OAI22_X1 port map( A1 => n67690, A2 => n63664, B1 => n68159, B2 => 
                           n67682, ZN => n5600);
   U47133 : OAI22_X1 port map( A1 => n67690, A2 => n63663, B1 => n68162, B2 => 
                           n67682, ZN => n5601);
   U47134 : OAI22_X1 port map( A1 => n67690, A2 => n63662, B1 => n68165, B2 => 
                           n67682, ZN => n5602);
   U47135 : OAI22_X1 port map( A1 => n67690, A2 => n63661, B1 => n68168, B2 => 
                           n67683, ZN => n5603);
   U47136 : OAI22_X1 port map( A1 => n67690, A2 => n63660, B1 => n68171, B2 => 
                           n67683, ZN => n5604);
   U47137 : OAI22_X1 port map( A1 => n67691, A2 => n63659, B1 => n68174, B2 => 
                           n67683, ZN => n5605);
   U47138 : OAI22_X1 port map( A1 => n67691, A2 => n63658, B1 => n68177, B2 => 
                           n67683, ZN => n5606);
   U47139 : OAI22_X1 port map( A1 => n67691, A2 => n63657, B1 => n68180, B2 => 
                           n67683, ZN => n5607);
   U47140 : OAI22_X1 port map( A1 => n67691, A2 => n63656, B1 => n68183, B2 => 
                           n67683, ZN => n5608);
   U47141 : OAI22_X1 port map( A1 => n67691, A2 => n63655, B1 => n68186, B2 => 
                           n67683, ZN => n5609);
   U47142 : OAI22_X1 port map( A1 => n67691, A2 => n63654, B1 => n68189, B2 => 
                           n67683, ZN => n5610);
   U47143 : OAI22_X1 port map( A1 => n67691, A2 => n63653, B1 => n68192, B2 => 
                           n67683, ZN => n5611);
   U47144 : OAI22_X1 port map( A1 => n67691, A2 => n63652, B1 => n68195, B2 => 
                           n67683, ZN => n5612);
   U47145 : OAI22_X1 port map( A1 => n67691, A2 => n63651, B1 => n68198, B2 => 
                           n67683, ZN => n5613);
   U47146 : OAI22_X1 port map( A1 => n67691, A2 => n63650, B1 => n68201, B2 => 
                           n67683, ZN => n5614);
   U47147 : OAI22_X1 port map( A1 => n67691, A2 => n63649, B1 => n68204, B2 => 
                           n67684, ZN => n5615);
   U47148 : OAI22_X1 port map( A1 => n67691, A2 => n63648, B1 => n68207, B2 => 
                           n67684, ZN => n5616);
   U47149 : OAI22_X1 port map( A1 => n67691, A2 => n63647, B1 => n68210, B2 => 
                           n67684, ZN => n5617);
   U47150 : OAI22_X1 port map( A1 => n67692, A2 => n63646, B1 => n68213, B2 => 
                           n67684, ZN => n5618);
   U47151 : OAI22_X1 port map( A1 => n67692, A2 => n63645, B1 => n68216, B2 => 
                           n67684, ZN => n5619);
   U47152 : OAI22_X1 port map( A1 => n67692, A2 => n63644, B1 => n68219, B2 => 
                           n67684, ZN => n5620);
   U47153 : OAI22_X1 port map( A1 => n67692, A2 => n63643, B1 => n68222, B2 => 
                           n67684, ZN => n5621);
   U47154 : OAI22_X1 port map( A1 => n67692, A2 => n63642, B1 => n68225, B2 => 
                           n67684, ZN => n5622);
   U47155 : OAI22_X1 port map( A1 => n67692, A2 => n63641, B1 => n68228, B2 => 
                           n67684, ZN => n5623);
   U47156 : OAI22_X1 port map( A1 => n67692, A2 => n63640, B1 => n68231, B2 => 
                           n67684, ZN => n5624);
   U47157 : OAI22_X1 port map( A1 => n67692, A2 => n63639, B1 => n68234, B2 => 
                           n67684, ZN => n5625);
   U47158 : OAI22_X1 port map( A1 => n67692, A2 => n63638, B1 => n68237, B2 => 
                           n67684, ZN => n5626);
   U47159 : OAI22_X1 port map( A1 => n67714, A2 => n63565, B1 => n68060, B2 => 
                           n67706, ZN => n5695);
   U47160 : OAI22_X1 port map( A1 => n67714, A2 => n63564, B1 => n68063, B2 => 
                           n67706, ZN => n5696);
   U47161 : OAI22_X1 port map( A1 => n67714, A2 => n63563, B1 => n68066, B2 => 
                           n67706, ZN => n5697);
   U47162 : OAI22_X1 port map( A1 => n67714, A2 => n63562, B1 => n68069, B2 => 
                           n67706, ZN => n5698);
   U47163 : OAI22_X1 port map( A1 => n67714, A2 => n63561, B1 => n68072, B2 => 
                           n67706, ZN => n5699);
   U47164 : OAI22_X1 port map( A1 => n67714, A2 => n63560, B1 => n68075, B2 => 
                           n67706, ZN => n5700);
   U47165 : OAI22_X1 port map( A1 => n67714, A2 => n63559, B1 => n68078, B2 => 
                           n67706, ZN => n5701);
   U47166 : OAI22_X1 port map( A1 => n67714, A2 => n63558, B1 => n68081, B2 => 
                           n67706, ZN => n5702);
   U47167 : OAI22_X1 port map( A1 => n67714, A2 => n63557, B1 => n68084, B2 => 
                           n67706, ZN => n5703);
   U47168 : OAI22_X1 port map( A1 => n67714, A2 => n63556, B1 => n68087, B2 => 
                           n67706, ZN => n5704);
   U47169 : OAI22_X1 port map( A1 => n67714, A2 => n63555, B1 => n68090, B2 => 
                           n67706, ZN => n5705);
   U47170 : OAI22_X1 port map( A1 => n67714, A2 => n63554, B1 => n68093, B2 => 
                           n67706, ZN => n5706);
   U47171 : OAI22_X1 port map( A1 => n67715, A2 => n63553, B1 => n68096, B2 => 
                           n67707, ZN => n5707);
   U47172 : OAI22_X1 port map( A1 => n67715, A2 => n63552, B1 => n68099, B2 => 
                           n67707, ZN => n5708);
   U47173 : OAI22_X1 port map( A1 => n67715, A2 => n63551, B1 => n68102, B2 => 
                           n67707, ZN => n5709);
   U47174 : OAI22_X1 port map( A1 => n67715, A2 => n63550, B1 => n68105, B2 => 
                           n67707, ZN => n5710);
   U47175 : OAI22_X1 port map( A1 => n67715, A2 => n63549, B1 => n68108, B2 => 
                           n67707, ZN => n5711);
   U47176 : OAI22_X1 port map( A1 => n67715, A2 => n63548, B1 => n68111, B2 => 
                           n67707, ZN => n5712);
   U47177 : OAI22_X1 port map( A1 => n67715, A2 => n63547, B1 => n68114, B2 => 
                           n67707, ZN => n5713);
   U47178 : OAI22_X1 port map( A1 => n67715, A2 => n63546, B1 => n68117, B2 => 
                           n67707, ZN => n5714);
   U47179 : OAI22_X1 port map( A1 => n67715, A2 => n63545, B1 => n68120, B2 => 
                           n67707, ZN => n5715);
   U47180 : OAI22_X1 port map( A1 => n67715, A2 => n63544, B1 => n68123, B2 => 
                           n67707, ZN => n5716);
   U47181 : OAI22_X1 port map( A1 => n67715, A2 => n63543, B1 => n68126, B2 => 
                           n67707, ZN => n5717);
   U47182 : OAI22_X1 port map( A1 => n67715, A2 => n63542, B1 => n68129, B2 => 
                           n67707, ZN => n5718);
   U47183 : OAI22_X1 port map( A1 => n67715, A2 => n63541, B1 => n68132, B2 => 
                           n67708, ZN => n5719);
   U47184 : OAI22_X1 port map( A1 => n67716, A2 => n63540, B1 => n68135, B2 => 
                           n67708, ZN => n5720);
   U47185 : OAI22_X1 port map( A1 => n67716, A2 => n63539, B1 => n68138, B2 => 
                           n67708, ZN => n5721);
   U47186 : OAI22_X1 port map( A1 => n67716, A2 => n63538, B1 => n68141, B2 => 
                           n67708, ZN => n5722);
   U47187 : OAI22_X1 port map( A1 => n67716, A2 => n63537, B1 => n68144, B2 => 
                           n67708, ZN => n5723);
   U47188 : OAI22_X1 port map( A1 => n67716, A2 => n63536, B1 => n68147, B2 => 
                           n67708, ZN => n5724);
   U47189 : OAI22_X1 port map( A1 => n67716, A2 => n63535, B1 => n68150, B2 => 
                           n67708, ZN => n5725);
   U47190 : OAI22_X1 port map( A1 => n67716, A2 => n63534, B1 => n68153, B2 => 
                           n67708, ZN => n5726);
   U47191 : OAI22_X1 port map( A1 => n67716, A2 => n63533, B1 => n68156, B2 => 
                           n67708, ZN => n5727);
   U47192 : OAI22_X1 port map( A1 => n67716, A2 => n63532, B1 => n68159, B2 => 
                           n67708, ZN => n5728);
   U47193 : OAI22_X1 port map( A1 => n67716, A2 => n63531, B1 => n68162, B2 => 
                           n67708, ZN => n5729);
   U47194 : OAI22_X1 port map( A1 => n67716, A2 => n63530, B1 => n68165, B2 => 
                           n67708, ZN => n5730);
   U47195 : OAI22_X1 port map( A1 => n67716, A2 => n63529, B1 => n68168, B2 => 
                           n67709, ZN => n5731);
   U47196 : OAI22_X1 port map( A1 => n67716, A2 => n63528, B1 => n68171, B2 => 
                           n67709, ZN => n5732);
   U47197 : OAI22_X1 port map( A1 => n67717, A2 => n63527, B1 => n68174, B2 => 
                           n67709, ZN => n5733);
   U47198 : OAI22_X1 port map( A1 => n67717, A2 => n63526, B1 => n68177, B2 => 
                           n67709, ZN => n5734);
   U47199 : OAI22_X1 port map( A1 => n67717, A2 => n63525, B1 => n68180, B2 => 
                           n67709, ZN => n5735);
   U47200 : OAI22_X1 port map( A1 => n67717, A2 => n63524, B1 => n68183, B2 => 
                           n67709, ZN => n5736);
   U47201 : OAI22_X1 port map( A1 => n67717, A2 => n63523, B1 => n68186, B2 => 
                           n67709, ZN => n5737);
   U47202 : OAI22_X1 port map( A1 => n67717, A2 => n63522, B1 => n68189, B2 => 
                           n67709, ZN => n5738);
   U47203 : OAI22_X1 port map( A1 => n67717, A2 => n63521, B1 => n68192, B2 => 
                           n67709, ZN => n5739);
   U47204 : OAI22_X1 port map( A1 => n67717, A2 => n63520, B1 => n68195, B2 => 
                           n67709, ZN => n5740);
   U47205 : OAI22_X1 port map( A1 => n67717, A2 => n63519, B1 => n68198, B2 => 
                           n67709, ZN => n5741);
   U47206 : OAI22_X1 port map( A1 => n67717, A2 => n63518, B1 => n68201, B2 => 
                           n67709, ZN => n5742);
   U47207 : OAI22_X1 port map( A1 => n67717, A2 => n63517, B1 => n68204, B2 => 
                           n67710, ZN => n5743);
   U47208 : OAI22_X1 port map( A1 => n67717, A2 => n63516, B1 => n68207, B2 => 
                           n67710, ZN => n5744);
   U47209 : OAI22_X1 port map( A1 => n67717, A2 => n63515, B1 => n68210, B2 => 
                           n67710, ZN => n5745);
   U47210 : OAI22_X1 port map( A1 => n67718, A2 => n63514, B1 => n68213, B2 => 
                           n67710, ZN => n5746);
   U47211 : OAI22_X1 port map( A1 => n67718, A2 => n63513, B1 => n68216, B2 => 
                           n67710, ZN => n5747);
   U47212 : OAI22_X1 port map( A1 => n67718, A2 => n63512, B1 => n68219, B2 => 
                           n67710, ZN => n5748);
   U47213 : OAI22_X1 port map( A1 => n67718, A2 => n63511, B1 => n68222, B2 => 
                           n67710, ZN => n5749);
   U47214 : OAI22_X1 port map( A1 => n67718, A2 => n63510, B1 => n68225, B2 => 
                           n67710, ZN => n5750);
   U47215 : OAI22_X1 port map( A1 => n67718, A2 => n63509, B1 => n68228, B2 => 
                           n67710, ZN => n5751);
   U47216 : OAI22_X1 port map( A1 => n67718, A2 => n63508, B1 => n68231, B2 => 
                           n67710, ZN => n5752);
   U47217 : OAI22_X1 port map( A1 => n67718, A2 => n63507, B1 => n68234, B2 => 
                           n67710, ZN => n5753);
   U47218 : OAI22_X1 port map( A1 => n67718, A2 => n63506, B1 => n68237, B2 => 
                           n67710, ZN => n5754);
   U47219 : OAI22_X1 port map( A1 => n67701, A2 => n63631, B1 => n68060, B2 => 
                           n67693, ZN => n5631);
   U47220 : OAI22_X1 port map( A1 => n67701, A2 => n63630, B1 => n68063, B2 => 
                           n67693, ZN => n5632);
   U47221 : OAI22_X1 port map( A1 => n67701, A2 => n63629, B1 => n68066, B2 => 
                           n67693, ZN => n5633);
   U47222 : OAI22_X1 port map( A1 => n67701, A2 => n63628, B1 => n68069, B2 => 
                           n67693, ZN => n5634);
   U47223 : OAI22_X1 port map( A1 => n67701, A2 => n63627, B1 => n68072, B2 => 
                           n67693, ZN => n5635);
   U47224 : OAI22_X1 port map( A1 => n67701, A2 => n63626, B1 => n68075, B2 => 
                           n67693, ZN => n5636);
   U47225 : OAI22_X1 port map( A1 => n67701, A2 => n63625, B1 => n68078, B2 => 
                           n67693, ZN => n5637);
   U47226 : OAI22_X1 port map( A1 => n67701, A2 => n63624, B1 => n68081, B2 => 
                           n67693, ZN => n5638);
   U47227 : OAI22_X1 port map( A1 => n67701, A2 => n63623, B1 => n68084, B2 => 
                           n67693, ZN => n5639);
   U47228 : OAI22_X1 port map( A1 => n67701, A2 => n63622, B1 => n68087, B2 => 
                           n67693, ZN => n5640);
   U47229 : OAI22_X1 port map( A1 => n67701, A2 => n63621, B1 => n68090, B2 => 
                           n67693, ZN => n5641);
   U47230 : OAI22_X1 port map( A1 => n67701, A2 => n63620, B1 => n68093, B2 => 
                           n67693, ZN => n5642);
   U47231 : OAI22_X1 port map( A1 => n67702, A2 => n63619, B1 => n68096, B2 => 
                           n67694, ZN => n5643);
   U47232 : OAI22_X1 port map( A1 => n67702, A2 => n63618, B1 => n68099, B2 => 
                           n67694, ZN => n5644);
   U47233 : OAI22_X1 port map( A1 => n67702, A2 => n63617, B1 => n68102, B2 => 
                           n67694, ZN => n5645);
   U47234 : OAI22_X1 port map( A1 => n67702, A2 => n63616, B1 => n68105, B2 => 
                           n67694, ZN => n5646);
   U47235 : OAI22_X1 port map( A1 => n67702, A2 => n63615, B1 => n68108, B2 => 
                           n67694, ZN => n5647);
   U47236 : OAI22_X1 port map( A1 => n67702, A2 => n63614, B1 => n68111, B2 => 
                           n67694, ZN => n5648);
   U47237 : OAI22_X1 port map( A1 => n67702, A2 => n63613, B1 => n68114, B2 => 
                           n67694, ZN => n5649);
   U47238 : OAI22_X1 port map( A1 => n67702, A2 => n63612, B1 => n68117, B2 => 
                           n67694, ZN => n5650);
   U47239 : OAI22_X1 port map( A1 => n67702, A2 => n63611, B1 => n68120, B2 => 
                           n67694, ZN => n5651);
   U47240 : OAI22_X1 port map( A1 => n67702, A2 => n63610, B1 => n68123, B2 => 
                           n67694, ZN => n5652);
   U47241 : OAI22_X1 port map( A1 => n67702, A2 => n63609, B1 => n68126, B2 => 
                           n67694, ZN => n5653);
   U47242 : OAI22_X1 port map( A1 => n67702, A2 => n63608, B1 => n68129, B2 => 
                           n67694, ZN => n5654);
   U47243 : OAI22_X1 port map( A1 => n67702, A2 => n63607, B1 => n68132, B2 => 
                           n67695, ZN => n5655);
   U47244 : OAI22_X1 port map( A1 => n67703, A2 => n63606, B1 => n68135, B2 => 
                           n67695, ZN => n5656);
   U47245 : OAI22_X1 port map( A1 => n67703, A2 => n63605, B1 => n68138, B2 => 
                           n67695, ZN => n5657);
   U47246 : OAI22_X1 port map( A1 => n67703, A2 => n63604, B1 => n68141, B2 => 
                           n67695, ZN => n5658);
   U47247 : OAI22_X1 port map( A1 => n67703, A2 => n63603, B1 => n68144, B2 => 
                           n67695, ZN => n5659);
   U47248 : OAI22_X1 port map( A1 => n67703, A2 => n63602, B1 => n68147, B2 => 
                           n67695, ZN => n5660);
   U47249 : OAI22_X1 port map( A1 => n67703, A2 => n63601, B1 => n68150, B2 => 
                           n67695, ZN => n5661);
   U47250 : OAI22_X1 port map( A1 => n67703, A2 => n63600, B1 => n68153, B2 => 
                           n67695, ZN => n5662);
   U47251 : OAI22_X1 port map( A1 => n67703, A2 => n63599, B1 => n68156, B2 => 
                           n67695, ZN => n5663);
   U47252 : OAI22_X1 port map( A1 => n67703, A2 => n63598, B1 => n68159, B2 => 
                           n67695, ZN => n5664);
   U47253 : OAI22_X1 port map( A1 => n67703, A2 => n63597, B1 => n68162, B2 => 
                           n67695, ZN => n5665);
   U47254 : OAI22_X1 port map( A1 => n67703, A2 => n63596, B1 => n68165, B2 => 
                           n67695, ZN => n5666);
   U47255 : OAI22_X1 port map( A1 => n67703, A2 => n63595, B1 => n68168, B2 => 
                           n67696, ZN => n5667);
   U47256 : OAI22_X1 port map( A1 => n67703, A2 => n63594, B1 => n68171, B2 => 
                           n67696, ZN => n5668);
   U47257 : OAI22_X1 port map( A1 => n67704, A2 => n63593, B1 => n68174, B2 => 
                           n67696, ZN => n5669);
   U47258 : OAI22_X1 port map( A1 => n67704, A2 => n63592, B1 => n68177, B2 => 
                           n67696, ZN => n5670);
   U47259 : OAI22_X1 port map( A1 => n67704, A2 => n63591, B1 => n68180, B2 => 
                           n67696, ZN => n5671);
   U47260 : OAI22_X1 port map( A1 => n67704, A2 => n63590, B1 => n68183, B2 => 
                           n67696, ZN => n5672);
   U47261 : OAI22_X1 port map( A1 => n67704, A2 => n63589, B1 => n68186, B2 => 
                           n67696, ZN => n5673);
   U47262 : OAI22_X1 port map( A1 => n67704, A2 => n63588, B1 => n68189, B2 => 
                           n67696, ZN => n5674);
   U47263 : OAI22_X1 port map( A1 => n67704, A2 => n63587, B1 => n68192, B2 => 
                           n67696, ZN => n5675);
   U47264 : OAI22_X1 port map( A1 => n67704, A2 => n63586, B1 => n68195, B2 => 
                           n67696, ZN => n5676);
   U47265 : OAI22_X1 port map( A1 => n67704, A2 => n63585, B1 => n68198, B2 => 
                           n67696, ZN => n5677);
   U47266 : OAI22_X1 port map( A1 => n67704, A2 => n63584, B1 => n68201, B2 => 
                           n67696, ZN => n5678);
   U47267 : OAI22_X1 port map( A1 => n67704, A2 => n63583, B1 => n68204, B2 => 
                           n67697, ZN => n5679);
   U47268 : OAI22_X1 port map( A1 => n67704, A2 => n63582, B1 => n68207, B2 => 
                           n67697, ZN => n5680);
   U47269 : OAI22_X1 port map( A1 => n67704, A2 => n63581, B1 => n68210, B2 => 
                           n67697, ZN => n5681);
   U47270 : OAI22_X1 port map( A1 => n67705, A2 => n63580, B1 => n68213, B2 => 
                           n67697, ZN => n5682);
   U47271 : OAI22_X1 port map( A1 => n67705, A2 => n63579, B1 => n68216, B2 => 
                           n67697, ZN => n5683);
   U47272 : OAI22_X1 port map( A1 => n67705, A2 => n63578, B1 => n68219, B2 => 
                           n67697, ZN => n5684);
   U47273 : OAI22_X1 port map( A1 => n67705, A2 => n63577, B1 => n68222, B2 => 
                           n67697, ZN => n5685);
   U47274 : OAI22_X1 port map( A1 => n67705, A2 => n63576, B1 => n68225, B2 => 
                           n67697, ZN => n5686);
   U47275 : OAI22_X1 port map( A1 => n67705, A2 => n63575, B1 => n68228, B2 => 
                           n67697, ZN => n5687);
   U47276 : OAI22_X1 port map( A1 => n67705, A2 => n63574, B1 => n68231, B2 => 
                           n67697, ZN => n5688);
   U47277 : OAI22_X1 port map( A1 => n67705, A2 => n63573, B1 => n68234, B2 => 
                           n67697, ZN => n5689);
   U47278 : OAI22_X1 port map( A1 => n67705, A2 => n63572, B1 => n68237, B2 => 
                           n67697, ZN => n5690);
   U47279 : NAND2_X1 port map( A1 => n66280, A2 => n66281, ZN => n65108);
   U47280 : NAND2_X1 port map( A1 => n66287, A2 => n66277, ZN => n65118);
   U47281 : AND2_X1 port map( A1 => n65085, A2 => n65074, ZN => n63790);
   U47282 : OAI22_X1 port map( A1 => n67943, A2 => n62691, B1 => n68058, B2 => 
                           n67935, ZN => n6847);
   U47283 : OAI22_X1 port map( A1 => n67943, A2 => n62690, B1 => n68061, B2 => 
                           n67935, ZN => n6848);
   U47284 : OAI22_X1 port map( A1 => n67943, A2 => n62689, B1 => n68064, B2 => 
                           n67935, ZN => n6849);
   U47285 : OAI22_X1 port map( A1 => n67943, A2 => n62688, B1 => n68067, B2 => 
                           n67935, ZN => n6850);
   U47286 : OAI22_X1 port map( A1 => n67943, A2 => n62687, B1 => n68070, B2 => 
                           n67935, ZN => n6851);
   U47287 : OAI22_X1 port map( A1 => n67943, A2 => n62686, B1 => n68073, B2 => 
                           n67935, ZN => n6852);
   U47288 : OAI22_X1 port map( A1 => n67943, A2 => n62685, B1 => n68076, B2 => 
                           n67935, ZN => n6853);
   U47289 : OAI22_X1 port map( A1 => n67943, A2 => n62684, B1 => n68079, B2 => 
                           n67935, ZN => n6854);
   U47290 : OAI22_X1 port map( A1 => n67943, A2 => n62683, B1 => n68082, B2 => 
                           n67935, ZN => n6855);
   U47291 : OAI22_X1 port map( A1 => n67943, A2 => n62682, B1 => n68085, B2 => 
                           n67935, ZN => n6856);
   U47292 : OAI22_X1 port map( A1 => n67943, A2 => n62681, B1 => n68088, B2 => 
                           n67935, ZN => n6857);
   U47293 : OAI22_X1 port map( A1 => n67943, A2 => n62680, B1 => n68091, B2 => 
                           n67935, ZN => n6858);
   U47294 : OAI22_X1 port map( A1 => n67944, A2 => n62679, B1 => n68094, B2 => 
                           n67936, ZN => n6859);
   U47295 : OAI22_X1 port map( A1 => n67944, A2 => n62678, B1 => n68097, B2 => 
                           n67936, ZN => n6860);
   U47296 : OAI22_X1 port map( A1 => n67944, A2 => n62677, B1 => n68100, B2 => 
                           n67936, ZN => n6861);
   U47297 : OAI22_X1 port map( A1 => n67944, A2 => n62676, B1 => n68103, B2 => 
                           n67936, ZN => n6862);
   U47298 : OAI22_X1 port map( A1 => n67944, A2 => n62675, B1 => n68106, B2 => 
                           n67936, ZN => n6863);
   U47299 : OAI22_X1 port map( A1 => n67944, A2 => n62674, B1 => n68109, B2 => 
                           n67936, ZN => n6864);
   U47300 : OAI22_X1 port map( A1 => n67944, A2 => n62673, B1 => n68112, B2 => 
                           n67936, ZN => n6865);
   U47301 : OAI22_X1 port map( A1 => n67944, A2 => n62672, B1 => n68115, B2 => 
                           n67936, ZN => n6866);
   U47302 : OAI22_X1 port map( A1 => n67944, A2 => n62671, B1 => n68118, B2 => 
                           n67936, ZN => n6867);
   U47303 : OAI22_X1 port map( A1 => n67944, A2 => n62670, B1 => n68121, B2 => 
                           n67936, ZN => n6868);
   U47304 : OAI22_X1 port map( A1 => n67944, A2 => n62669, B1 => n68124, B2 => 
                           n67936, ZN => n6869);
   U47305 : OAI22_X1 port map( A1 => n67944, A2 => n62668, B1 => n68127, B2 => 
                           n67936, ZN => n6870);
   U47306 : OAI22_X1 port map( A1 => n67944, A2 => n62667, B1 => n68130, B2 => 
                           n67937, ZN => n6871);
   U47307 : OAI22_X1 port map( A1 => n67945, A2 => n62666, B1 => n68133, B2 => 
                           n67937, ZN => n6872);
   U47308 : OAI22_X1 port map( A1 => n67945, A2 => n62665, B1 => n68136, B2 => 
                           n67937, ZN => n6873);
   U47309 : OAI22_X1 port map( A1 => n67945, A2 => n62664, B1 => n68139, B2 => 
                           n67937, ZN => n6874);
   U47310 : OAI22_X1 port map( A1 => n67945, A2 => n62663, B1 => n68142, B2 => 
                           n67937, ZN => n6875);
   U47311 : OAI22_X1 port map( A1 => n67945, A2 => n62662, B1 => n68145, B2 => 
                           n67937, ZN => n6876);
   U47312 : OAI22_X1 port map( A1 => n67945, A2 => n62661, B1 => n68148, B2 => 
                           n67937, ZN => n6877);
   U47313 : OAI22_X1 port map( A1 => n67945, A2 => n62660, B1 => n68151, B2 => 
                           n67937, ZN => n6878);
   U47314 : OAI22_X1 port map( A1 => n67945, A2 => n62659, B1 => n68154, B2 => 
                           n67937, ZN => n6879);
   U47315 : OAI22_X1 port map( A1 => n67945, A2 => n62658, B1 => n68157, B2 => 
                           n67937, ZN => n6880);
   U47316 : OAI22_X1 port map( A1 => n67945, A2 => n62657, B1 => n68160, B2 => 
                           n67937, ZN => n6881);
   U47317 : OAI22_X1 port map( A1 => n67945, A2 => n62656, B1 => n68163, B2 => 
                           n67937, ZN => n6882);
   U47318 : OAI22_X1 port map( A1 => n67945, A2 => n62655, B1 => n68166, B2 => 
                           n67938, ZN => n6883);
   U47319 : OAI22_X1 port map( A1 => n67945, A2 => n62654, B1 => n68169, B2 => 
                           n67938, ZN => n6884);
   U47320 : OAI22_X1 port map( A1 => n67946, A2 => n62653, B1 => n68172, B2 => 
                           n67938, ZN => n6885);
   U47321 : OAI22_X1 port map( A1 => n67946, A2 => n62652, B1 => n68175, B2 => 
                           n67938, ZN => n6886);
   U47322 : OAI22_X1 port map( A1 => n67946, A2 => n62651, B1 => n68178, B2 => 
                           n67938, ZN => n6887);
   U47323 : OAI22_X1 port map( A1 => n67946, A2 => n62650, B1 => n68181, B2 => 
                           n67938, ZN => n6888);
   U47324 : OAI22_X1 port map( A1 => n67946, A2 => n62649, B1 => n68184, B2 => 
                           n67938, ZN => n6889);
   U47325 : OAI22_X1 port map( A1 => n67946, A2 => n62648, B1 => n68187, B2 => 
                           n67938, ZN => n6890);
   U47326 : OAI22_X1 port map( A1 => n67946, A2 => n62647, B1 => n68190, B2 => 
                           n67938, ZN => n6891);
   U47327 : OAI22_X1 port map( A1 => n67946, A2 => n62646, B1 => n68193, B2 => 
                           n67938, ZN => n6892);
   U47328 : OAI22_X1 port map( A1 => n67946, A2 => n62645, B1 => n68196, B2 => 
                           n67938, ZN => n6893);
   U47329 : OAI22_X1 port map( A1 => n67946, A2 => n62644, B1 => n68199, B2 => 
                           n67938, ZN => n6894);
   U47330 : OAI22_X1 port map( A1 => n67946, A2 => n62643, B1 => n68202, B2 => 
                           n67939, ZN => n6895);
   U47331 : OAI22_X1 port map( A1 => n67946, A2 => n62642, B1 => n68205, B2 => 
                           n67939, ZN => n6896);
   U47332 : OAI22_X1 port map( A1 => n67946, A2 => n62641, B1 => n68208, B2 => 
                           n67939, ZN => n6897);
   U47333 : OAI22_X1 port map( A1 => n67947, A2 => n62640, B1 => n68211, B2 => 
                           n67939, ZN => n6898);
   U47334 : OAI22_X1 port map( A1 => n67947, A2 => n62639, B1 => n68214, B2 => 
                           n67939, ZN => n6899);
   U47335 : OAI22_X1 port map( A1 => n67947, A2 => n62638, B1 => n68217, B2 => 
                           n67939, ZN => n6900);
   U47336 : OAI22_X1 port map( A1 => n67947, A2 => n62637, B1 => n68220, B2 => 
                           n67939, ZN => n6901);
   U47337 : OAI22_X1 port map( A1 => n67947, A2 => n62636, B1 => n68223, B2 => 
                           n67939, ZN => n6902);
   U47338 : OAI22_X1 port map( A1 => n67947, A2 => n62635, B1 => n68226, B2 => 
                           n67939, ZN => n6903);
   U47339 : OAI22_X1 port map( A1 => n67947, A2 => n62634, B1 => n68229, B2 => 
                           n67939, ZN => n6904);
   U47340 : OAI22_X1 port map( A1 => n67947, A2 => n62633, B1 => n68232, B2 => 
                           n67939, ZN => n6905);
   U47341 : OAI22_X1 port map( A1 => n67947, A2 => n62632, B1 => n68235, B2 => 
                           n67939, ZN => n6906);
   U47342 : OAI22_X1 port map( A1 => n67956, A2 => n62624, B1 => n68058, B2 => 
                           n67948, ZN => n6911);
   U47343 : OAI22_X1 port map( A1 => n67956, A2 => n62623, B1 => n68061, B2 => 
                           n67948, ZN => n6912);
   U47344 : OAI22_X1 port map( A1 => n67956, A2 => n62622, B1 => n68064, B2 => 
                           n67948, ZN => n6913);
   U47345 : OAI22_X1 port map( A1 => n67956, A2 => n62621, B1 => n68067, B2 => 
                           n67948, ZN => n6914);
   U47346 : OAI22_X1 port map( A1 => n67956, A2 => n62620, B1 => n68070, B2 => 
                           n67948, ZN => n6915);
   U47347 : OAI22_X1 port map( A1 => n67956, A2 => n62619, B1 => n68073, B2 => 
                           n67948, ZN => n6916);
   U47348 : OAI22_X1 port map( A1 => n67956, A2 => n62618, B1 => n68076, B2 => 
                           n67948, ZN => n6917);
   U47349 : OAI22_X1 port map( A1 => n67956, A2 => n62617, B1 => n68079, B2 => 
                           n67948, ZN => n6918);
   U47350 : OAI22_X1 port map( A1 => n67956, A2 => n62616, B1 => n68082, B2 => 
                           n67948, ZN => n6919);
   U47351 : OAI22_X1 port map( A1 => n67956, A2 => n62615, B1 => n68085, B2 => 
                           n67948, ZN => n6920);
   U47352 : OAI22_X1 port map( A1 => n67956, A2 => n62614, B1 => n68088, B2 => 
                           n67948, ZN => n6921);
   U47353 : OAI22_X1 port map( A1 => n67956, A2 => n62613, B1 => n68091, B2 => 
                           n67948, ZN => n6922);
   U47354 : OAI22_X1 port map( A1 => n67957, A2 => n62612, B1 => n68094, B2 => 
                           n67949, ZN => n6923);
   U47355 : OAI22_X1 port map( A1 => n67957, A2 => n62611, B1 => n68097, B2 => 
                           n67949, ZN => n6924);
   U47356 : OAI22_X1 port map( A1 => n67957, A2 => n62610, B1 => n68100, B2 => 
                           n67949, ZN => n6925);
   U47357 : OAI22_X1 port map( A1 => n67957, A2 => n62609, B1 => n68103, B2 => 
                           n67949, ZN => n6926);
   U47358 : OAI22_X1 port map( A1 => n67957, A2 => n62608, B1 => n68106, B2 => 
                           n67949, ZN => n6927);
   U47359 : OAI22_X1 port map( A1 => n67957, A2 => n62607, B1 => n68109, B2 => 
                           n67949, ZN => n6928);
   U47360 : OAI22_X1 port map( A1 => n67957, A2 => n62606, B1 => n68112, B2 => 
                           n67949, ZN => n6929);
   U47361 : OAI22_X1 port map( A1 => n67957, A2 => n62605, B1 => n68115, B2 => 
                           n67949, ZN => n6930);
   U47362 : OAI22_X1 port map( A1 => n67957, A2 => n62604, B1 => n68118, B2 => 
                           n67949, ZN => n6931);
   U47363 : OAI22_X1 port map( A1 => n67957, A2 => n62603, B1 => n68121, B2 => 
                           n67949, ZN => n6932);
   U47364 : OAI22_X1 port map( A1 => n67957, A2 => n62602, B1 => n68124, B2 => 
                           n67949, ZN => n6933);
   U47365 : OAI22_X1 port map( A1 => n67957, A2 => n62601, B1 => n68127, B2 => 
                           n67949, ZN => n6934);
   U47366 : OAI22_X1 port map( A1 => n67957, A2 => n62600, B1 => n68130, B2 => 
                           n67950, ZN => n6935);
   U47367 : OAI22_X1 port map( A1 => n67958, A2 => n62599, B1 => n68133, B2 => 
                           n67950, ZN => n6936);
   U47368 : OAI22_X1 port map( A1 => n67958, A2 => n62598, B1 => n68136, B2 => 
                           n67950, ZN => n6937);
   U47369 : OAI22_X1 port map( A1 => n67958, A2 => n62597, B1 => n68139, B2 => 
                           n67950, ZN => n6938);
   U47370 : OAI22_X1 port map( A1 => n67958, A2 => n62596, B1 => n68142, B2 => 
                           n67950, ZN => n6939);
   U47371 : OAI22_X1 port map( A1 => n67958, A2 => n62595, B1 => n68145, B2 => 
                           n67950, ZN => n6940);
   U47372 : OAI22_X1 port map( A1 => n67958, A2 => n62594, B1 => n68148, B2 => 
                           n67950, ZN => n6941);
   U47373 : OAI22_X1 port map( A1 => n67958, A2 => n62593, B1 => n68151, B2 => 
                           n67950, ZN => n6942);
   U47374 : OAI22_X1 port map( A1 => n67958, A2 => n62592, B1 => n68154, B2 => 
                           n67950, ZN => n6943);
   U47375 : OAI22_X1 port map( A1 => n67958, A2 => n62591, B1 => n68157, B2 => 
                           n67950, ZN => n6944);
   U47376 : OAI22_X1 port map( A1 => n67958, A2 => n62590, B1 => n68160, B2 => 
                           n67950, ZN => n6945);
   U47377 : OAI22_X1 port map( A1 => n67958, A2 => n62589, B1 => n68163, B2 => 
                           n67950, ZN => n6946);
   U47378 : OAI22_X1 port map( A1 => n67958, A2 => n62588, B1 => n68166, B2 => 
                           n67951, ZN => n6947);
   U47379 : OAI22_X1 port map( A1 => n67958, A2 => n62587, B1 => n68169, B2 => 
                           n67951, ZN => n6948);
   U47380 : OAI22_X1 port map( A1 => n67959, A2 => n62586, B1 => n68172, B2 => 
                           n67951, ZN => n6949);
   U47381 : OAI22_X1 port map( A1 => n67959, A2 => n62585, B1 => n68175, B2 => 
                           n67951, ZN => n6950);
   U47382 : OAI22_X1 port map( A1 => n67959, A2 => n62584, B1 => n68178, B2 => 
                           n67951, ZN => n6951);
   U47383 : OAI22_X1 port map( A1 => n67959, A2 => n62583, B1 => n68181, B2 => 
                           n67951, ZN => n6952);
   U47384 : OAI22_X1 port map( A1 => n67959, A2 => n62582, B1 => n68184, B2 => 
                           n67951, ZN => n6953);
   U47385 : OAI22_X1 port map( A1 => n67959, A2 => n62581, B1 => n68187, B2 => 
                           n67951, ZN => n6954);
   U47386 : OAI22_X1 port map( A1 => n67959, A2 => n62580, B1 => n68190, B2 => 
                           n67951, ZN => n6955);
   U47387 : OAI22_X1 port map( A1 => n67959, A2 => n62579, B1 => n68193, B2 => 
                           n67951, ZN => n6956);
   U47388 : OAI22_X1 port map( A1 => n67959, A2 => n62578, B1 => n68196, B2 => 
                           n67951, ZN => n6957);
   U47389 : OAI22_X1 port map( A1 => n67959, A2 => n62577, B1 => n68199, B2 => 
                           n67951, ZN => n6958);
   U47390 : OAI22_X1 port map( A1 => n67959, A2 => n62576, B1 => n68202, B2 => 
                           n67952, ZN => n6959);
   U47391 : OAI22_X1 port map( A1 => n67959, A2 => n62575, B1 => n68205, B2 => 
                           n67952, ZN => n6960);
   U47392 : OAI22_X1 port map( A1 => n67959, A2 => n62574, B1 => n68208, B2 => 
                           n67952, ZN => n6961);
   U47393 : OAI22_X1 port map( A1 => n67960, A2 => n62573, B1 => n68211, B2 => 
                           n67952, ZN => n6962);
   U47394 : OAI22_X1 port map( A1 => n67960, A2 => n62572, B1 => n68214, B2 => 
                           n67952, ZN => n6963);
   U47395 : OAI22_X1 port map( A1 => n67960, A2 => n62571, B1 => n68217, B2 => 
                           n67952, ZN => n6964);
   U47396 : OAI22_X1 port map( A1 => n67960, A2 => n62570, B1 => n68220, B2 => 
                           n67952, ZN => n6965);
   U47397 : OAI22_X1 port map( A1 => n67960, A2 => n62569, B1 => n68223, B2 => 
                           n67952, ZN => n6966);
   U47398 : OAI22_X1 port map( A1 => n67960, A2 => n62568, B1 => n68226, B2 => 
                           n67952, ZN => n6967);
   U47399 : OAI22_X1 port map( A1 => n67960, A2 => n62567, B1 => n68229, B2 => 
                           n67952, ZN => n6968);
   U47400 : OAI22_X1 port map( A1 => n67960, A2 => n62566, B1 => n68232, B2 => 
                           n67952, ZN => n6969);
   U47401 : OAI22_X1 port map( A1 => n67960, A2 => n62565, B1 => n68235, B2 => 
                           n67952, ZN => n6970);
   U47402 : OAI22_X1 port map( A1 => n68047, A2 => n62155, B1 => n68058, B2 => 
                           n68039, ZN => n7359);
   U47403 : OAI22_X1 port map( A1 => n68047, A2 => n62154, B1 => n68061, B2 => 
                           n68039, ZN => n7360);
   U47404 : OAI22_X1 port map( A1 => n68047, A2 => n62153, B1 => n68064, B2 => 
                           n68039, ZN => n7361);
   U47405 : OAI22_X1 port map( A1 => n68047, A2 => n62152, B1 => n68067, B2 => 
                           n68039, ZN => n7362);
   U47406 : OAI22_X1 port map( A1 => n68047, A2 => n62151, B1 => n68070, B2 => 
                           n68039, ZN => n7363);
   U47407 : OAI22_X1 port map( A1 => n68047, A2 => n62150, B1 => n68073, B2 => 
                           n68039, ZN => n7364);
   U47408 : OAI22_X1 port map( A1 => n68047, A2 => n62149, B1 => n68076, B2 => 
                           n68039, ZN => n7365);
   U47409 : OAI22_X1 port map( A1 => n68047, A2 => n62148, B1 => n68079, B2 => 
                           n68039, ZN => n7366);
   U47410 : OAI22_X1 port map( A1 => n68047, A2 => n62147, B1 => n68082, B2 => 
                           n68039, ZN => n7367);
   U47411 : OAI22_X1 port map( A1 => n68047, A2 => n62146, B1 => n68085, B2 => 
                           n68039, ZN => n7368);
   U47412 : OAI22_X1 port map( A1 => n68047, A2 => n62145, B1 => n68088, B2 => 
                           n68039, ZN => n7369);
   U47413 : OAI22_X1 port map( A1 => n68047, A2 => n62144, B1 => n68091, B2 => 
                           n68039, ZN => n7370);
   U47414 : OAI22_X1 port map( A1 => n68048, A2 => n62143, B1 => n68094, B2 => 
                           n68040, ZN => n7371);
   U47415 : OAI22_X1 port map( A1 => n68048, A2 => n62142, B1 => n68097, B2 => 
                           n68040, ZN => n7372);
   U47416 : OAI22_X1 port map( A1 => n68048, A2 => n62141, B1 => n68100, B2 => 
                           n68040, ZN => n7373);
   U47417 : OAI22_X1 port map( A1 => n68048, A2 => n62140, B1 => n68103, B2 => 
                           n68040, ZN => n7374);
   U47418 : OAI22_X1 port map( A1 => n68048, A2 => n62139, B1 => n68106, B2 => 
                           n68040, ZN => n7375);
   U47419 : OAI22_X1 port map( A1 => n68048, A2 => n62138, B1 => n68109, B2 => 
                           n68040, ZN => n7376);
   U47420 : OAI22_X1 port map( A1 => n68048, A2 => n62137, B1 => n68112, B2 => 
                           n68040, ZN => n7377);
   U47421 : OAI22_X1 port map( A1 => n68048, A2 => n62136, B1 => n68115, B2 => 
                           n68040, ZN => n7378);
   U47422 : OAI22_X1 port map( A1 => n68048, A2 => n62135, B1 => n68118, B2 => 
                           n68040, ZN => n7379);
   U47423 : OAI22_X1 port map( A1 => n68048, A2 => n62134, B1 => n68121, B2 => 
                           n68040, ZN => n7380);
   U47424 : OAI22_X1 port map( A1 => n68048, A2 => n62133, B1 => n68124, B2 => 
                           n68040, ZN => n7381);
   U47425 : OAI22_X1 port map( A1 => n68048, A2 => n62132, B1 => n68127, B2 => 
                           n68040, ZN => n7382);
   U47426 : OAI22_X1 port map( A1 => n68048, A2 => n62131, B1 => n68130, B2 => 
                           n68041, ZN => n7383);
   U47427 : OAI22_X1 port map( A1 => n68049, A2 => n62130, B1 => n68133, B2 => 
                           n68041, ZN => n7384);
   U47428 : OAI22_X1 port map( A1 => n68049, A2 => n62129, B1 => n68136, B2 => 
                           n68041, ZN => n7385);
   U47429 : OAI22_X1 port map( A1 => n68049, A2 => n62128, B1 => n68139, B2 => 
                           n68041, ZN => n7386);
   U47430 : OAI22_X1 port map( A1 => n68049, A2 => n62127, B1 => n68142, B2 => 
                           n68041, ZN => n7387);
   U47431 : OAI22_X1 port map( A1 => n68049, A2 => n62126, B1 => n68145, B2 => 
                           n68041, ZN => n7388);
   U47432 : OAI22_X1 port map( A1 => n68049, A2 => n62125, B1 => n68148, B2 => 
                           n68041, ZN => n7389);
   U47433 : OAI22_X1 port map( A1 => n68049, A2 => n62124, B1 => n68151, B2 => 
                           n68041, ZN => n7390);
   U47434 : OAI22_X1 port map( A1 => n68049, A2 => n62123, B1 => n68154, B2 => 
                           n68041, ZN => n7391);
   U47435 : OAI22_X1 port map( A1 => n68049, A2 => n62122, B1 => n68157, B2 => 
                           n68041, ZN => n7392);
   U47436 : OAI22_X1 port map( A1 => n68049, A2 => n62121, B1 => n68160, B2 => 
                           n68041, ZN => n7393);
   U47437 : OAI22_X1 port map( A1 => n68049, A2 => n62120, B1 => n68163, B2 => 
                           n68041, ZN => n7394);
   U47438 : OAI22_X1 port map( A1 => n68049, A2 => n62119, B1 => n68166, B2 => 
                           n68042, ZN => n7395);
   U47439 : OAI22_X1 port map( A1 => n68049, A2 => n62118, B1 => n68169, B2 => 
                           n68042, ZN => n7396);
   U47440 : OAI22_X1 port map( A1 => n68050, A2 => n62117, B1 => n68172, B2 => 
                           n68042, ZN => n7397);
   U47441 : OAI22_X1 port map( A1 => n68050, A2 => n62116, B1 => n68175, B2 => 
                           n68042, ZN => n7398);
   U47442 : OAI22_X1 port map( A1 => n68050, A2 => n62115, B1 => n68178, B2 => 
                           n68042, ZN => n7399);
   U47443 : OAI22_X1 port map( A1 => n68050, A2 => n62114, B1 => n68181, B2 => 
                           n68042, ZN => n7400);
   U47444 : OAI22_X1 port map( A1 => n68050, A2 => n62113, B1 => n68184, B2 => 
                           n68042, ZN => n7401);
   U47445 : OAI22_X1 port map( A1 => n68050, A2 => n62112, B1 => n68187, B2 => 
                           n68042, ZN => n7402);
   U47446 : OAI22_X1 port map( A1 => n68050, A2 => n62111, B1 => n68190, B2 => 
                           n68042, ZN => n7403);
   U47447 : OAI22_X1 port map( A1 => n68050, A2 => n62110, B1 => n68193, B2 => 
                           n68042, ZN => n7404);
   U47448 : OAI22_X1 port map( A1 => n68050, A2 => n62109, B1 => n68196, B2 => 
                           n68042, ZN => n7405);
   U47449 : OAI22_X1 port map( A1 => n68050, A2 => n62108, B1 => n68199, B2 => 
                           n68042, ZN => n7406);
   U47450 : OAI22_X1 port map( A1 => n68050, A2 => n62107, B1 => n68202, B2 => 
                           n68043, ZN => n7407);
   U47451 : OAI22_X1 port map( A1 => n68050, A2 => n62106, B1 => n68205, B2 => 
                           n68043, ZN => n7408);
   U47452 : OAI22_X1 port map( A1 => n68050, A2 => n62105, B1 => n68208, B2 => 
                           n68043, ZN => n7409);
   U47453 : OAI22_X1 port map( A1 => n68051, A2 => n62104, B1 => n68211, B2 => 
                           n68043, ZN => n7410);
   U47454 : OAI22_X1 port map( A1 => n68051, A2 => n62103, B1 => n68214, B2 => 
                           n68043, ZN => n7411);
   U47455 : OAI22_X1 port map( A1 => n68051, A2 => n62102, B1 => n68217, B2 => 
                           n68043, ZN => n7412);
   U47456 : OAI22_X1 port map( A1 => n68051, A2 => n62101, B1 => n68220, B2 => 
                           n68043, ZN => n7413);
   U47457 : OAI22_X1 port map( A1 => n68051, A2 => n62100, B1 => n68223, B2 => 
                           n68043, ZN => n7414);
   U47458 : OAI22_X1 port map( A1 => n68051, A2 => n62099, B1 => n68226, B2 => 
                           n68043, ZN => n7415);
   U47459 : OAI22_X1 port map( A1 => n68051, A2 => n62098, B1 => n68229, B2 => 
                           n68043, ZN => n7416);
   U47460 : OAI22_X1 port map( A1 => n68051, A2 => n62097, B1 => n68232, B2 => 
                           n68043, ZN => n7417);
   U47461 : OAI22_X1 port map( A1 => n68051, A2 => n62096, B1 => n68235, B2 => 
                           n68043, ZN => n7418);
   U47462 : OAI22_X1 port map( A1 => n68008, A2 => n62355, B1 => n68058, B2 => 
                           n68000, ZN => n7167);
   U47463 : OAI22_X1 port map( A1 => n68008, A2 => n62354, B1 => n68061, B2 => 
                           n68000, ZN => n7168);
   U47464 : OAI22_X1 port map( A1 => n68008, A2 => n62353, B1 => n68064, B2 => 
                           n68000, ZN => n7169);
   U47465 : OAI22_X1 port map( A1 => n68008, A2 => n62352, B1 => n68067, B2 => 
                           n68000, ZN => n7170);
   U47466 : OAI22_X1 port map( A1 => n68008, A2 => n62351, B1 => n68070, B2 => 
                           n68000, ZN => n7171);
   U47467 : OAI22_X1 port map( A1 => n68008, A2 => n62350, B1 => n68073, B2 => 
                           n68000, ZN => n7172);
   U47468 : OAI22_X1 port map( A1 => n68008, A2 => n62349, B1 => n68076, B2 => 
                           n68000, ZN => n7173);
   U47469 : OAI22_X1 port map( A1 => n68008, A2 => n62348, B1 => n68079, B2 => 
                           n68000, ZN => n7174);
   U47470 : OAI22_X1 port map( A1 => n68008, A2 => n62347, B1 => n68082, B2 => 
                           n68000, ZN => n7175);
   U47471 : OAI22_X1 port map( A1 => n68008, A2 => n62346, B1 => n68085, B2 => 
                           n68000, ZN => n7176);
   U47472 : OAI22_X1 port map( A1 => n68008, A2 => n62345, B1 => n68088, B2 => 
                           n68000, ZN => n7177);
   U47473 : OAI22_X1 port map( A1 => n68008, A2 => n62344, B1 => n68091, B2 => 
                           n68000, ZN => n7178);
   U47474 : OAI22_X1 port map( A1 => n68009, A2 => n62343, B1 => n68094, B2 => 
                           n68001, ZN => n7179);
   U47475 : OAI22_X1 port map( A1 => n68009, A2 => n62342, B1 => n68097, B2 => 
                           n68001, ZN => n7180);
   U47476 : OAI22_X1 port map( A1 => n68009, A2 => n62341, B1 => n68100, B2 => 
                           n68001, ZN => n7181);
   U47477 : OAI22_X1 port map( A1 => n68009, A2 => n62340, B1 => n68103, B2 => 
                           n68001, ZN => n7182);
   U47478 : OAI22_X1 port map( A1 => n68009, A2 => n62339, B1 => n68106, B2 => 
                           n68001, ZN => n7183);
   U47479 : OAI22_X1 port map( A1 => n68009, A2 => n62338, B1 => n68109, B2 => 
                           n68001, ZN => n7184);
   U47480 : OAI22_X1 port map( A1 => n68009, A2 => n62337, B1 => n68112, B2 => 
                           n68001, ZN => n7185);
   U47481 : OAI22_X1 port map( A1 => n68009, A2 => n62336, B1 => n68115, B2 => 
                           n68001, ZN => n7186);
   U47482 : OAI22_X1 port map( A1 => n68009, A2 => n62335, B1 => n68118, B2 => 
                           n68001, ZN => n7187);
   U47483 : OAI22_X1 port map( A1 => n68009, A2 => n62334, B1 => n68121, B2 => 
                           n68001, ZN => n7188);
   U47484 : OAI22_X1 port map( A1 => n68009, A2 => n62333, B1 => n68124, B2 => 
                           n68001, ZN => n7189);
   U47485 : OAI22_X1 port map( A1 => n68009, A2 => n62332, B1 => n68127, B2 => 
                           n68001, ZN => n7190);
   U47486 : OAI22_X1 port map( A1 => n68009, A2 => n62331, B1 => n68130, B2 => 
                           n68002, ZN => n7191);
   U47487 : OAI22_X1 port map( A1 => n68010, A2 => n62330, B1 => n68133, B2 => 
                           n68002, ZN => n7192);
   U47488 : OAI22_X1 port map( A1 => n68010, A2 => n62329, B1 => n68136, B2 => 
                           n68002, ZN => n7193);
   U47489 : OAI22_X1 port map( A1 => n68010, A2 => n62328, B1 => n68139, B2 => 
                           n68002, ZN => n7194);
   U47490 : OAI22_X1 port map( A1 => n68010, A2 => n62327, B1 => n68142, B2 => 
                           n68002, ZN => n7195);
   U47491 : OAI22_X1 port map( A1 => n68010, A2 => n62326, B1 => n68145, B2 => 
                           n68002, ZN => n7196);
   U47492 : OAI22_X1 port map( A1 => n68010, A2 => n62325, B1 => n68148, B2 => 
                           n68002, ZN => n7197);
   U47493 : OAI22_X1 port map( A1 => n68010, A2 => n62324, B1 => n68151, B2 => 
                           n68002, ZN => n7198);
   U47494 : OAI22_X1 port map( A1 => n68010, A2 => n62323, B1 => n68154, B2 => 
                           n68002, ZN => n7199);
   U47495 : OAI22_X1 port map( A1 => n68010, A2 => n62322, B1 => n68157, B2 => 
                           n68002, ZN => n7200);
   U47496 : OAI22_X1 port map( A1 => n68010, A2 => n62321, B1 => n68160, B2 => 
                           n68002, ZN => n7201);
   U47497 : OAI22_X1 port map( A1 => n68010, A2 => n62320, B1 => n68163, B2 => 
                           n68002, ZN => n7202);
   U47498 : OAI22_X1 port map( A1 => n68010, A2 => n62319, B1 => n68166, B2 => 
                           n68003, ZN => n7203);
   U47499 : OAI22_X1 port map( A1 => n68010, A2 => n62318, B1 => n68169, B2 => 
                           n68003, ZN => n7204);
   U47500 : OAI22_X1 port map( A1 => n68011, A2 => n62317, B1 => n68172, B2 => 
                           n68003, ZN => n7205);
   U47501 : OAI22_X1 port map( A1 => n68011, A2 => n62316, B1 => n68175, B2 => 
                           n68003, ZN => n7206);
   U47502 : OAI22_X1 port map( A1 => n68011, A2 => n62315, B1 => n68178, B2 => 
                           n68003, ZN => n7207);
   U47503 : OAI22_X1 port map( A1 => n68011, A2 => n62314, B1 => n68181, B2 => 
                           n68003, ZN => n7208);
   U47504 : OAI22_X1 port map( A1 => n68011, A2 => n62313, B1 => n68184, B2 => 
                           n68003, ZN => n7209);
   U47505 : OAI22_X1 port map( A1 => n68011, A2 => n62312, B1 => n68187, B2 => 
                           n68003, ZN => n7210);
   U47506 : OAI22_X1 port map( A1 => n68011, A2 => n62311, B1 => n68190, B2 => 
                           n68003, ZN => n7211);
   U47507 : OAI22_X1 port map( A1 => n68011, A2 => n62310, B1 => n68193, B2 => 
                           n68003, ZN => n7212);
   U47508 : OAI22_X1 port map( A1 => n68011, A2 => n62309, B1 => n68196, B2 => 
                           n68003, ZN => n7213);
   U47509 : OAI22_X1 port map( A1 => n68011, A2 => n62308, B1 => n68199, B2 => 
                           n68003, ZN => n7214);
   U47510 : OAI22_X1 port map( A1 => n68011, A2 => n62307, B1 => n68202, B2 => 
                           n68004, ZN => n7215);
   U47511 : OAI22_X1 port map( A1 => n68011, A2 => n62306, B1 => n68205, B2 => 
                           n68004, ZN => n7216);
   U47512 : OAI22_X1 port map( A1 => n68011, A2 => n62305, B1 => n68208, B2 => 
                           n68004, ZN => n7217);
   U47513 : OAI22_X1 port map( A1 => n68012, A2 => n62304, B1 => n68211, B2 => 
                           n68004, ZN => n7218);
   U47514 : OAI22_X1 port map( A1 => n68012, A2 => n62303, B1 => n68214, B2 => 
                           n68004, ZN => n7219);
   U47515 : OAI22_X1 port map( A1 => n68012, A2 => n62302, B1 => n68217, B2 => 
                           n68004, ZN => n7220);
   U47516 : OAI22_X1 port map( A1 => n68012, A2 => n62301, B1 => n68220, B2 => 
                           n68004, ZN => n7221);
   U47517 : OAI22_X1 port map( A1 => n68012, A2 => n62300, B1 => n68223, B2 => 
                           n68004, ZN => n7222);
   U47518 : OAI22_X1 port map( A1 => n68012, A2 => n62299, B1 => n68226, B2 => 
                           n68004, ZN => n7223);
   U47519 : OAI22_X1 port map( A1 => n68012, A2 => n62298, B1 => n68229, B2 => 
                           n68004, ZN => n7224);
   U47520 : OAI22_X1 port map( A1 => n68012, A2 => n62297, B1 => n68232, B2 => 
                           n68004, ZN => n7225);
   U47521 : OAI22_X1 port map( A1 => n68012, A2 => n62296, B1 => n68235, B2 => 
                           n68004, ZN => n7226);
   U47522 : OAI22_X1 port map( A1 => n67969, A2 => n62558, B1 => n68058, B2 => 
                           n67961, ZN => n6975);
   U47523 : OAI22_X1 port map( A1 => n67969, A2 => n62557, B1 => n68061, B2 => 
                           n67961, ZN => n6976);
   U47524 : OAI22_X1 port map( A1 => n67969, A2 => n62556, B1 => n68064, B2 => 
                           n67961, ZN => n6977);
   U47525 : OAI22_X1 port map( A1 => n67969, A2 => n62555, B1 => n68067, B2 => 
                           n67961, ZN => n6978);
   U47526 : OAI22_X1 port map( A1 => n67969, A2 => n62554, B1 => n68070, B2 => 
                           n67961, ZN => n6979);
   U47527 : OAI22_X1 port map( A1 => n67969, A2 => n62553, B1 => n68073, B2 => 
                           n67961, ZN => n6980);
   U47528 : OAI22_X1 port map( A1 => n67969, A2 => n62552, B1 => n68076, B2 => 
                           n67961, ZN => n6981);
   U47529 : OAI22_X1 port map( A1 => n67969, A2 => n62551, B1 => n68079, B2 => 
                           n67961, ZN => n6982);
   U47530 : OAI22_X1 port map( A1 => n67969, A2 => n62550, B1 => n68082, B2 => 
                           n67961, ZN => n6983);
   U47531 : OAI22_X1 port map( A1 => n67969, A2 => n62549, B1 => n68085, B2 => 
                           n67961, ZN => n6984);
   U47532 : OAI22_X1 port map( A1 => n67969, A2 => n62548, B1 => n68088, B2 => 
                           n67961, ZN => n6985);
   U47533 : OAI22_X1 port map( A1 => n67969, A2 => n62547, B1 => n68091, B2 => 
                           n67961, ZN => n6986);
   U47534 : OAI22_X1 port map( A1 => n67970, A2 => n62546, B1 => n68094, B2 => 
                           n67962, ZN => n6987);
   U47535 : OAI22_X1 port map( A1 => n67970, A2 => n62545, B1 => n68097, B2 => 
                           n67962, ZN => n6988);
   U47536 : OAI22_X1 port map( A1 => n67970, A2 => n62544, B1 => n68100, B2 => 
                           n67962, ZN => n6989);
   U47537 : OAI22_X1 port map( A1 => n67970, A2 => n62543, B1 => n68103, B2 => 
                           n67962, ZN => n6990);
   U47538 : OAI22_X1 port map( A1 => n67970, A2 => n62542, B1 => n68106, B2 => 
                           n67962, ZN => n6991);
   U47539 : OAI22_X1 port map( A1 => n67970, A2 => n62541, B1 => n68109, B2 => 
                           n67962, ZN => n6992);
   U47540 : OAI22_X1 port map( A1 => n67970, A2 => n62540, B1 => n68112, B2 => 
                           n67962, ZN => n6993);
   U47541 : OAI22_X1 port map( A1 => n67970, A2 => n62539, B1 => n68115, B2 => 
                           n67962, ZN => n6994);
   U47542 : OAI22_X1 port map( A1 => n67970, A2 => n62538, B1 => n68118, B2 => 
                           n67962, ZN => n6995);
   U47543 : OAI22_X1 port map( A1 => n67970, A2 => n62537, B1 => n68121, B2 => 
                           n67962, ZN => n6996);
   U47544 : OAI22_X1 port map( A1 => n67970, A2 => n62536, B1 => n68124, B2 => 
                           n67962, ZN => n6997);
   U47545 : OAI22_X1 port map( A1 => n67970, A2 => n62535, B1 => n68127, B2 => 
                           n67962, ZN => n6998);
   U47546 : OAI22_X1 port map( A1 => n67970, A2 => n62534, B1 => n68130, B2 => 
                           n67963, ZN => n6999);
   U47547 : OAI22_X1 port map( A1 => n67971, A2 => n62533, B1 => n68133, B2 => 
                           n67963, ZN => n7000);
   U47548 : OAI22_X1 port map( A1 => n67971, A2 => n62532, B1 => n68136, B2 => 
                           n67963, ZN => n7001);
   U47549 : OAI22_X1 port map( A1 => n67971, A2 => n62531, B1 => n68139, B2 => 
                           n67963, ZN => n7002);
   U47550 : OAI22_X1 port map( A1 => n67971, A2 => n62530, B1 => n68142, B2 => 
                           n67963, ZN => n7003);
   U47551 : OAI22_X1 port map( A1 => n67971, A2 => n62529, B1 => n68145, B2 => 
                           n67963, ZN => n7004);
   U47552 : OAI22_X1 port map( A1 => n67971, A2 => n62528, B1 => n68148, B2 => 
                           n67963, ZN => n7005);
   U47553 : OAI22_X1 port map( A1 => n67971, A2 => n62527, B1 => n68151, B2 => 
                           n67963, ZN => n7006);
   U47554 : OAI22_X1 port map( A1 => n67971, A2 => n62526, B1 => n68154, B2 => 
                           n67963, ZN => n7007);
   U47555 : OAI22_X1 port map( A1 => n67971, A2 => n62525, B1 => n68157, B2 => 
                           n67963, ZN => n7008);
   U47556 : OAI22_X1 port map( A1 => n67971, A2 => n62524, B1 => n68160, B2 => 
                           n67963, ZN => n7009);
   U47557 : OAI22_X1 port map( A1 => n67971, A2 => n62523, B1 => n68163, B2 => 
                           n67963, ZN => n7010);
   U47558 : OAI22_X1 port map( A1 => n67971, A2 => n62522, B1 => n68166, B2 => 
                           n67964, ZN => n7011);
   U47559 : OAI22_X1 port map( A1 => n67971, A2 => n62521, B1 => n68169, B2 => 
                           n67964, ZN => n7012);
   U47560 : OAI22_X1 port map( A1 => n67972, A2 => n62520, B1 => n68172, B2 => 
                           n67964, ZN => n7013);
   U47561 : OAI22_X1 port map( A1 => n67972, A2 => n62519, B1 => n68175, B2 => 
                           n67964, ZN => n7014);
   U47562 : OAI22_X1 port map( A1 => n67972, A2 => n62518, B1 => n68178, B2 => 
                           n67964, ZN => n7015);
   U47563 : OAI22_X1 port map( A1 => n67972, A2 => n62517, B1 => n68181, B2 => 
                           n67964, ZN => n7016);
   U47564 : OAI22_X1 port map( A1 => n67972, A2 => n62516, B1 => n68184, B2 => 
                           n67964, ZN => n7017);
   U47565 : OAI22_X1 port map( A1 => n67972, A2 => n62515, B1 => n68187, B2 => 
                           n67964, ZN => n7018);
   U47566 : OAI22_X1 port map( A1 => n67972, A2 => n62514, B1 => n68190, B2 => 
                           n67964, ZN => n7019);
   U47567 : OAI22_X1 port map( A1 => n67972, A2 => n62513, B1 => n68193, B2 => 
                           n67964, ZN => n7020);
   U47568 : OAI22_X1 port map( A1 => n67972, A2 => n62512, B1 => n68196, B2 => 
                           n67964, ZN => n7021);
   U47569 : OAI22_X1 port map( A1 => n67972, A2 => n62511, B1 => n68199, B2 => 
                           n67964, ZN => n7022);
   U47570 : OAI22_X1 port map( A1 => n67972, A2 => n62510, B1 => n68202, B2 => 
                           n67965, ZN => n7023);
   U47571 : OAI22_X1 port map( A1 => n67972, A2 => n62509, B1 => n68205, B2 => 
                           n67965, ZN => n7024);
   U47572 : OAI22_X1 port map( A1 => n67972, A2 => n62508, B1 => n68208, B2 => 
                           n67965, ZN => n7025);
   U47573 : OAI22_X1 port map( A1 => n67973, A2 => n62507, B1 => n68211, B2 => 
                           n67965, ZN => n7026);
   U47574 : OAI22_X1 port map( A1 => n67973, A2 => n62506, B1 => n68214, B2 => 
                           n67965, ZN => n7027);
   U47575 : OAI22_X1 port map( A1 => n67973, A2 => n62505, B1 => n68217, B2 => 
                           n67965, ZN => n7028);
   U47576 : OAI22_X1 port map( A1 => n67973, A2 => n62504, B1 => n68220, B2 => 
                           n67965, ZN => n7029);
   U47577 : OAI22_X1 port map( A1 => n67973, A2 => n62503, B1 => n68223, B2 => 
                           n67965, ZN => n7030);
   U47578 : OAI22_X1 port map( A1 => n67973, A2 => n62502, B1 => n68226, B2 => 
                           n67965, ZN => n7031);
   U47579 : OAI22_X1 port map( A1 => n67973, A2 => n62501, B1 => n68229, B2 => 
                           n67965, ZN => n7032);
   U47580 : OAI22_X1 port map( A1 => n67973, A2 => n62500, B1 => n68232, B2 => 
                           n67965, ZN => n7033);
   U47581 : OAI22_X1 port map( A1 => n67973, A2 => n62499, B1 => n68235, B2 => 
                           n67965, ZN => n7034);
   U47582 : OAI22_X1 port map( A1 => n67803, A2 => n63226, B1 => n68059, B2 => 
                           n67795, ZN => n6143);
   U47583 : OAI22_X1 port map( A1 => n67803, A2 => n63225, B1 => n68062, B2 => 
                           n67795, ZN => n6144);
   U47584 : OAI22_X1 port map( A1 => n67803, A2 => n63224, B1 => n68065, B2 => 
                           n67795, ZN => n6145);
   U47585 : OAI22_X1 port map( A1 => n67803, A2 => n63223, B1 => n68068, B2 => 
                           n67795, ZN => n6146);
   U47586 : OAI22_X1 port map( A1 => n67803, A2 => n63222, B1 => n68071, B2 => 
                           n67795, ZN => n6147);
   U47587 : OAI22_X1 port map( A1 => n67803, A2 => n63221, B1 => n68074, B2 => 
                           n67795, ZN => n6148);
   U47588 : OAI22_X1 port map( A1 => n67803, A2 => n63220, B1 => n68077, B2 => 
                           n67795, ZN => n6149);
   U47589 : OAI22_X1 port map( A1 => n67803, A2 => n63219, B1 => n68080, B2 => 
                           n67795, ZN => n6150);
   U47590 : OAI22_X1 port map( A1 => n67803, A2 => n63218, B1 => n68083, B2 => 
                           n67795, ZN => n6151);
   U47591 : OAI22_X1 port map( A1 => n67803, A2 => n63217, B1 => n68086, B2 => 
                           n67795, ZN => n6152);
   U47592 : OAI22_X1 port map( A1 => n67803, A2 => n63216, B1 => n68089, B2 => 
                           n67795, ZN => n6153);
   U47593 : OAI22_X1 port map( A1 => n67803, A2 => n63215, B1 => n68092, B2 => 
                           n67795, ZN => n6154);
   U47594 : OAI22_X1 port map( A1 => n67804, A2 => n63214, B1 => n68095, B2 => 
                           n67796, ZN => n6155);
   U47595 : OAI22_X1 port map( A1 => n67804, A2 => n63213, B1 => n68098, B2 => 
                           n67796, ZN => n6156);
   U47596 : OAI22_X1 port map( A1 => n67804, A2 => n63212, B1 => n68101, B2 => 
                           n67796, ZN => n6157);
   U47597 : OAI22_X1 port map( A1 => n67804, A2 => n63211, B1 => n68104, B2 => 
                           n67796, ZN => n6158);
   U47598 : OAI22_X1 port map( A1 => n67804, A2 => n63210, B1 => n68107, B2 => 
                           n67796, ZN => n6159);
   U47599 : OAI22_X1 port map( A1 => n67804, A2 => n63209, B1 => n68110, B2 => 
                           n67796, ZN => n6160);
   U47600 : OAI22_X1 port map( A1 => n67804, A2 => n63208, B1 => n68113, B2 => 
                           n67796, ZN => n6161);
   U47601 : OAI22_X1 port map( A1 => n67804, A2 => n63207, B1 => n68116, B2 => 
                           n67796, ZN => n6162);
   U47602 : OAI22_X1 port map( A1 => n67804, A2 => n63206, B1 => n68119, B2 => 
                           n67796, ZN => n6163);
   U47603 : OAI22_X1 port map( A1 => n67804, A2 => n63205, B1 => n68122, B2 => 
                           n67796, ZN => n6164);
   U47604 : OAI22_X1 port map( A1 => n67804, A2 => n63204, B1 => n68125, B2 => 
                           n67796, ZN => n6165);
   U47605 : OAI22_X1 port map( A1 => n67804, A2 => n63203, B1 => n68128, B2 => 
                           n67796, ZN => n6166);
   U47606 : OAI22_X1 port map( A1 => n67804, A2 => n63202, B1 => n68131, B2 => 
                           n67797, ZN => n6167);
   U47607 : OAI22_X1 port map( A1 => n67805, A2 => n63201, B1 => n68134, B2 => 
                           n67797, ZN => n6168);
   U47608 : OAI22_X1 port map( A1 => n67805, A2 => n63200, B1 => n68137, B2 => 
                           n67797, ZN => n6169);
   U47609 : OAI22_X1 port map( A1 => n67805, A2 => n63199, B1 => n68140, B2 => 
                           n67797, ZN => n6170);
   U47610 : OAI22_X1 port map( A1 => n67805, A2 => n63198, B1 => n68143, B2 => 
                           n67797, ZN => n6171);
   U47611 : OAI22_X1 port map( A1 => n67805, A2 => n63197, B1 => n68146, B2 => 
                           n67797, ZN => n6172);
   U47612 : OAI22_X1 port map( A1 => n67805, A2 => n63196, B1 => n68149, B2 => 
                           n67797, ZN => n6173);
   U47613 : OAI22_X1 port map( A1 => n67805, A2 => n63195, B1 => n68152, B2 => 
                           n67797, ZN => n6174);
   U47614 : OAI22_X1 port map( A1 => n67805, A2 => n63194, B1 => n68155, B2 => 
                           n67797, ZN => n6175);
   U47615 : OAI22_X1 port map( A1 => n67805, A2 => n63193, B1 => n68158, B2 => 
                           n67797, ZN => n6176);
   U47616 : OAI22_X1 port map( A1 => n67805, A2 => n63192, B1 => n68161, B2 => 
                           n67797, ZN => n6177);
   U47617 : OAI22_X1 port map( A1 => n67805, A2 => n63191, B1 => n68164, B2 => 
                           n67797, ZN => n6178);
   U47618 : OAI22_X1 port map( A1 => n67805, A2 => n63190, B1 => n68167, B2 => 
                           n67798, ZN => n6179);
   U47619 : OAI22_X1 port map( A1 => n67805, A2 => n63189, B1 => n68170, B2 => 
                           n67798, ZN => n6180);
   U47620 : OAI22_X1 port map( A1 => n67806, A2 => n63188, B1 => n68173, B2 => 
                           n67798, ZN => n6181);
   U47621 : OAI22_X1 port map( A1 => n67806, A2 => n63187, B1 => n68176, B2 => 
                           n67798, ZN => n6182);
   U47622 : OAI22_X1 port map( A1 => n67806, A2 => n63186, B1 => n68179, B2 => 
                           n67798, ZN => n6183);
   U47623 : OAI22_X1 port map( A1 => n67806, A2 => n63185, B1 => n68182, B2 => 
                           n67798, ZN => n6184);
   U47624 : OAI22_X1 port map( A1 => n67806, A2 => n63184, B1 => n68185, B2 => 
                           n67798, ZN => n6185);
   U47625 : OAI22_X1 port map( A1 => n67806, A2 => n63183, B1 => n68188, B2 => 
                           n67798, ZN => n6186);
   U47626 : OAI22_X1 port map( A1 => n67806, A2 => n63182, B1 => n68191, B2 => 
                           n67798, ZN => n6187);
   U47627 : OAI22_X1 port map( A1 => n67806, A2 => n63181, B1 => n68194, B2 => 
                           n67798, ZN => n6188);
   U47628 : OAI22_X1 port map( A1 => n67806, A2 => n63180, B1 => n68197, B2 => 
                           n67798, ZN => n6189);
   U47629 : OAI22_X1 port map( A1 => n67806, A2 => n63179, B1 => n68200, B2 => 
                           n67798, ZN => n6190);
   U47630 : OAI22_X1 port map( A1 => n67806, A2 => n63178, B1 => n68203, B2 => 
                           n67799, ZN => n6191);
   U47631 : OAI22_X1 port map( A1 => n67806, A2 => n63177, B1 => n68206, B2 => 
                           n67799, ZN => n6192);
   U47632 : OAI22_X1 port map( A1 => n67806, A2 => n63176, B1 => n68209, B2 => 
                           n67799, ZN => n6193);
   U47633 : OAI22_X1 port map( A1 => n67807, A2 => n63175, B1 => n68212, B2 => 
                           n67799, ZN => n6194);
   U47634 : OAI22_X1 port map( A1 => n67807, A2 => n63174, B1 => n68215, B2 => 
                           n67799, ZN => n6195);
   U47635 : OAI22_X1 port map( A1 => n67807, A2 => n63173, B1 => n68218, B2 => 
                           n67799, ZN => n6196);
   U47636 : OAI22_X1 port map( A1 => n67807, A2 => n63172, B1 => n68221, B2 => 
                           n67799, ZN => n6197);
   U47637 : OAI22_X1 port map( A1 => n67807, A2 => n63171, B1 => n68224, B2 => 
                           n67799, ZN => n6198);
   U47638 : OAI22_X1 port map( A1 => n67807, A2 => n63170, B1 => n68227, B2 => 
                           n67799, ZN => n6199);
   U47639 : OAI22_X1 port map( A1 => n67807, A2 => n63169, B1 => n68230, B2 => 
                           n67799, ZN => n6200);
   U47640 : OAI22_X1 port map( A1 => n67807, A2 => n63168, B1 => n68233, B2 => 
                           n67799, ZN => n6201);
   U47641 : OAI22_X1 port map( A1 => n67807, A2 => n63167, B1 => n68236, B2 => 
                           n67799, ZN => n6202);
   U47642 : OAI22_X1 port map( A1 => n67854, A2 => n63024, B1 => n68059, B2 => 
                           n67846, ZN => n6399);
   U47643 : OAI22_X1 port map( A1 => n67854, A2 => n63023, B1 => n68062, B2 => 
                           n67846, ZN => n6400);
   U47644 : OAI22_X1 port map( A1 => n67854, A2 => n63022, B1 => n68065, B2 => 
                           n67846, ZN => n6401);
   U47645 : OAI22_X1 port map( A1 => n67854, A2 => n63021, B1 => n68068, B2 => 
                           n67846, ZN => n6402);
   U47646 : OAI22_X1 port map( A1 => n67854, A2 => n63020, B1 => n68071, B2 => 
                           n67846, ZN => n6403);
   U47647 : OAI22_X1 port map( A1 => n67854, A2 => n63019, B1 => n68074, B2 => 
                           n67846, ZN => n6404);
   U47648 : OAI22_X1 port map( A1 => n67854, A2 => n63018, B1 => n68077, B2 => 
                           n67846, ZN => n6405);
   U47649 : OAI22_X1 port map( A1 => n67854, A2 => n63017, B1 => n68080, B2 => 
                           n67846, ZN => n6406);
   U47650 : OAI22_X1 port map( A1 => n67854, A2 => n63016, B1 => n68083, B2 => 
                           n67846, ZN => n6407);
   U47651 : OAI22_X1 port map( A1 => n67854, A2 => n63015, B1 => n68086, B2 => 
                           n67846, ZN => n6408);
   U47652 : OAI22_X1 port map( A1 => n67854, A2 => n63014, B1 => n68089, B2 => 
                           n67846, ZN => n6409);
   U47653 : OAI22_X1 port map( A1 => n67854, A2 => n63013, B1 => n68092, B2 => 
                           n67846, ZN => n6410);
   U47654 : OAI22_X1 port map( A1 => n67855, A2 => n63012, B1 => n68095, B2 => 
                           n67847, ZN => n6411);
   U47655 : OAI22_X1 port map( A1 => n67855, A2 => n63011, B1 => n68098, B2 => 
                           n67847, ZN => n6412);
   U47656 : OAI22_X1 port map( A1 => n67855, A2 => n63010, B1 => n68101, B2 => 
                           n67847, ZN => n6413);
   U47657 : OAI22_X1 port map( A1 => n67855, A2 => n63009, B1 => n68104, B2 => 
                           n67847, ZN => n6414);
   U47658 : OAI22_X1 port map( A1 => n67855, A2 => n63008, B1 => n68107, B2 => 
                           n67847, ZN => n6415);
   U47659 : OAI22_X1 port map( A1 => n67855, A2 => n63007, B1 => n68110, B2 => 
                           n67847, ZN => n6416);
   U47660 : OAI22_X1 port map( A1 => n67855, A2 => n63006, B1 => n68113, B2 => 
                           n67847, ZN => n6417);
   U47661 : OAI22_X1 port map( A1 => n67855, A2 => n63005, B1 => n68116, B2 => 
                           n67847, ZN => n6418);
   U47662 : OAI22_X1 port map( A1 => n67855, A2 => n63004, B1 => n68119, B2 => 
                           n67847, ZN => n6419);
   U47663 : OAI22_X1 port map( A1 => n67855, A2 => n63003, B1 => n68122, B2 => 
                           n67847, ZN => n6420);
   U47664 : OAI22_X1 port map( A1 => n67855, A2 => n63002, B1 => n68125, B2 => 
                           n67847, ZN => n6421);
   U47665 : OAI22_X1 port map( A1 => n67855, A2 => n63001, B1 => n68128, B2 => 
                           n67847, ZN => n6422);
   U47666 : OAI22_X1 port map( A1 => n67855, A2 => n63000, B1 => n68131, B2 => 
                           n67848, ZN => n6423);
   U47667 : OAI22_X1 port map( A1 => n67856, A2 => n62999, B1 => n68134, B2 => 
                           n67848, ZN => n6424);
   U47668 : OAI22_X1 port map( A1 => n67856, A2 => n62998, B1 => n68137, B2 => 
                           n67848, ZN => n6425);
   U47669 : OAI22_X1 port map( A1 => n67856, A2 => n62997, B1 => n68140, B2 => 
                           n67848, ZN => n6426);
   U47670 : OAI22_X1 port map( A1 => n67856, A2 => n62996, B1 => n68143, B2 => 
                           n67848, ZN => n6427);
   U47671 : OAI22_X1 port map( A1 => n67856, A2 => n62995, B1 => n68146, B2 => 
                           n67848, ZN => n6428);
   U47672 : OAI22_X1 port map( A1 => n67856, A2 => n62994, B1 => n68149, B2 => 
                           n67848, ZN => n6429);
   U47673 : OAI22_X1 port map( A1 => n67856, A2 => n62993, B1 => n68152, B2 => 
                           n67848, ZN => n6430);
   U47674 : OAI22_X1 port map( A1 => n67856, A2 => n62992, B1 => n68155, B2 => 
                           n67848, ZN => n6431);
   U47675 : OAI22_X1 port map( A1 => n67856, A2 => n62991, B1 => n68158, B2 => 
                           n67848, ZN => n6432);
   U47676 : OAI22_X1 port map( A1 => n67856, A2 => n62990, B1 => n68161, B2 => 
                           n67848, ZN => n6433);
   U47677 : OAI22_X1 port map( A1 => n67856, A2 => n62989, B1 => n68164, B2 => 
                           n67848, ZN => n6434);
   U47678 : OAI22_X1 port map( A1 => n67856, A2 => n62988, B1 => n68167, B2 => 
                           n67849, ZN => n6435);
   U47679 : OAI22_X1 port map( A1 => n67856, A2 => n62987, B1 => n68170, B2 => 
                           n67849, ZN => n6436);
   U47680 : OAI22_X1 port map( A1 => n67857, A2 => n62986, B1 => n68173, B2 => 
                           n67849, ZN => n6437);
   U47681 : OAI22_X1 port map( A1 => n67857, A2 => n62985, B1 => n68176, B2 => 
                           n67849, ZN => n6438);
   U47682 : OAI22_X1 port map( A1 => n67857, A2 => n62984, B1 => n68179, B2 => 
                           n67849, ZN => n6439);
   U47683 : OAI22_X1 port map( A1 => n67857, A2 => n62983, B1 => n68182, B2 => 
                           n67849, ZN => n6440);
   U47684 : OAI22_X1 port map( A1 => n67857, A2 => n62982, B1 => n68185, B2 => 
                           n67849, ZN => n6441);
   U47685 : OAI22_X1 port map( A1 => n67857, A2 => n62981, B1 => n68188, B2 => 
                           n67849, ZN => n6442);
   U47686 : OAI22_X1 port map( A1 => n67857, A2 => n62980, B1 => n68191, B2 => 
                           n67849, ZN => n6443);
   U47687 : OAI22_X1 port map( A1 => n67857, A2 => n62979, B1 => n68194, B2 => 
                           n67849, ZN => n6444);
   U47688 : OAI22_X1 port map( A1 => n67857, A2 => n62978, B1 => n68197, B2 => 
                           n67849, ZN => n6445);
   U47689 : OAI22_X1 port map( A1 => n67857, A2 => n62977, B1 => n68200, B2 => 
                           n67849, ZN => n6446);
   U47690 : OAI22_X1 port map( A1 => n67857, A2 => n62976, B1 => n68203, B2 => 
                           n67850, ZN => n6447);
   U47691 : OAI22_X1 port map( A1 => n67857, A2 => n62975, B1 => n68206, B2 => 
                           n67850, ZN => n6448);
   U47692 : OAI22_X1 port map( A1 => n67857, A2 => n62974, B1 => n68209, B2 => 
                           n67850, ZN => n6449);
   U47693 : OAI22_X1 port map( A1 => n67858, A2 => n62973, B1 => n68212, B2 => 
                           n67850, ZN => n6450);
   U47694 : OAI22_X1 port map( A1 => n67858, A2 => n62972, B1 => n68215, B2 => 
                           n67850, ZN => n6451);
   U47695 : OAI22_X1 port map( A1 => n67858, A2 => n62971, B1 => n68218, B2 => 
                           n67850, ZN => n6452);
   U47696 : OAI22_X1 port map( A1 => n67858, A2 => n62970, B1 => n68221, B2 => 
                           n67850, ZN => n6453);
   U47697 : OAI22_X1 port map( A1 => n67858, A2 => n62969, B1 => n68224, B2 => 
                           n67850, ZN => n6454);
   U47698 : OAI22_X1 port map( A1 => n67858, A2 => n62968, B1 => n68227, B2 => 
                           n67850, ZN => n6455);
   U47699 : OAI22_X1 port map( A1 => n67858, A2 => n62967, B1 => n68230, B2 => 
                           n67850, ZN => n6456);
   U47700 : OAI22_X1 port map( A1 => n67858, A2 => n62966, B1 => n68233, B2 => 
                           n67850, ZN => n6457);
   U47701 : OAI22_X1 port map( A1 => n67858, A2 => n62965, B1 => n68236, B2 => 
                           n67850, ZN => n6458);
   U47702 : OAI22_X1 port map( A1 => n67841, A2 => n63091, B1 => n68059, B2 => 
                           n67833, ZN => n6335);
   U47703 : OAI22_X1 port map( A1 => n67841, A2 => n63090, B1 => n68062, B2 => 
                           n67833, ZN => n6336);
   U47704 : OAI22_X1 port map( A1 => n67841, A2 => n63089, B1 => n68065, B2 => 
                           n67833, ZN => n6337);
   U47705 : OAI22_X1 port map( A1 => n67841, A2 => n63088, B1 => n68068, B2 => 
                           n67833, ZN => n6338);
   U47706 : OAI22_X1 port map( A1 => n67841, A2 => n63087, B1 => n68071, B2 => 
                           n67833, ZN => n6339);
   U47707 : OAI22_X1 port map( A1 => n67841, A2 => n63086, B1 => n68074, B2 => 
                           n67833, ZN => n6340);
   U47708 : OAI22_X1 port map( A1 => n67841, A2 => n63085, B1 => n68077, B2 => 
                           n67833, ZN => n6341);
   U47709 : OAI22_X1 port map( A1 => n67841, A2 => n63084, B1 => n68080, B2 => 
                           n67833, ZN => n6342);
   U47710 : OAI22_X1 port map( A1 => n67841, A2 => n63083, B1 => n68083, B2 => 
                           n67833, ZN => n6343);
   U47711 : OAI22_X1 port map( A1 => n67841, A2 => n63082, B1 => n68086, B2 => 
                           n67833, ZN => n6344);
   U47712 : OAI22_X1 port map( A1 => n67841, A2 => n63081, B1 => n68089, B2 => 
                           n67833, ZN => n6345);
   U47713 : OAI22_X1 port map( A1 => n67841, A2 => n63080, B1 => n68092, B2 => 
                           n67833, ZN => n6346);
   U47714 : OAI22_X1 port map( A1 => n67842, A2 => n63079, B1 => n68095, B2 => 
                           n67834, ZN => n6347);
   U47715 : OAI22_X1 port map( A1 => n67842, A2 => n63078, B1 => n68098, B2 => 
                           n67834, ZN => n6348);
   U47716 : OAI22_X1 port map( A1 => n67842, A2 => n63077, B1 => n68101, B2 => 
                           n67834, ZN => n6349);
   U47717 : OAI22_X1 port map( A1 => n67842, A2 => n63076, B1 => n68104, B2 => 
                           n67834, ZN => n6350);
   U47718 : OAI22_X1 port map( A1 => n67842, A2 => n63075, B1 => n68107, B2 => 
                           n67834, ZN => n6351);
   U47719 : OAI22_X1 port map( A1 => n67842, A2 => n63074, B1 => n68110, B2 => 
                           n67834, ZN => n6352);
   U47720 : OAI22_X1 port map( A1 => n67842, A2 => n63073, B1 => n68113, B2 => 
                           n67834, ZN => n6353);
   U47721 : OAI22_X1 port map( A1 => n67842, A2 => n63072, B1 => n68116, B2 => 
                           n67834, ZN => n6354);
   U47722 : OAI22_X1 port map( A1 => n67842, A2 => n63071, B1 => n68119, B2 => 
                           n67834, ZN => n6355);
   U47723 : OAI22_X1 port map( A1 => n67842, A2 => n63070, B1 => n68122, B2 => 
                           n67834, ZN => n6356);
   U47724 : OAI22_X1 port map( A1 => n67842, A2 => n63069, B1 => n68125, B2 => 
                           n67834, ZN => n6357);
   U47725 : OAI22_X1 port map( A1 => n67842, A2 => n63068, B1 => n68128, B2 => 
                           n67834, ZN => n6358);
   U47726 : OAI22_X1 port map( A1 => n67842, A2 => n63067, B1 => n68131, B2 => 
                           n67835, ZN => n6359);
   U47727 : OAI22_X1 port map( A1 => n67843, A2 => n63066, B1 => n68134, B2 => 
                           n67835, ZN => n6360);
   U47728 : OAI22_X1 port map( A1 => n67843, A2 => n63065, B1 => n68137, B2 => 
                           n67835, ZN => n6361);
   U47729 : OAI22_X1 port map( A1 => n67843, A2 => n63064, B1 => n68140, B2 => 
                           n67835, ZN => n6362);
   U47730 : OAI22_X1 port map( A1 => n67843, A2 => n63063, B1 => n68143, B2 => 
                           n67835, ZN => n6363);
   U47731 : OAI22_X1 port map( A1 => n67843, A2 => n63062, B1 => n68146, B2 => 
                           n67835, ZN => n6364);
   U47732 : OAI22_X1 port map( A1 => n67843, A2 => n63061, B1 => n68149, B2 => 
                           n67835, ZN => n6365);
   U47733 : OAI22_X1 port map( A1 => n67843, A2 => n63060, B1 => n68152, B2 => 
                           n67835, ZN => n6366);
   U47734 : OAI22_X1 port map( A1 => n67843, A2 => n63059, B1 => n68155, B2 => 
                           n67835, ZN => n6367);
   U47735 : OAI22_X1 port map( A1 => n67843, A2 => n63058, B1 => n68158, B2 => 
                           n67835, ZN => n6368);
   U47736 : OAI22_X1 port map( A1 => n67843, A2 => n63057, B1 => n68161, B2 => 
                           n67835, ZN => n6369);
   U47737 : OAI22_X1 port map( A1 => n67843, A2 => n63056, B1 => n68164, B2 => 
                           n67835, ZN => n6370);
   U47738 : OAI22_X1 port map( A1 => n67843, A2 => n63055, B1 => n68167, B2 => 
                           n67836, ZN => n6371);
   U47739 : OAI22_X1 port map( A1 => n67843, A2 => n63054, B1 => n68170, B2 => 
                           n67836, ZN => n6372);
   U47740 : OAI22_X1 port map( A1 => n67844, A2 => n63053, B1 => n68173, B2 => 
                           n67836, ZN => n6373);
   U47741 : OAI22_X1 port map( A1 => n67844, A2 => n63052, B1 => n68176, B2 => 
                           n67836, ZN => n6374);
   U47742 : OAI22_X1 port map( A1 => n67844, A2 => n63051, B1 => n68179, B2 => 
                           n67836, ZN => n6375);
   U47743 : OAI22_X1 port map( A1 => n67844, A2 => n63050, B1 => n68182, B2 => 
                           n67836, ZN => n6376);
   U47744 : OAI22_X1 port map( A1 => n67844, A2 => n63049, B1 => n68185, B2 => 
                           n67836, ZN => n6377);
   U47745 : OAI22_X1 port map( A1 => n67844, A2 => n63048, B1 => n68188, B2 => 
                           n67836, ZN => n6378);
   U47746 : OAI22_X1 port map( A1 => n67844, A2 => n63047, B1 => n68191, B2 => 
                           n67836, ZN => n6379);
   U47747 : OAI22_X1 port map( A1 => n67844, A2 => n63046, B1 => n68194, B2 => 
                           n67836, ZN => n6380);
   U47748 : OAI22_X1 port map( A1 => n67844, A2 => n63045, B1 => n68197, B2 => 
                           n67836, ZN => n6381);
   U47749 : OAI22_X1 port map( A1 => n67844, A2 => n63044, B1 => n68200, B2 => 
                           n67836, ZN => n6382);
   U47750 : OAI22_X1 port map( A1 => n67844, A2 => n63043, B1 => n68203, B2 => 
                           n67837, ZN => n6383);
   U47751 : OAI22_X1 port map( A1 => n67844, A2 => n63042, B1 => n68206, B2 => 
                           n67837, ZN => n6384);
   U47752 : OAI22_X1 port map( A1 => n67844, A2 => n63041, B1 => n68209, B2 => 
                           n67837, ZN => n6385);
   U47753 : OAI22_X1 port map( A1 => n67845, A2 => n63040, B1 => n68212, B2 => 
                           n67837, ZN => n6386);
   U47754 : OAI22_X1 port map( A1 => n67845, A2 => n63039, B1 => n68215, B2 => 
                           n67837, ZN => n6387);
   U47755 : OAI22_X1 port map( A1 => n67845, A2 => n63038, B1 => n68218, B2 => 
                           n67837, ZN => n6388);
   U47756 : OAI22_X1 port map( A1 => n67845, A2 => n63037, B1 => n68221, B2 => 
                           n67837, ZN => n6389);
   U47757 : OAI22_X1 port map( A1 => n67845, A2 => n63036, B1 => n68224, B2 => 
                           n67837, ZN => n6390);
   U47758 : OAI22_X1 port map( A1 => n67845, A2 => n63035, B1 => n68227, B2 => 
                           n67837, ZN => n6391);
   U47759 : OAI22_X1 port map( A1 => n67845, A2 => n63034, B1 => n68230, B2 => 
                           n67837, ZN => n6392);
   U47760 : OAI22_X1 port map( A1 => n67845, A2 => n63033, B1 => n68233, B2 => 
                           n67837, ZN => n6393);
   U47761 : OAI22_X1 port map( A1 => n67845, A2 => n63032, B1 => n68236, B2 => 
                           n67837, ZN => n6394);
   U47762 : OAI22_X1 port map( A1 => n67752, A2 => n63427, B1 => n68059, B2 => 
                           n67744, ZN => n5887);
   U47763 : OAI22_X1 port map( A1 => n67752, A2 => n63426, B1 => n68062, B2 => 
                           n67744, ZN => n5888);
   U47764 : OAI22_X1 port map( A1 => n67752, A2 => n63425, B1 => n68065, B2 => 
                           n67744, ZN => n5889);
   U47765 : OAI22_X1 port map( A1 => n67752, A2 => n63424, B1 => n68068, B2 => 
                           n67744, ZN => n5890);
   U47766 : OAI22_X1 port map( A1 => n67752, A2 => n63423, B1 => n68071, B2 => 
                           n67744, ZN => n5891);
   U47767 : OAI22_X1 port map( A1 => n67752, A2 => n63422, B1 => n68074, B2 => 
                           n67744, ZN => n5892);
   U47768 : OAI22_X1 port map( A1 => n67752, A2 => n63421, B1 => n68077, B2 => 
                           n67744, ZN => n5893);
   U47769 : OAI22_X1 port map( A1 => n67752, A2 => n63420, B1 => n68080, B2 => 
                           n67744, ZN => n5894);
   U47770 : OAI22_X1 port map( A1 => n67752, A2 => n63419, B1 => n68083, B2 => 
                           n67744, ZN => n5895);
   U47771 : OAI22_X1 port map( A1 => n67752, A2 => n63418, B1 => n68086, B2 => 
                           n67744, ZN => n5896);
   U47772 : OAI22_X1 port map( A1 => n67752, A2 => n63417, B1 => n68089, B2 => 
                           n67744, ZN => n5897);
   U47773 : OAI22_X1 port map( A1 => n67752, A2 => n63416, B1 => n68092, B2 => 
                           n67744, ZN => n5898);
   U47774 : OAI22_X1 port map( A1 => n67753, A2 => n63415, B1 => n68095, B2 => 
                           n67745, ZN => n5899);
   U47775 : OAI22_X1 port map( A1 => n67753, A2 => n63414, B1 => n68098, B2 => 
                           n67745, ZN => n5900);
   U47776 : OAI22_X1 port map( A1 => n67753, A2 => n63413, B1 => n68101, B2 => 
                           n67745, ZN => n5901);
   U47777 : OAI22_X1 port map( A1 => n67753, A2 => n63412, B1 => n68104, B2 => 
                           n67745, ZN => n5902);
   U47778 : OAI22_X1 port map( A1 => n67753, A2 => n63411, B1 => n68107, B2 => 
                           n67745, ZN => n5903);
   U47779 : OAI22_X1 port map( A1 => n67753, A2 => n63410, B1 => n68110, B2 => 
                           n67745, ZN => n5904);
   U47780 : OAI22_X1 port map( A1 => n67753, A2 => n63409, B1 => n68113, B2 => 
                           n67745, ZN => n5905);
   U47781 : OAI22_X1 port map( A1 => n67753, A2 => n63408, B1 => n68116, B2 => 
                           n67745, ZN => n5906);
   U47782 : OAI22_X1 port map( A1 => n67753, A2 => n63407, B1 => n68119, B2 => 
                           n67745, ZN => n5907);
   U47783 : OAI22_X1 port map( A1 => n67753, A2 => n63406, B1 => n68122, B2 => 
                           n67745, ZN => n5908);
   U47784 : OAI22_X1 port map( A1 => n67753, A2 => n63405, B1 => n68125, B2 => 
                           n67745, ZN => n5909);
   U47785 : OAI22_X1 port map( A1 => n67753, A2 => n63404, B1 => n68128, B2 => 
                           n67745, ZN => n5910);
   U47786 : OAI22_X1 port map( A1 => n67753, A2 => n63403, B1 => n68131, B2 => 
                           n67746, ZN => n5911);
   U47787 : OAI22_X1 port map( A1 => n67754, A2 => n63402, B1 => n68134, B2 => 
                           n67746, ZN => n5912);
   U47788 : OAI22_X1 port map( A1 => n67754, A2 => n63401, B1 => n68137, B2 => 
                           n67746, ZN => n5913);
   U47789 : OAI22_X1 port map( A1 => n67754, A2 => n63400, B1 => n68140, B2 => 
                           n67746, ZN => n5914);
   U47790 : OAI22_X1 port map( A1 => n67754, A2 => n63399, B1 => n68143, B2 => 
                           n67746, ZN => n5915);
   U47791 : OAI22_X1 port map( A1 => n67754, A2 => n63398, B1 => n68146, B2 => 
                           n67746, ZN => n5916);
   U47792 : OAI22_X1 port map( A1 => n67754, A2 => n63397, B1 => n68149, B2 => 
                           n67746, ZN => n5917);
   U47793 : OAI22_X1 port map( A1 => n67754, A2 => n63396, B1 => n68152, B2 => 
                           n67746, ZN => n5918);
   U47794 : OAI22_X1 port map( A1 => n67754, A2 => n63395, B1 => n68155, B2 => 
                           n67746, ZN => n5919);
   U47795 : OAI22_X1 port map( A1 => n67754, A2 => n63394, B1 => n68158, B2 => 
                           n67746, ZN => n5920);
   U47796 : OAI22_X1 port map( A1 => n67754, A2 => n63393, B1 => n68161, B2 => 
                           n67746, ZN => n5921);
   U47797 : OAI22_X1 port map( A1 => n67754, A2 => n63392, B1 => n68164, B2 => 
                           n67746, ZN => n5922);
   U47798 : OAI22_X1 port map( A1 => n67754, A2 => n63391, B1 => n68167, B2 => 
                           n67747, ZN => n5923);
   U47799 : OAI22_X1 port map( A1 => n67754, A2 => n63390, B1 => n68170, B2 => 
                           n67747, ZN => n5924);
   U47800 : OAI22_X1 port map( A1 => n67755, A2 => n63389, B1 => n68173, B2 => 
                           n67747, ZN => n5925);
   U47801 : OAI22_X1 port map( A1 => n67755, A2 => n63388, B1 => n68176, B2 => 
                           n67747, ZN => n5926);
   U47802 : OAI22_X1 port map( A1 => n67755, A2 => n63387, B1 => n68179, B2 => 
                           n67747, ZN => n5927);
   U47803 : OAI22_X1 port map( A1 => n67755, A2 => n63386, B1 => n68182, B2 => 
                           n67747, ZN => n5928);
   U47804 : OAI22_X1 port map( A1 => n67755, A2 => n63385, B1 => n68185, B2 => 
                           n67747, ZN => n5929);
   U47805 : OAI22_X1 port map( A1 => n67755, A2 => n63384, B1 => n68188, B2 => 
                           n67747, ZN => n5930);
   U47806 : OAI22_X1 port map( A1 => n67755, A2 => n63383, B1 => n68191, B2 => 
                           n67747, ZN => n5931);
   U47807 : OAI22_X1 port map( A1 => n67755, A2 => n63382, B1 => n68194, B2 => 
                           n67747, ZN => n5932);
   U47808 : OAI22_X1 port map( A1 => n67755, A2 => n63381, B1 => n68197, B2 => 
                           n67747, ZN => n5933);
   U47809 : OAI22_X1 port map( A1 => n67755, A2 => n63380, B1 => n68200, B2 => 
                           n67747, ZN => n5934);
   U47810 : OAI22_X1 port map( A1 => n67755, A2 => n63379, B1 => n68203, B2 => 
                           n67748, ZN => n5935);
   U47811 : OAI22_X1 port map( A1 => n67755, A2 => n63378, B1 => n68206, B2 => 
                           n67748, ZN => n5936);
   U47812 : OAI22_X1 port map( A1 => n67755, A2 => n63377, B1 => n68209, B2 => 
                           n67748, ZN => n5937);
   U47813 : OAI22_X1 port map( A1 => n67756, A2 => n63376, B1 => n68212, B2 => 
                           n67748, ZN => n5938);
   U47814 : OAI22_X1 port map( A1 => n67756, A2 => n63375, B1 => n68215, B2 => 
                           n67748, ZN => n5939);
   U47815 : OAI22_X1 port map( A1 => n67756, A2 => n63374, B1 => n68218, B2 => 
                           n67748, ZN => n5940);
   U47816 : OAI22_X1 port map( A1 => n67756, A2 => n63373, B1 => n68221, B2 => 
                           n67748, ZN => n5941);
   U47817 : OAI22_X1 port map( A1 => n67756, A2 => n63372, B1 => n68224, B2 => 
                           n67748, ZN => n5942);
   U47818 : OAI22_X1 port map( A1 => n67756, A2 => n63371, B1 => n68227, B2 => 
                           n67748, ZN => n5943);
   U47819 : OAI22_X1 port map( A1 => n67756, A2 => n63370, B1 => n68230, B2 => 
                           n67748, ZN => n5944);
   U47820 : OAI22_X1 port map( A1 => n67756, A2 => n63369, B1 => n68233, B2 => 
                           n67748, ZN => n5945);
   U47821 : OAI22_X1 port map( A1 => n67756, A2 => n63368, B1 => n68236, B2 => 
                           n67748, ZN => n5946);
   U47822 : OAI22_X1 port map( A1 => n67880, A2 => n62891, B1 => n68059, B2 => 
                           n67872, ZN => n6527);
   U47823 : OAI22_X1 port map( A1 => n67880, A2 => n62890, B1 => n68062, B2 => 
                           n67872, ZN => n6528);
   U47824 : OAI22_X1 port map( A1 => n67880, A2 => n62889, B1 => n68065, B2 => 
                           n67872, ZN => n6529);
   U47825 : OAI22_X1 port map( A1 => n67880, A2 => n62888, B1 => n68068, B2 => 
                           n67872, ZN => n6530);
   U47826 : OAI22_X1 port map( A1 => n67880, A2 => n62887, B1 => n68071, B2 => 
                           n67872, ZN => n6531);
   U47827 : OAI22_X1 port map( A1 => n67880, A2 => n62886, B1 => n68074, B2 => 
                           n67872, ZN => n6532);
   U47828 : OAI22_X1 port map( A1 => n67880, A2 => n62885, B1 => n68077, B2 => 
                           n67872, ZN => n6533);
   U47829 : OAI22_X1 port map( A1 => n67880, A2 => n62884, B1 => n68080, B2 => 
                           n67872, ZN => n6534);
   U47830 : OAI22_X1 port map( A1 => n67880, A2 => n62883, B1 => n68083, B2 => 
                           n67872, ZN => n6535);
   U47831 : OAI22_X1 port map( A1 => n67880, A2 => n62882, B1 => n68086, B2 => 
                           n67872, ZN => n6536);
   U47832 : OAI22_X1 port map( A1 => n67880, A2 => n62881, B1 => n68089, B2 => 
                           n67872, ZN => n6537);
   U47833 : OAI22_X1 port map( A1 => n67880, A2 => n62880, B1 => n68092, B2 => 
                           n67872, ZN => n6538);
   U47834 : OAI22_X1 port map( A1 => n67881, A2 => n62879, B1 => n68095, B2 => 
                           n67873, ZN => n6539);
   U47835 : OAI22_X1 port map( A1 => n67881, A2 => n62878, B1 => n68098, B2 => 
                           n67873, ZN => n6540);
   U47836 : OAI22_X1 port map( A1 => n67881, A2 => n62877, B1 => n68101, B2 => 
                           n67873, ZN => n6541);
   U47837 : OAI22_X1 port map( A1 => n67881, A2 => n62876, B1 => n68104, B2 => 
                           n67873, ZN => n6542);
   U47838 : OAI22_X1 port map( A1 => n67881, A2 => n62875, B1 => n68107, B2 => 
                           n67873, ZN => n6543);
   U47839 : OAI22_X1 port map( A1 => n67881, A2 => n62874, B1 => n68110, B2 => 
                           n67873, ZN => n6544);
   U47840 : OAI22_X1 port map( A1 => n67881, A2 => n62873, B1 => n68113, B2 => 
                           n67873, ZN => n6545);
   U47841 : OAI22_X1 port map( A1 => n67881, A2 => n62872, B1 => n68116, B2 => 
                           n67873, ZN => n6546);
   U47842 : OAI22_X1 port map( A1 => n67881, A2 => n62871, B1 => n68119, B2 => 
                           n67873, ZN => n6547);
   U47843 : OAI22_X1 port map( A1 => n67881, A2 => n62870, B1 => n68122, B2 => 
                           n67873, ZN => n6548);
   U47844 : OAI22_X1 port map( A1 => n67881, A2 => n62869, B1 => n68125, B2 => 
                           n67873, ZN => n6549);
   U47845 : OAI22_X1 port map( A1 => n67881, A2 => n62868, B1 => n68128, B2 => 
                           n67873, ZN => n6550);
   U47846 : OAI22_X1 port map( A1 => n67881, A2 => n62867, B1 => n68131, B2 => 
                           n67874, ZN => n6551);
   U47847 : OAI22_X1 port map( A1 => n67882, A2 => n62866, B1 => n68134, B2 => 
                           n67874, ZN => n6552);
   U47848 : OAI22_X1 port map( A1 => n67882, A2 => n62865, B1 => n68137, B2 => 
                           n67874, ZN => n6553);
   U47849 : OAI22_X1 port map( A1 => n67882, A2 => n62864, B1 => n68140, B2 => 
                           n67874, ZN => n6554);
   U47850 : OAI22_X1 port map( A1 => n67882, A2 => n62863, B1 => n68143, B2 => 
                           n67874, ZN => n6555);
   U47851 : OAI22_X1 port map( A1 => n67882, A2 => n62862, B1 => n68146, B2 => 
                           n67874, ZN => n6556);
   U47852 : OAI22_X1 port map( A1 => n67882, A2 => n62861, B1 => n68149, B2 => 
                           n67874, ZN => n6557);
   U47853 : OAI22_X1 port map( A1 => n67882, A2 => n62860, B1 => n68152, B2 => 
                           n67874, ZN => n6558);
   U47854 : OAI22_X1 port map( A1 => n67882, A2 => n62859, B1 => n68155, B2 => 
                           n67874, ZN => n6559);
   U47855 : OAI22_X1 port map( A1 => n67882, A2 => n62858, B1 => n68158, B2 => 
                           n67874, ZN => n6560);
   U47856 : OAI22_X1 port map( A1 => n67882, A2 => n62857, B1 => n68161, B2 => 
                           n67874, ZN => n6561);
   U47857 : OAI22_X1 port map( A1 => n67882, A2 => n62856, B1 => n68164, B2 => 
                           n67874, ZN => n6562);
   U47858 : OAI22_X1 port map( A1 => n67882, A2 => n62855, B1 => n68167, B2 => 
                           n67875, ZN => n6563);
   U47859 : OAI22_X1 port map( A1 => n67882, A2 => n62854, B1 => n68170, B2 => 
                           n67875, ZN => n6564);
   U47860 : OAI22_X1 port map( A1 => n67883, A2 => n62853, B1 => n68173, B2 => 
                           n67875, ZN => n6565);
   U47861 : OAI22_X1 port map( A1 => n67883, A2 => n62852, B1 => n68176, B2 => 
                           n67875, ZN => n6566);
   U47862 : OAI22_X1 port map( A1 => n67883, A2 => n62851, B1 => n68179, B2 => 
                           n67875, ZN => n6567);
   U47863 : OAI22_X1 port map( A1 => n67883, A2 => n62850, B1 => n68182, B2 => 
                           n67875, ZN => n6568);
   U47864 : OAI22_X1 port map( A1 => n67883, A2 => n62849, B1 => n68185, B2 => 
                           n67875, ZN => n6569);
   U47865 : OAI22_X1 port map( A1 => n67883, A2 => n62848, B1 => n68188, B2 => 
                           n67875, ZN => n6570);
   U47866 : OAI22_X1 port map( A1 => n67883, A2 => n62847, B1 => n68191, B2 => 
                           n67875, ZN => n6571);
   U47867 : OAI22_X1 port map( A1 => n67883, A2 => n62846, B1 => n68194, B2 => 
                           n67875, ZN => n6572);
   U47868 : OAI22_X1 port map( A1 => n67883, A2 => n62845, B1 => n68197, B2 => 
                           n67875, ZN => n6573);
   U47869 : OAI22_X1 port map( A1 => n67883, A2 => n62844, B1 => n68200, B2 => 
                           n67875, ZN => n6574);
   U47870 : OAI22_X1 port map( A1 => n67883, A2 => n62843, B1 => n68203, B2 => 
                           n67876, ZN => n6575);
   U47871 : OAI22_X1 port map( A1 => n67883, A2 => n62842, B1 => n68206, B2 => 
                           n67876, ZN => n6576);
   U47872 : OAI22_X1 port map( A1 => n67883, A2 => n62841, B1 => n68209, B2 => 
                           n67876, ZN => n6577);
   U47873 : OAI22_X1 port map( A1 => n67884, A2 => n62840, B1 => n68212, B2 => 
                           n67876, ZN => n6578);
   U47874 : OAI22_X1 port map( A1 => n67884, A2 => n62839, B1 => n68215, B2 => 
                           n67876, ZN => n6579);
   U47875 : OAI22_X1 port map( A1 => n67884, A2 => n62838, B1 => n68218, B2 => 
                           n67876, ZN => n6580);
   U47876 : OAI22_X1 port map( A1 => n67884, A2 => n62837, B1 => n68221, B2 => 
                           n67876, ZN => n6581);
   U47877 : OAI22_X1 port map( A1 => n67884, A2 => n62836, B1 => n68224, B2 => 
                           n67876, ZN => n6582);
   U47878 : OAI22_X1 port map( A1 => n67884, A2 => n62835, B1 => n68227, B2 => 
                           n67876, ZN => n6583);
   U47879 : OAI22_X1 port map( A1 => n67884, A2 => n62834, B1 => n68230, B2 => 
                           n67876, ZN => n6584);
   U47880 : OAI22_X1 port map( A1 => n67884, A2 => n62833, B1 => n68233, B2 => 
                           n67876, ZN => n6585);
   U47881 : OAI22_X1 port map( A1 => n67884, A2 => n62832, B1 => n68236, B2 => 
                           n67876, ZN => n6586);
   U47882 : OAI22_X1 port map( A1 => n68034, A2 => n62222, B1 => n68058, B2 => 
                           n68026, ZN => n7295);
   U47883 : OAI22_X1 port map( A1 => n68034, A2 => n62221, B1 => n68061, B2 => 
                           n68026, ZN => n7296);
   U47884 : OAI22_X1 port map( A1 => n68034, A2 => n62220, B1 => n68064, B2 => 
                           n68026, ZN => n7297);
   U47885 : OAI22_X1 port map( A1 => n68034, A2 => n62219, B1 => n68067, B2 => 
                           n68026, ZN => n7298);
   U47886 : OAI22_X1 port map( A1 => n68034, A2 => n62218, B1 => n68070, B2 => 
                           n68026, ZN => n7299);
   U47887 : OAI22_X1 port map( A1 => n68034, A2 => n62217, B1 => n68073, B2 => 
                           n68026, ZN => n7300);
   U47888 : OAI22_X1 port map( A1 => n68034, A2 => n62216, B1 => n68076, B2 => 
                           n68026, ZN => n7301);
   U47889 : OAI22_X1 port map( A1 => n68034, A2 => n62215, B1 => n68079, B2 => 
                           n68026, ZN => n7302);
   U47890 : OAI22_X1 port map( A1 => n68034, A2 => n62214, B1 => n68082, B2 => 
                           n68026, ZN => n7303);
   U47891 : OAI22_X1 port map( A1 => n68034, A2 => n62213, B1 => n68085, B2 => 
                           n68026, ZN => n7304);
   U47892 : OAI22_X1 port map( A1 => n68034, A2 => n62212, B1 => n68088, B2 => 
                           n68026, ZN => n7305);
   U47893 : OAI22_X1 port map( A1 => n68034, A2 => n62211, B1 => n68091, B2 => 
                           n68026, ZN => n7306);
   U47894 : OAI22_X1 port map( A1 => n68035, A2 => n62210, B1 => n68094, B2 => 
                           n68027, ZN => n7307);
   U47895 : OAI22_X1 port map( A1 => n68035, A2 => n62209, B1 => n68097, B2 => 
                           n68027, ZN => n7308);
   U47896 : OAI22_X1 port map( A1 => n68035, A2 => n62208, B1 => n68100, B2 => 
                           n68027, ZN => n7309);
   U47897 : OAI22_X1 port map( A1 => n68035, A2 => n62207, B1 => n68103, B2 => 
                           n68027, ZN => n7310);
   U47898 : OAI22_X1 port map( A1 => n68035, A2 => n62206, B1 => n68106, B2 => 
                           n68027, ZN => n7311);
   U47899 : OAI22_X1 port map( A1 => n68035, A2 => n62205, B1 => n68109, B2 => 
                           n68027, ZN => n7312);
   U47900 : OAI22_X1 port map( A1 => n68035, A2 => n62204, B1 => n68112, B2 => 
                           n68027, ZN => n7313);
   U47901 : OAI22_X1 port map( A1 => n68035, A2 => n62203, B1 => n68115, B2 => 
                           n68027, ZN => n7314);
   U47902 : OAI22_X1 port map( A1 => n68035, A2 => n62202, B1 => n68118, B2 => 
                           n68027, ZN => n7315);
   U47903 : OAI22_X1 port map( A1 => n68035, A2 => n62201, B1 => n68121, B2 => 
                           n68027, ZN => n7316);
   U47904 : OAI22_X1 port map( A1 => n68035, A2 => n62200, B1 => n68124, B2 => 
                           n68027, ZN => n7317);
   U47905 : OAI22_X1 port map( A1 => n68035, A2 => n62199, B1 => n68127, B2 => 
                           n68027, ZN => n7318);
   U47906 : OAI22_X1 port map( A1 => n68035, A2 => n62198, B1 => n68130, B2 => 
                           n68028, ZN => n7319);
   U47907 : OAI22_X1 port map( A1 => n68036, A2 => n62197, B1 => n68133, B2 => 
                           n68028, ZN => n7320);
   U47908 : OAI22_X1 port map( A1 => n68036, A2 => n62196, B1 => n68136, B2 => 
                           n68028, ZN => n7321);
   U47909 : OAI22_X1 port map( A1 => n68036, A2 => n62195, B1 => n68139, B2 => 
                           n68028, ZN => n7322);
   U47910 : OAI22_X1 port map( A1 => n68036, A2 => n62194, B1 => n68142, B2 => 
                           n68028, ZN => n7323);
   U47911 : OAI22_X1 port map( A1 => n68036, A2 => n62193, B1 => n68145, B2 => 
                           n68028, ZN => n7324);
   U47912 : OAI22_X1 port map( A1 => n68036, A2 => n62192, B1 => n68148, B2 => 
                           n68028, ZN => n7325);
   U47913 : OAI22_X1 port map( A1 => n68036, A2 => n62191, B1 => n68151, B2 => 
                           n68028, ZN => n7326);
   U47914 : OAI22_X1 port map( A1 => n68036, A2 => n62190, B1 => n68154, B2 => 
                           n68028, ZN => n7327);
   U47915 : OAI22_X1 port map( A1 => n68036, A2 => n62189, B1 => n68157, B2 => 
                           n68028, ZN => n7328);
   U47916 : OAI22_X1 port map( A1 => n68036, A2 => n62188, B1 => n68160, B2 => 
                           n68028, ZN => n7329);
   U47917 : OAI22_X1 port map( A1 => n68036, A2 => n62187, B1 => n68163, B2 => 
                           n68028, ZN => n7330);
   U47918 : OAI22_X1 port map( A1 => n68036, A2 => n62186, B1 => n68166, B2 => 
                           n68029, ZN => n7331);
   U47919 : OAI22_X1 port map( A1 => n68036, A2 => n62185, B1 => n68169, B2 => 
                           n68029, ZN => n7332);
   U47920 : OAI22_X1 port map( A1 => n68037, A2 => n62184, B1 => n68172, B2 => 
                           n68029, ZN => n7333);
   U47921 : OAI22_X1 port map( A1 => n68037, A2 => n62183, B1 => n68175, B2 => 
                           n68029, ZN => n7334);
   U47922 : OAI22_X1 port map( A1 => n68037, A2 => n62182, B1 => n68178, B2 => 
                           n68029, ZN => n7335);
   U47923 : OAI22_X1 port map( A1 => n68037, A2 => n62181, B1 => n68181, B2 => 
                           n68029, ZN => n7336);
   U47924 : OAI22_X1 port map( A1 => n68037, A2 => n62180, B1 => n68184, B2 => 
                           n68029, ZN => n7337);
   U47925 : OAI22_X1 port map( A1 => n68037, A2 => n62179, B1 => n68187, B2 => 
                           n68029, ZN => n7338);
   U47926 : OAI22_X1 port map( A1 => n68037, A2 => n62178, B1 => n68190, B2 => 
                           n68029, ZN => n7339);
   U47927 : OAI22_X1 port map( A1 => n68037, A2 => n62177, B1 => n68193, B2 => 
                           n68029, ZN => n7340);
   U47928 : OAI22_X1 port map( A1 => n68037, A2 => n62176, B1 => n68196, B2 => 
                           n68029, ZN => n7341);
   U47929 : OAI22_X1 port map( A1 => n68037, A2 => n62175, B1 => n68199, B2 => 
                           n68029, ZN => n7342);
   U47930 : OAI22_X1 port map( A1 => n68037, A2 => n62174, B1 => n68202, B2 => 
                           n68030, ZN => n7343);
   U47931 : OAI22_X1 port map( A1 => n68037, A2 => n62173, B1 => n68205, B2 => 
                           n68030, ZN => n7344);
   U47932 : OAI22_X1 port map( A1 => n68037, A2 => n62172, B1 => n68208, B2 => 
                           n68030, ZN => n7345);
   U47933 : OAI22_X1 port map( A1 => n68038, A2 => n62171, B1 => n68211, B2 => 
                           n68030, ZN => n7346);
   U47934 : OAI22_X1 port map( A1 => n68038, A2 => n62170, B1 => n68214, B2 => 
                           n68030, ZN => n7347);
   U47935 : OAI22_X1 port map( A1 => n68038, A2 => n62169, B1 => n68217, B2 => 
                           n68030, ZN => n7348);
   U47936 : OAI22_X1 port map( A1 => n68038, A2 => n62168, B1 => n68220, B2 => 
                           n68030, ZN => n7349);
   U47937 : OAI22_X1 port map( A1 => n68038, A2 => n62167, B1 => n68223, B2 => 
                           n68030, ZN => n7350);
   U47938 : OAI22_X1 port map( A1 => n68038, A2 => n62166, B1 => n68226, B2 => 
                           n68030, ZN => n7351);
   U47939 : OAI22_X1 port map( A1 => n68038, A2 => n62165, B1 => n68229, B2 => 
                           n68030, ZN => n7352);
   U47940 : OAI22_X1 port map( A1 => n68038, A2 => n62164, B1 => n68232, B2 => 
                           n68030, ZN => n7353);
   U47941 : OAI22_X1 port map( A1 => n68038, A2 => n62163, B1 => n68235, B2 => 
                           n68030, ZN => n7354);
   U47942 : OAI22_X1 port map( A1 => n68021, A2 => n62289, B1 => n68058, B2 => 
                           n68013, ZN => n7231);
   U47943 : OAI22_X1 port map( A1 => n68021, A2 => n62288, B1 => n68061, B2 => 
                           n68013, ZN => n7232);
   U47944 : OAI22_X1 port map( A1 => n68021, A2 => n62287, B1 => n68064, B2 => 
                           n68013, ZN => n7233);
   U47945 : OAI22_X1 port map( A1 => n68021, A2 => n62286, B1 => n68067, B2 => 
                           n68013, ZN => n7234);
   U47946 : OAI22_X1 port map( A1 => n68021, A2 => n62285, B1 => n68070, B2 => 
                           n68013, ZN => n7235);
   U47947 : OAI22_X1 port map( A1 => n68021, A2 => n62284, B1 => n68073, B2 => 
                           n68013, ZN => n7236);
   U47948 : OAI22_X1 port map( A1 => n68021, A2 => n62283, B1 => n68076, B2 => 
                           n68013, ZN => n7237);
   U47949 : OAI22_X1 port map( A1 => n68021, A2 => n62282, B1 => n68079, B2 => 
                           n68013, ZN => n7238);
   U47950 : OAI22_X1 port map( A1 => n68021, A2 => n62281, B1 => n68082, B2 => 
                           n68013, ZN => n7239);
   U47951 : OAI22_X1 port map( A1 => n68021, A2 => n62280, B1 => n68085, B2 => 
                           n68013, ZN => n7240);
   U47952 : OAI22_X1 port map( A1 => n68021, A2 => n62279, B1 => n68088, B2 => 
                           n68013, ZN => n7241);
   U47953 : OAI22_X1 port map( A1 => n68021, A2 => n62278, B1 => n68091, B2 => 
                           n68013, ZN => n7242);
   U47954 : OAI22_X1 port map( A1 => n68022, A2 => n62277, B1 => n68094, B2 => 
                           n68014, ZN => n7243);
   U47955 : OAI22_X1 port map( A1 => n68022, A2 => n62276, B1 => n68097, B2 => 
                           n68014, ZN => n7244);
   U47956 : OAI22_X1 port map( A1 => n68022, A2 => n62275, B1 => n68100, B2 => 
                           n68014, ZN => n7245);
   U47957 : OAI22_X1 port map( A1 => n68022, A2 => n62274, B1 => n68103, B2 => 
                           n68014, ZN => n7246);
   U47958 : OAI22_X1 port map( A1 => n68022, A2 => n62273, B1 => n68106, B2 => 
                           n68014, ZN => n7247);
   U47959 : OAI22_X1 port map( A1 => n68022, A2 => n62272, B1 => n68109, B2 => 
                           n68014, ZN => n7248);
   U47960 : OAI22_X1 port map( A1 => n68022, A2 => n62271, B1 => n68112, B2 => 
                           n68014, ZN => n7249);
   U47961 : OAI22_X1 port map( A1 => n68022, A2 => n62270, B1 => n68115, B2 => 
                           n68014, ZN => n7250);
   U47962 : OAI22_X1 port map( A1 => n68022, A2 => n62269, B1 => n68118, B2 => 
                           n68014, ZN => n7251);
   U47963 : OAI22_X1 port map( A1 => n68022, A2 => n62268, B1 => n68121, B2 => 
                           n68014, ZN => n7252);
   U47964 : OAI22_X1 port map( A1 => n68022, A2 => n62267, B1 => n68124, B2 => 
                           n68014, ZN => n7253);
   U47965 : OAI22_X1 port map( A1 => n68022, A2 => n62266, B1 => n68127, B2 => 
                           n68014, ZN => n7254);
   U47966 : OAI22_X1 port map( A1 => n68022, A2 => n62265, B1 => n68130, B2 => 
                           n68015, ZN => n7255);
   U47967 : OAI22_X1 port map( A1 => n68023, A2 => n62264, B1 => n68133, B2 => 
                           n68015, ZN => n7256);
   U47968 : OAI22_X1 port map( A1 => n68023, A2 => n62263, B1 => n68136, B2 => 
                           n68015, ZN => n7257);
   U47969 : OAI22_X1 port map( A1 => n68023, A2 => n62262, B1 => n68139, B2 => 
                           n68015, ZN => n7258);
   U47970 : OAI22_X1 port map( A1 => n68023, A2 => n62261, B1 => n68142, B2 => 
                           n68015, ZN => n7259);
   U47971 : OAI22_X1 port map( A1 => n68023, A2 => n62260, B1 => n68145, B2 => 
                           n68015, ZN => n7260);
   U47972 : OAI22_X1 port map( A1 => n68023, A2 => n62259, B1 => n68148, B2 => 
                           n68015, ZN => n7261);
   U47973 : OAI22_X1 port map( A1 => n68023, A2 => n62258, B1 => n68151, B2 => 
                           n68015, ZN => n7262);
   U47974 : OAI22_X1 port map( A1 => n68023, A2 => n62257, B1 => n68154, B2 => 
                           n68015, ZN => n7263);
   U47975 : OAI22_X1 port map( A1 => n68023, A2 => n62256, B1 => n68157, B2 => 
                           n68015, ZN => n7264);
   U47976 : OAI22_X1 port map( A1 => n68023, A2 => n62255, B1 => n68160, B2 => 
                           n68015, ZN => n7265);
   U47977 : OAI22_X1 port map( A1 => n68023, A2 => n62254, B1 => n68163, B2 => 
                           n68015, ZN => n7266);
   U47978 : OAI22_X1 port map( A1 => n68023, A2 => n62253, B1 => n68166, B2 => 
                           n68016, ZN => n7267);
   U47979 : OAI22_X1 port map( A1 => n68023, A2 => n62252, B1 => n68169, B2 => 
                           n68016, ZN => n7268);
   U47980 : OAI22_X1 port map( A1 => n68024, A2 => n62251, B1 => n68172, B2 => 
                           n68016, ZN => n7269);
   U47981 : OAI22_X1 port map( A1 => n68024, A2 => n62250, B1 => n68175, B2 => 
                           n68016, ZN => n7270);
   U47982 : OAI22_X1 port map( A1 => n68024, A2 => n62249, B1 => n68178, B2 => 
                           n68016, ZN => n7271);
   U47983 : OAI22_X1 port map( A1 => n68024, A2 => n62248, B1 => n68181, B2 => 
                           n68016, ZN => n7272);
   U47984 : OAI22_X1 port map( A1 => n68024, A2 => n62247, B1 => n68184, B2 => 
                           n68016, ZN => n7273);
   U47985 : OAI22_X1 port map( A1 => n68024, A2 => n62246, B1 => n68187, B2 => 
                           n68016, ZN => n7274);
   U47986 : OAI22_X1 port map( A1 => n68024, A2 => n62245, B1 => n68190, B2 => 
                           n68016, ZN => n7275);
   U47987 : OAI22_X1 port map( A1 => n68024, A2 => n62244, B1 => n68193, B2 => 
                           n68016, ZN => n7276);
   U47988 : OAI22_X1 port map( A1 => n68024, A2 => n62243, B1 => n68196, B2 => 
                           n68016, ZN => n7277);
   U47989 : OAI22_X1 port map( A1 => n68024, A2 => n62242, B1 => n68199, B2 => 
                           n68016, ZN => n7278);
   U47990 : OAI22_X1 port map( A1 => n68024, A2 => n62241, B1 => n68202, B2 => 
                           n68017, ZN => n7279);
   U47991 : OAI22_X1 port map( A1 => n68024, A2 => n62240, B1 => n68205, B2 => 
                           n68017, ZN => n7280);
   U47992 : OAI22_X1 port map( A1 => n68024, A2 => n62239, B1 => n68208, B2 => 
                           n68017, ZN => n7281);
   U47993 : OAI22_X1 port map( A1 => n68025, A2 => n62238, B1 => n68211, B2 => 
                           n68017, ZN => n7282);
   U47994 : OAI22_X1 port map( A1 => n68025, A2 => n62237, B1 => n68214, B2 => 
                           n68017, ZN => n7283);
   U47995 : OAI22_X1 port map( A1 => n68025, A2 => n62236, B1 => n68217, B2 => 
                           n68017, ZN => n7284);
   U47996 : OAI22_X1 port map( A1 => n68025, A2 => n62235, B1 => n68220, B2 => 
                           n68017, ZN => n7285);
   U47997 : OAI22_X1 port map( A1 => n68025, A2 => n62234, B1 => n68223, B2 => 
                           n68017, ZN => n7286);
   U47998 : OAI22_X1 port map( A1 => n68025, A2 => n62233, B1 => n68226, B2 => 
                           n68017, ZN => n7287);
   U47999 : OAI22_X1 port map( A1 => n68025, A2 => n62232, B1 => n68229, B2 => 
                           n68017, ZN => n7288);
   U48000 : OAI22_X1 port map( A1 => n68025, A2 => n62231, B1 => n68232, B2 => 
                           n68017, ZN => n7289);
   U48001 : OAI22_X1 port map( A1 => n68025, A2 => n62230, B1 => n68235, B2 => 
                           n68017, ZN => n7290);
   U48002 : OAI22_X1 port map( A1 => n67995, A2 => n62422, B1 => n68058, B2 => 
                           n67987, ZN => n7103);
   U48003 : OAI22_X1 port map( A1 => n67995, A2 => n62421, B1 => n68061, B2 => 
                           n67987, ZN => n7104);
   U48004 : OAI22_X1 port map( A1 => n67995, A2 => n62420, B1 => n68064, B2 => 
                           n67987, ZN => n7105);
   U48005 : OAI22_X1 port map( A1 => n67995, A2 => n62419, B1 => n68067, B2 => 
                           n67987, ZN => n7106);
   U48006 : OAI22_X1 port map( A1 => n67995, A2 => n62418, B1 => n68070, B2 => 
                           n67987, ZN => n7107);
   U48007 : OAI22_X1 port map( A1 => n67995, A2 => n62417, B1 => n68073, B2 => 
                           n67987, ZN => n7108);
   U48008 : OAI22_X1 port map( A1 => n67995, A2 => n62416, B1 => n68076, B2 => 
                           n67987, ZN => n7109);
   U48009 : OAI22_X1 port map( A1 => n67995, A2 => n62415, B1 => n68079, B2 => 
                           n67987, ZN => n7110);
   U48010 : OAI22_X1 port map( A1 => n67995, A2 => n62414, B1 => n68082, B2 => 
                           n67987, ZN => n7111);
   U48011 : OAI22_X1 port map( A1 => n67995, A2 => n62413, B1 => n68085, B2 => 
                           n67987, ZN => n7112);
   U48012 : OAI22_X1 port map( A1 => n67995, A2 => n62412, B1 => n68088, B2 => 
                           n67987, ZN => n7113);
   U48013 : OAI22_X1 port map( A1 => n67995, A2 => n62411, B1 => n68091, B2 => 
                           n67987, ZN => n7114);
   U48014 : OAI22_X1 port map( A1 => n67996, A2 => n62410, B1 => n68094, B2 => 
                           n67988, ZN => n7115);
   U48015 : OAI22_X1 port map( A1 => n67996, A2 => n62409, B1 => n68097, B2 => 
                           n67988, ZN => n7116);
   U48016 : OAI22_X1 port map( A1 => n67996, A2 => n62408, B1 => n68100, B2 => 
                           n67988, ZN => n7117);
   U48017 : OAI22_X1 port map( A1 => n67996, A2 => n62407, B1 => n68103, B2 => 
                           n67988, ZN => n7118);
   U48018 : OAI22_X1 port map( A1 => n67996, A2 => n62406, B1 => n68106, B2 => 
                           n67988, ZN => n7119);
   U48019 : OAI22_X1 port map( A1 => n67996, A2 => n62405, B1 => n68109, B2 => 
                           n67988, ZN => n7120);
   U48020 : OAI22_X1 port map( A1 => n67996, A2 => n62404, B1 => n68112, B2 => 
                           n67988, ZN => n7121);
   U48021 : OAI22_X1 port map( A1 => n67996, A2 => n62403, B1 => n68115, B2 => 
                           n67988, ZN => n7122);
   U48022 : OAI22_X1 port map( A1 => n67996, A2 => n62402, B1 => n68118, B2 => 
                           n67988, ZN => n7123);
   U48023 : OAI22_X1 port map( A1 => n67996, A2 => n62401, B1 => n68121, B2 => 
                           n67988, ZN => n7124);
   U48024 : OAI22_X1 port map( A1 => n67996, A2 => n62400, B1 => n68124, B2 => 
                           n67988, ZN => n7125);
   U48025 : OAI22_X1 port map( A1 => n67996, A2 => n62399, B1 => n68127, B2 => 
                           n67988, ZN => n7126);
   U48026 : OAI22_X1 port map( A1 => n67996, A2 => n62398, B1 => n68130, B2 => 
                           n67989, ZN => n7127);
   U48027 : OAI22_X1 port map( A1 => n67997, A2 => n62397, B1 => n68133, B2 => 
                           n67989, ZN => n7128);
   U48028 : OAI22_X1 port map( A1 => n67997, A2 => n62396, B1 => n68136, B2 => 
                           n67989, ZN => n7129);
   U48029 : OAI22_X1 port map( A1 => n67997, A2 => n62395, B1 => n68139, B2 => 
                           n67989, ZN => n7130);
   U48030 : OAI22_X1 port map( A1 => n67997, A2 => n62394, B1 => n68142, B2 => 
                           n67989, ZN => n7131);
   U48031 : OAI22_X1 port map( A1 => n67997, A2 => n62393, B1 => n68145, B2 => 
                           n67989, ZN => n7132);
   U48032 : OAI22_X1 port map( A1 => n67997, A2 => n62392, B1 => n68148, B2 => 
                           n67989, ZN => n7133);
   U48033 : OAI22_X1 port map( A1 => n67997, A2 => n62391, B1 => n68151, B2 => 
                           n67989, ZN => n7134);
   U48034 : OAI22_X1 port map( A1 => n67997, A2 => n62390, B1 => n68154, B2 => 
                           n67989, ZN => n7135);
   U48035 : OAI22_X1 port map( A1 => n67997, A2 => n62389, B1 => n68157, B2 => 
                           n67989, ZN => n7136);
   U48036 : OAI22_X1 port map( A1 => n67997, A2 => n62388, B1 => n68160, B2 => 
                           n67989, ZN => n7137);
   U48037 : OAI22_X1 port map( A1 => n67997, A2 => n62387, B1 => n68163, B2 => 
                           n67989, ZN => n7138);
   U48038 : OAI22_X1 port map( A1 => n67997, A2 => n62386, B1 => n68166, B2 => 
                           n67990, ZN => n7139);
   U48039 : OAI22_X1 port map( A1 => n67997, A2 => n62385, B1 => n68169, B2 => 
                           n67990, ZN => n7140);
   U48040 : OAI22_X1 port map( A1 => n67998, A2 => n62384, B1 => n68172, B2 => 
                           n67990, ZN => n7141);
   U48041 : OAI22_X1 port map( A1 => n67998, A2 => n62383, B1 => n68175, B2 => 
                           n67990, ZN => n7142);
   U48042 : OAI22_X1 port map( A1 => n67998, A2 => n62382, B1 => n68178, B2 => 
                           n67990, ZN => n7143);
   U48043 : OAI22_X1 port map( A1 => n67998, A2 => n62381, B1 => n68181, B2 => 
                           n67990, ZN => n7144);
   U48044 : OAI22_X1 port map( A1 => n67998, A2 => n62380, B1 => n68184, B2 => 
                           n67990, ZN => n7145);
   U48045 : OAI22_X1 port map( A1 => n67998, A2 => n62379, B1 => n68187, B2 => 
                           n67990, ZN => n7146);
   U48046 : OAI22_X1 port map( A1 => n67998, A2 => n62378, B1 => n68190, B2 => 
                           n67990, ZN => n7147);
   U48047 : OAI22_X1 port map( A1 => n67998, A2 => n62377, B1 => n68193, B2 => 
                           n67990, ZN => n7148);
   U48048 : OAI22_X1 port map( A1 => n67998, A2 => n62376, B1 => n68196, B2 => 
                           n67990, ZN => n7149);
   U48049 : OAI22_X1 port map( A1 => n67998, A2 => n62375, B1 => n68199, B2 => 
                           n67990, ZN => n7150);
   U48050 : OAI22_X1 port map( A1 => n67998, A2 => n62374, B1 => n68202, B2 => 
                           n67991, ZN => n7151);
   U48051 : OAI22_X1 port map( A1 => n67998, A2 => n62373, B1 => n68205, B2 => 
                           n67991, ZN => n7152);
   U48052 : OAI22_X1 port map( A1 => n67998, A2 => n62372, B1 => n68208, B2 => 
                           n67991, ZN => n7153);
   U48053 : OAI22_X1 port map( A1 => n67999, A2 => n62371, B1 => n68211, B2 => 
                           n67991, ZN => n7154);
   U48054 : OAI22_X1 port map( A1 => n67999, A2 => n62370, B1 => n68214, B2 => 
                           n67991, ZN => n7155);
   U48055 : OAI22_X1 port map( A1 => n67999, A2 => n62369, B1 => n68217, B2 => 
                           n67991, ZN => n7156);
   U48056 : OAI22_X1 port map( A1 => n67999, A2 => n62368, B1 => n68220, B2 => 
                           n67991, ZN => n7157);
   U48057 : OAI22_X1 port map( A1 => n67999, A2 => n62367, B1 => n68223, B2 => 
                           n67991, ZN => n7158);
   U48058 : OAI22_X1 port map( A1 => n67999, A2 => n62366, B1 => n68226, B2 => 
                           n67991, ZN => n7159);
   U48059 : OAI22_X1 port map( A1 => n67999, A2 => n62365, B1 => n68229, B2 => 
                           n67991, ZN => n7160);
   U48060 : OAI22_X1 port map( A1 => n67999, A2 => n62364, B1 => n68232, B2 => 
                           n67991, ZN => n7161);
   U48061 : OAI22_X1 port map( A1 => n67999, A2 => n62363, B1 => n68235, B2 => 
                           n67991, ZN => n7162);
   U48062 : OAI22_X1 port map( A1 => n67816, A2 => n63160, B1 => n68059, B2 => 
                           n67808, ZN => n6207);
   U48063 : OAI22_X1 port map( A1 => n67816, A2 => n63159, B1 => n68062, B2 => 
                           n67808, ZN => n6208);
   U48064 : OAI22_X1 port map( A1 => n67816, A2 => n63158, B1 => n68065, B2 => 
                           n67808, ZN => n6209);
   U48065 : OAI22_X1 port map( A1 => n67816, A2 => n63157, B1 => n68068, B2 => 
                           n67808, ZN => n6210);
   U48066 : OAI22_X1 port map( A1 => n67816, A2 => n63156, B1 => n68071, B2 => 
                           n67808, ZN => n6211);
   U48067 : OAI22_X1 port map( A1 => n67816, A2 => n63155, B1 => n68074, B2 => 
                           n67808, ZN => n6212);
   U48068 : OAI22_X1 port map( A1 => n67816, A2 => n63154, B1 => n68077, B2 => 
                           n67808, ZN => n6213);
   U48069 : OAI22_X1 port map( A1 => n67816, A2 => n63153, B1 => n68080, B2 => 
                           n67808, ZN => n6214);
   U48070 : OAI22_X1 port map( A1 => n67816, A2 => n63152, B1 => n68083, B2 => 
                           n67808, ZN => n6215);
   U48071 : OAI22_X1 port map( A1 => n67816, A2 => n63151, B1 => n68086, B2 => 
                           n67808, ZN => n6216);
   U48072 : OAI22_X1 port map( A1 => n67816, A2 => n63150, B1 => n68089, B2 => 
                           n67808, ZN => n6217);
   U48073 : OAI22_X1 port map( A1 => n67816, A2 => n63149, B1 => n68092, B2 => 
                           n67808, ZN => n6218);
   U48074 : OAI22_X1 port map( A1 => n67817, A2 => n63148, B1 => n68095, B2 => 
                           n67809, ZN => n6219);
   U48075 : OAI22_X1 port map( A1 => n67817, A2 => n63147, B1 => n68098, B2 => 
                           n67809, ZN => n6220);
   U48076 : OAI22_X1 port map( A1 => n67817, A2 => n63146, B1 => n68101, B2 => 
                           n67809, ZN => n6221);
   U48077 : OAI22_X1 port map( A1 => n67817, A2 => n63145, B1 => n68104, B2 => 
                           n67809, ZN => n6222);
   U48078 : OAI22_X1 port map( A1 => n67817, A2 => n63144, B1 => n68107, B2 => 
                           n67809, ZN => n6223);
   U48079 : OAI22_X1 port map( A1 => n67817, A2 => n63143, B1 => n68110, B2 => 
                           n67809, ZN => n6224);
   U48080 : OAI22_X1 port map( A1 => n67817, A2 => n63142, B1 => n68113, B2 => 
                           n67809, ZN => n6225);
   U48081 : OAI22_X1 port map( A1 => n67817, A2 => n63141, B1 => n68116, B2 => 
                           n67809, ZN => n6226);
   U48082 : OAI22_X1 port map( A1 => n67817, A2 => n63140, B1 => n68119, B2 => 
                           n67809, ZN => n6227);
   U48083 : OAI22_X1 port map( A1 => n67817, A2 => n63139, B1 => n68122, B2 => 
                           n67809, ZN => n6228);
   U48084 : OAI22_X1 port map( A1 => n67817, A2 => n63138, B1 => n68125, B2 => 
                           n67809, ZN => n6229);
   U48085 : OAI22_X1 port map( A1 => n67817, A2 => n63137, B1 => n68128, B2 => 
                           n67809, ZN => n6230);
   U48086 : OAI22_X1 port map( A1 => n67817, A2 => n63136, B1 => n68131, B2 => 
                           n67810, ZN => n6231);
   U48087 : OAI22_X1 port map( A1 => n67818, A2 => n63135, B1 => n68134, B2 => 
                           n67810, ZN => n6232);
   U48088 : OAI22_X1 port map( A1 => n67818, A2 => n63134, B1 => n68137, B2 => 
                           n67810, ZN => n6233);
   U48089 : OAI22_X1 port map( A1 => n67818, A2 => n63133, B1 => n68140, B2 => 
                           n67810, ZN => n6234);
   U48090 : OAI22_X1 port map( A1 => n67818, A2 => n63132, B1 => n68143, B2 => 
                           n67810, ZN => n6235);
   U48091 : OAI22_X1 port map( A1 => n67818, A2 => n63131, B1 => n68146, B2 => 
                           n67810, ZN => n6236);
   U48092 : OAI22_X1 port map( A1 => n67818, A2 => n63130, B1 => n68149, B2 => 
                           n67810, ZN => n6237);
   U48093 : OAI22_X1 port map( A1 => n67818, A2 => n63129, B1 => n68152, B2 => 
                           n67810, ZN => n6238);
   U48094 : OAI22_X1 port map( A1 => n67818, A2 => n63128, B1 => n68155, B2 => 
                           n67810, ZN => n6239);
   U48095 : OAI22_X1 port map( A1 => n67818, A2 => n63127, B1 => n68158, B2 => 
                           n67810, ZN => n6240);
   U48096 : OAI22_X1 port map( A1 => n67818, A2 => n63126, B1 => n68161, B2 => 
                           n67810, ZN => n6241);
   U48097 : OAI22_X1 port map( A1 => n67818, A2 => n63125, B1 => n68164, B2 => 
                           n67810, ZN => n6242);
   U48098 : OAI22_X1 port map( A1 => n67818, A2 => n63124, B1 => n68167, B2 => 
                           n67811, ZN => n6243);
   U48099 : OAI22_X1 port map( A1 => n67818, A2 => n63123, B1 => n68170, B2 => 
                           n67811, ZN => n6244);
   U48100 : OAI22_X1 port map( A1 => n67819, A2 => n63122, B1 => n68173, B2 => 
                           n67811, ZN => n6245);
   U48101 : OAI22_X1 port map( A1 => n67819, A2 => n63121, B1 => n68176, B2 => 
                           n67811, ZN => n6246);
   U48102 : OAI22_X1 port map( A1 => n67819, A2 => n63120, B1 => n68179, B2 => 
                           n67811, ZN => n6247);
   U48103 : OAI22_X1 port map( A1 => n67819, A2 => n63119, B1 => n68182, B2 => 
                           n67811, ZN => n6248);
   U48104 : OAI22_X1 port map( A1 => n67819, A2 => n63118, B1 => n68185, B2 => 
                           n67811, ZN => n6249);
   U48105 : OAI22_X1 port map( A1 => n67819, A2 => n63117, B1 => n68188, B2 => 
                           n67811, ZN => n6250);
   U48106 : OAI22_X1 port map( A1 => n67819, A2 => n63116, B1 => n68191, B2 => 
                           n67811, ZN => n6251);
   U48107 : OAI22_X1 port map( A1 => n67819, A2 => n63115, B1 => n68194, B2 => 
                           n67811, ZN => n6252);
   U48108 : OAI22_X1 port map( A1 => n67819, A2 => n63114, B1 => n68197, B2 => 
                           n67811, ZN => n6253);
   U48109 : OAI22_X1 port map( A1 => n67819, A2 => n63113, B1 => n68200, B2 => 
                           n67811, ZN => n6254);
   U48110 : OAI22_X1 port map( A1 => n67819, A2 => n63112, B1 => n68203, B2 => 
                           n67812, ZN => n6255);
   U48111 : OAI22_X1 port map( A1 => n67819, A2 => n63111, B1 => n68206, B2 => 
                           n67812, ZN => n6256);
   U48112 : OAI22_X1 port map( A1 => n67819, A2 => n63110, B1 => n68209, B2 => 
                           n67812, ZN => n6257);
   U48113 : OAI22_X1 port map( A1 => n67820, A2 => n63109, B1 => n68212, B2 => 
                           n67812, ZN => n6258);
   U48114 : OAI22_X1 port map( A1 => n67820, A2 => n63108, B1 => n68215, B2 => 
                           n67812, ZN => n6259);
   U48115 : OAI22_X1 port map( A1 => n67820, A2 => n63107, B1 => n68218, B2 => 
                           n67812, ZN => n6260);
   U48116 : OAI22_X1 port map( A1 => n67820, A2 => n63106, B1 => n68221, B2 => 
                           n67812, ZN => n6261);
   U48117 : OAI22_X1 port map( A1 => n67820, A2 => n63105, B1 => n68224, B2 => 
                           n67812, ZN => n6262);
   U48118 : OAI22_X1 port map( A1 => n67820, A2 => n63104, B1 => n68227, B2 => 
                           n67812, ZN => n6263);
   U48119 : OAI22_X1 port map( A1 => n67820, A2 => n63103, B1 => n68230, B2 => 
                           n67812, ZN => n6264);
   U48120 : OAI22_X1 port map( A1 => n67820, A2 => n63102, B1 => n68233, B2 => 
                           n67812, ZN => n6265);
   U48121 : OAI22_X1 port map( A1 => n67820, A2 => n63101, B1 => n68236, B2 => 
                           n67812, ZN => n6266);
   U48122 : OAI22_X1 port map( A1 => n67982, A2 => n62488, B1 => n68058, B2 => 
                           n67974, ZN => n7039);
   U48123 : OAI22_X1 port map( A1 => n67982, A2 => n62487, B1 => n68061, B2 => 
                           n67974, ZN => n7040);
   U48124 : OAI22_X1 port map( A1 => n67982, A2 => n62486, B1 => n68064, B2 => 
                           n67974, ZN => n7041);
   U48125 : OAI22_X1 port map( A1 => n67982, A2 => n62485, B1 => n68067, B2 => 
                           n67974, ZN => n7042);
   U48126 : OAI22_X1 port map( A1 => n67982, A2 => n62484, B1 => n68070, B2 => 
                           n67974, ZN => n7043);
   U48127 : OAI22_X1 port map( A1 => n67982, A2 => n62483, B1 => n68073, B2 => 
                           n67974, ZN => n7044);
   U48128 : OAI22_X1 port map( A1 => n67982, A2 => n62482, B1 => n68076, B2 => 
                           n67974, ZN => n7045);
   U48129 : OAI22_X1 port map( A1 => n67982, A2 => n62481, B1 => n68079, B2 => 
                           n67974, ZN => n7046);
   U48130 : OAI22_X1 port map( A1 => n67982, A2 => n62480, B1 => n68082, B2 => 
                           n67974, ZN => n7047);
   U48131 : OAI22_X1 port map( A1 => n67982, A2 => n62479, B1 => n68085, B2 => 
                           n67974, ZN => n7048);
   U48132 : OAI22_X1 port map( A1 => n67982, A2 => n62478, B1 => n68088, B2 => 
                           n67974, ZN => n7049);
   U48133 : OAI22_X1 port map( A1 => n67982, A2 => n62477, B1 => n68091, B2 => 
                           n67974, ZN => n7050);
   U48134 : OAI22_X1 port map( A1 => n67983, A2 => n62476, B1 => n68094, B2 => 
                           n67975, ZN => n7051);
   U48135 : OAI22_X1 port map( A1 => n67983, A2 => n62475, B1 => n68097, B2 => 
                           n67975, ZN => n7052);
   U48136 : OAI22_X1 port map( A1 => n67983, A2 => n62474, B1 => n68100, B2 => 
                           n67975, ZN => n7053);
   U48137 : OAI22_X1 port map( A1 => n67983, A2 => n62473, B1 => n68103, B2 => 
                           n67975, ZN => n7054);
   U48138 : OAI22_X1 port map( A1 => n67983, A2 => n62472, B1 => n68106, B2 => 
                           n67975, ZN => n7055);
   U48139 : OAI22_X1 port map( A1 => n67983, A2 => n62471, B1 => n68109, B2 => 
                           n67975, ZN => n7056);
   U48140 : OAI22_X1 port map( A1 => n67983, A2 => n62470, B1 => n68112, B2 => 
                           n67975, ZN => n7057);
   U48141 : OAI22_X1 port map( A1 => n67983, A2 => n62469, B1 => n68115, B2 => 
                           n67975, ZN => n7058);
   U48142 : OAI22_X1 port map( A1 => n67983, A2 => n62468, B1 => n68118, B2 => 
                           n67975, ZN => n7059);
   U48143 : OAI22_X1 port map( A1 => n67983, A2 => n62467, B1 => n68121, B2 => 
                           n67975, ZN => n7060);
   U48144 : OAI22_X1 port map( A1 => n67983, A2 => n62466, B1 => n68124, B2 => 
                           n67975, ZN => n7061);
   U48145 : OAI22_X1 port map( A1 => n67983, A2 => n62465, B1 => n68127, B2 => 
                           n67975, ZN => n7062);
   U48146 : OAI22_X1 port map( A1 => n67983, A2 => n62464, B1 => n68130, B2 => 
                           n67976, ZN => n7063);
   U48147 : OAI22_X1 port map( A1 => n67984, A2 => n62463, B1 => n68133, B2 => 
                           n67976, ZN => n7064);
   U48148 : OAI22_X1 port map( A1 => n67984, A2 => n62462, B1 => n68136, B2 => 
                           n67976, ZN => n7065);
   U48149 : OAI22_X1 port map( A1 => n67984, A2 => n62461, B1 => n68139, B2 => 
                           n67976, ZN => n7066);
   U48150 : OAI22_X1 port map( A1 => n67984, A2 => n62460, B1 => n68142, B2 => 
                           n67976, ZN => n7067);
   U48151 : OAI22_X1 port map( A1 => n67984, A2 => n62459, B1 => n68145, B2 => 
                           n67976, ZN => n7068);
   U48152 : OAI22_X1 port map( A1 => n67984, A2 => n62458, B1 => n68148, B2 => 
                           n67976, ZN => n7069);
   U48153 : OAI22_X1 port map( A1 => n67984, A2 => n62457, B1 => n68151, B2 => 
                           n67976, ZN => n7070);
   U48154 : OAI22_X1 port map( A1 => n67984, A2 => n62456, B1 => n68154, B2 => 
                           n67976, ZN => n7071);
   U48155 : OAI22_X1 port map( A1 => n67984, A2 => n62455, B1 => n68157, B2 => 
                           n67976, ZN => n7072);
   U48156 : OAI22_X1 port map( A1 => n67984, A2 => n62454, B1 => n68160, B2 => 
                           n67976, ZN => n7073);
   U48157 : OAI22_X1 port map( A1 => n67984, A2 => n62453, B1 => n68163, B2 => 
                           n67976, ZN => n7074);
   U48158 : OAI22_X1 port map( A1 => n67984, A2 => n62452, B1 => n68166, B2 => 
                           n67977, ZN => n7075);
   U48159 : OAI22_X1 port map( A1 => n67984, A2 => n62451, B1 => n68169, B2 => 
                           n67977, ZN => n7076);
   U48160 : OAI22_X1 port map( A1 => n67985, A2 => n62450, B1 => n68172, B2 => 
                           n67977, ZN => n7077);
   U48161 : OAI22_X1 port map( A1 => n67985, A2 => n62449, B1 => n68175, B2 => 
                           n67977, ZN => n7078);
   U48162 : OAI22_X1 port map( A1 => n67985, A2 => n62448, B1 => n68178, B2 => 
                           n67977, ZN => n7079);
   U48163 : OAI22_X1 port map( A1 => n67985, A2 => n62447, B1 => n68181, B2 => 
                           n67977, ZN => n7080);
   U48164 : OAI22_X1 port map( A1 => n67985, A2 => n62446, B1 => n68184, B2 => 
                           n67977, ZN => n7081);
   U48165 : OAI22_X1 port map( A1 => n67985, A2 => n62445, B1 => n68187, B2 => 
                           n67977, ZN => n7082);
   U48166 : OAI22_X1 port map( A1 => n67985, A2 => n62444, B1 => n68190, B2 => 
                           n67977, ZN => n7083);
   U48167 : OAI22_X1 port map( A1 => n67985, A2 => n62443, B1 => n68193, B2 => 
                           n67977, ZN => n7084);
   U48168 : OAI22_X1 port map( A1 => n67985, A2 => n62442, B1 => n68196, B2 => 
                           n67977, ZN => n7085);
   U48169 : OAI22_X1 port map( A1 => n67985, A2 => n62441, B1 => n68199, B2 => 
                           n67977, ZN => n7086);
   U48170 : OAI22_X1 port map( A1 => n67985, A2 => n62440, B1 => n68202, B2 => 
                           n67978, ZN => n7087);
   U48171 : OAI22_X1 port map( A1 => n67985, A2 => n62439, B1 => n68205, B2 => 
                           n67978, ZN => n7088);
   U48172 : OAI22_X1 port map( A1 => n67985, A2 => n62438, B1 => n68208, B2 => 
                           n67978, ZN => n7089);
   U48173 : OAI22_X1 port map( A1 => n67986, A2 => n62437, B1 => n68211, B2 => 
                           n67978, ZN => n7090);
   U48174 : OAI22_X1 port map( A1 => n67986, A2 => n62436, B1 => n68214, B2 => 
                           n67978, ZN => n7091);
   U48175 : OAI22_X1 port map( A1 => n67986, A2 => n62435, B1 => n68217, B2 => 
                           n67978, ZN => n7092);
   U48176 : OAI22_X1 port map( A1 => n67986, A2 => n62434, B1 => n68220, B2 => 
                           n67978, ZN => n7093);
   U48177 : OAI22_X1 port map( A1 => n67986, A2 => n62433, B1 => n68223, B2 => 
                           n67978, ZN => n7094);
   U48178 : OAI22_X1 port map( A1 => n67986, A2 => n62432, B1 => n68226, B2 => 
                           n67978, ZN => n7095);
   U48179 : OAI22_X1 port map( A1 => n67986, A2 => n62431, B1 => n68229, B2 => 
                           n67978, ZN => n7096);
   U48180 : OAI22_X1 port map( A1 => n67986, A2 => n62430, B1 => n68232, B2 => 
                           n67978, ZN => n7097);
   U48181 : OAI22_X1 port map( A1 => n67986, A2 => n62429, B1 => n68235, B2 => 
                           n67978, ZN => n7098);
   U48182 : OAI22_X1 port map( A1 => n67765, A2 => n63361, B1 => n68059, B2 => 
                           n67757, ZN => n5951);
   U48183 : OAI22_X1 port map( A1 => n67765, A2 => n63360, B1 => n68062, B2 => 
                           n67757, ZN => n5952);
   U48184 : OAI22_X1 port map( A1 => n67765, A2 => n63359, B1 => n68065, B2 => 
                           n67757, ZN => n5953);
   U48185 : OAI22_X1 port map( A1 => n67765, A2 => n63358, B1 => n68068, B2 => 
                           n67757, ZN => n5954);
   U48186 : OAI22_X1 port map( A1 => n67765, A2 => n63357, B1 => n68071, B2 => 
                           n67757, ZN => n5955);
   U48187 : OAI22_X1 port map( A1 => n67765, A2 => n63356, B1 => n68074, B2 => 
                           n67757, ZN => n5956);
   U48188 : OAI22_X1 port map( A1 => n67765, A2 => n63355, B1 => n68077, B2 => 
                           n67757, ZN => n5957);
   U48189 : OAI22_X1 port map( A1 => n67765, A2 => n63354, B1 => n68080, B2 => 
                           n67757, ZN => n5958);
   U48190 : OAI22_X1 port map( A1 => n67765, A2 => n63353, B1 => n68083, B2 => 
                           n67757, ZN => n5959);
   U48191 : OAI22_X1 port map( A1 => n67765, A2 => n63352, B1 => n68086, B2 => 
                           n67757, ZN => n5960);
   U48192 : OAI22_X1 port map( A1 => n67765, A2 => n63351, B1 => n68089, B2 => 
                           n67757, ZN => n5961);
   U48193 : OAI22_X1 port map( A1 => n67765, A2 => n63350, B1 => n68092, B2 => 
                           n67757, ZN => n5962);
   U48194 : OAI22_X1 port map( A1 => n67766, A2 => n63349, B1 => n68095, B2 => 
                           n67758, ZN => n5963);
   U48195 : OAI22_X1 port map( A1 => n67766, A2 => n63348, B1 => n68098, B2 => 
                           n67758, ZN => n5964);
   U48196 : OAI22_X1 port map( A1 => n67766, A2 => n63347, B1 => n68101, B2 => 
                           n67758, ZN => n5965);
   U48197 : OAI22_X1 port map( A1 => n67766, A2 => n63346, B1 => n68104, B2 => 
                           n67758, ZN => n5966);
   U48198 : OAI22_X1 port map( A1 => n67766, A2 => n63345, B1 => n68107, B2 => 
                           n67758, ZN => n5967);
   U48199 : OAI22_X1 port map( A1 => n67766, A2 => n63344, B1 => n68110, B2 => 
                           n67758, ZN => n5968);
   U48200 : OAI22_X1 port map( A1 => n67766, A2 => n63343, B1 => n68113, B2 => 
                           n67758, ZN => n5969);
   U48201 : OAI22_X1 port map( A1 => n67766, A2 => n63342, B1 => n68116, B2 => 
                           n67758, ZN => n5970);
   U48202 : OAI22_X1 port map( A1 => n67766, A2 => n63341, B1 => n68119, B2 => 
                           n67758, ZN => n5971);
   U48203 : OAI22_X1 port map( A1 => n67766, A2 => n63340, B1 => n68122, B2 => 
                           n67758, ZN => n5972);
   U48204 : OAI22_X1 port map( A1 => n67766, A2 => n63339, B1 => n68125, B2 => 
                           n67758, ZN => n5973);
   U48205 : OAI22_X1 port map( A1 => n67766, A2 => n63338, B1 => n68128, B2 => 
                           n67758, ZN => n5974);
   U48206 : OAI22_X1 port map( A1 => n67766, A2 => n63337, B1 => n68131, B2 => 
                           n67759, ZN => n5975);
   U48207 : OAI22_X1 port map( A1 => n67767, A2 => n63336, B1 => n68134, B2 => 
                           n67759, ZN => n5976);
   U48208 : OAI22_X1 port map( A1 => n67767, A2 => n63335, B1 => n68137, B2 => 
                           n67759, ZN => n5977);
   U48209 : OAI22_X1 port map( A1 => n67767, A2 => n63334, B1 => n68140, B2 => 
                           n67759, ZN => n5978);
   U48210 : OAI22_X1 port map( A1 => n67767, A2 => n63333, B1 => n68143, B2 => 
                           n67759, ZN => n5979);
   U48211 : OAI22_X1 port map( A1 => n67767, A2 => n63332, B1 => n68146, B2 => 
                           n67759, ZN => n5980);
   U48212 : OAI22_X1 port map( A1 => n67767, A2 => n63331, B1 => n68149, B2 => 
                           n67759, ZN => n5981);
   U48213 : OAI22_X1 port map( A1 => n67767, A2 => n63330, B1 => n68152, B2 => 
                           n67759, ZN => n5982);
   U48214 : OAI22_X1 port map( A1 => n67767, A2 => n63329, B1 => n68155, B2 => 
                           n67759, ZN => n5983);
   U48215 : OAI22_X1 port map( A1 => n67767, A2 => n63328, B1 => n68158, B2 => 
                           n67759, ZN => n5984);
   U48216 : OAI22_X1 port map( A1 => n67767, A2 => n63327, B1 => n68161, B2 => 
                           n67759, ZN => n5985);
   U48217 : OAI22_X1 port map( A1 => n67767, A2 => n63326, B1 => n68164, B2 => 
                           n67759, ZN => n5986);
   U48218 : OAI22_X1 port map( A1 => n67767, A2 => n63325, B1 => n68167, B2 => 
                           n67760, ZN => n5987);
   U48219 : OAI22_X1 port map( A1 => n67767, A2 => n63324, B1 => n68170, B2 => 
                           n67760, ZN => n5988);
   U48220 : OAI22_X1 port map( A1 => n67768, A2 => n63323, B1 => n68173, B2 => 
                           n67760, ZN => n5989);
   U48221 : OAI22_X1 port map( A1 => n67768, A2 => n63322, B1 => n68176, B2 => 
                           n67760, ZN => n5990);
   U48222 : OAI22_X1 port map( A1 => n67768, A2 => n63321, B1 => n68179, B2 => 
                           n67760, ZN => n5991);
   U48223 : OAI22_X1 port map( A1 => n67768, A2 => n63320, B1 => n68182, B2 => 
                           n67760, ZN => n5992);
   U48224 : OAI22_X1 port map( A1 => n67768, A2 => n63319, B1 => n68185, B2 => 
                           n67760, ZN => n5993);
   U48225 : OAI22_X1 port map( A1 => n67768, A2 => n63318, B1 => n68188, B2 => 
                           n67760, ZN => n5994);
   U48226 : OAI22_X1 port map( A1 => n67768, A2 => n63317, B1 => n68191, B2 => 
                           n67760, ZN => n5995);
   U48227 : OAI22_X1 port map( A1 => n67768, A2 => n63316, B1 => n68194, B2 => 
                           n67760, ZN => n5996);
   U48228 : OAI22_X1 port map( A1 => n67768, A2 => n63315, B1 => n68197, B2 => 
                           n67760, ZN => n5997);
   U48229 : OAI22_X1 port map( A1 => n67768, A2 => n63314, B1 => n68200, B2 => 
                           n67760, ZN => n5998);
   U48230 : OAI22_X1 port map( A1 => n67768, A2 => n63313, B1 => n68203, B2 => 
                           n67761, ZN => n5999);
   U48231 : OAI22_X1 port map( A1 => n67768, A2 => n63312, B1 => n68206, B2 => 
                           n67761, ZN => n6000);
   U48232 : OAI22_X1 port map( A1 => n67768, A2 => n63311, B1 => n68209, B2 => 
                           n67761, ZN => n6001);
   U48233 : OAI22_X1 port map( A1 => n67769, A2 => n63310, B1 => n68212, B2 => 
                           n67761, ZN => n6002);
   U48234 : OAI22_X1 port map( A1 => n67769, A2 => n63309, B1 => n68215, B2 => 
                           n67761, ZN => n6003);
   U48235 : OAI22_X1 port map( A1 => n67769, A2 => n63308, B1 => n68218, B2 => 
                           n67761, ZN => n6004);
   U48236 : OAI22_X1 port map( A1 => n67769, A2 => n63307, B1 => n68221, B2 => 
                           n67761, ZN => n6005);
   U48237 : OAI22_X1 port map( A1 => n67769, A2 => n63306, B1 => n68224, B2 => 
                           n67761, ZN => n6006);
   U48238 : OAI22_X1 port map( A1 => n67769, A2 => n63305, B1 => n68227, B2 => 
                           n67761, ZN => n6007);
   U48239 : OAI22_X1 port map( A1 => n67769, A2 => n63304, B1 => n68230, B2 => 
                           n67761, ZN => n6008);
   U48240 : OAI22_X1 port map( A1 => n67769, A2 => n63303, B1 => n68233, B2 => 
                           n67761, ZN => n6009);
   U48241 : OAI22_X1 port map( A1 => n67769, A2 => n63302, B1 => n68236, B2 => 
                           n67761, ZN => n6010);
   U48242 : OAI22_X1 port map( A1 => n67867, A2 => n62957, B1 => n68059, B2 => 
                           n67859, ZN => n6463);
   U48243 : OAI22_X1 port map( A1 => n67867, A2 => n62956, B1 => n68062, B2 => 
                           n67859, ZN => n6464);
   U48244 : OAI22_X1 port map( A1 => n67867, A2 => n62955, B1 => n68065, B2 => 
                           n67859, ZN => n6465);
   U48245 : OAI22_X1 port map( A1 => n67867, A2 => n62954, B1 => n68068, B2 => 
                           n67859, ZN => n6466);
   U48246 : OAI22_X1 port map( A1 => n67867, A2 => n62953, B1 => n68071, B2 => 
                           n67859, ZN => n6467);
   U48247 : OAI22_X1 port map( A1 => n67867, A2 => n62952, B1 => n68074, B2 => 
                           n67859, ZN => n6468);
   U48248 : OAI22_X1 port map( A1 => n67867, A2 => n62951, B1 => n68077, B2 => 
                           n67859, ZN => n6469);
   U48249 : OAI22_X1 port map( A1 => n67867, A2 => n62950, B1 => n68080, B2 => 
                           n67859, ZN => n6470);
   U48250 : OAI22_X1 port map( A1 => n67867, A2 => n62949, B1 => n68083, B2 => 
                           n67859, ZN => n6471);
   U48251 : OAI22_X1 port map( A1 => n67867, A2 => n62948, B1 => n68086, B2 => 
                           n67859, ZN => n6472);
   U48252 : OAI22_X1 port map( A1 => n67867, A2 => n62947, B1 => n68089, B2 => 
                           n67859, ZN => n6473);
   U48253 : OAI22_X1 port map( A1 => n67867, A2 => n62946, B1 => n68092, B2 => 
                           n67859, ZN => n6474);
   U48254 : OAI22_X1 port map( A1 => n67868, A2 => n62945, B1 => n68095, B2 => 
                           n67860, ZN => n6475);
   U48255 : OAI22_X1 port map( A1 => n67868, A2 => n62944, B1 => n68098, B2 => 
                           n67860, ZN => n6476);
   U48256 : OAI22_X1 port map( A1 => n67868, A2 => n62943, B1 => n68101, B2 => 
                           n67860, ZN => n6477);
   U48257 : OAI22_X1 port map( A1 => n67868, A2 => n62942, B1 => n68104, B2 => 
                           n67860, ZN => n6478);
   U48258 : OAI22_X1 port map( A1 => n67868, A2 => n62941, B1 => n68107, B2 => 
                           n67860, ZN => n6479);
   U48259 : OAI22_X1 port map( A1 => n67868, A2 => n62940, B1 => n68110, B2 => 
                           n67860, ZN => n6480);
   U48260 : OAI22_X1 port map( A1 => n67868, A2 => n62939, B1 => n68113, B2 => 
                           n67860, ZN => n6481);
   U48261 : OAI22_X1 port map( A1 => n67868, A2 => n62938, B1 => n68116, B2 => 
                           n67860, ZN => n6482);
   U48262 : OAI22_X1 port map( A1 => n67868, A2 => n62937, B1 => n68119, B2 => 
                           n67860, ZN => n6483);
   U48263 : OAI22_X1 port map( A1 => n67868, A2 => n62936, B1 => n68122, B2 => 
                           n67860, ZN => n6484);
   U48264 : OAI22_X1 port map( A1 => n67868, A2 => n62935, B1 => n68125, B2 => 
                           n67860, ZN => n6485);
   U48265 : OAI22_X1 port map( A1 => n67868, A2 => n62934, B1 => n68128, B2 => 
                           n67860, ZN => n6486);
   U48266 : OAI22_X1 port map( A1 => n67868, A2 => n62933, B1 => n68131, B2 => 
                           n67861, ZN => n6487);
   U48267 : OAI22_X1 port map( A1 => n67869, A2 => n62932, B1 => n68134, B2 => 
                           n67861, ZN => n6488);
   U48268 : OAI22_X1 port map( A1 => n67869, A2 => n62931, B1 => n68137, B2 => 
                           n67861, ZN => n6489);
   U48269 : OAI22_X1 port map( A1 => n67869, A2 => n62930, B1 => n68140, B2 => 
                           n67861, ZN => n6490);
   U48270 : OAI22_X1 port map( A1 => n67869, A2 => n62929, B1 => n68143, B2 => 
                           n67861, ZN => n6491);
   U48271 : OAI22_X1 port map( A1 => n67869, A2 => n62928, B1 => n68146, B2 => 
                           n67861, ZN => n6492);
   U48272 : OAI22_X1 port map( A1 => n67869, A2 => n62927, B1 => n68149, B2 => 
                           n67861, ZN => n6493);
   U48273 : OAI22_X1 port map( A1 => n67869, A2 => n62926, B1 => n68152, B2 => 
                           n67861, ZN => n6494);
   U48274 : OAI22_X1 port map( A1 => n67869, A2 => n62925, B1 => n68155, B2 => 
                           n67861, ZN => n6495);
   U48275 : OAI22_X1 port map( A1 => n67869, A2 => n62924, B1 => n68158, B2 => 
                           n67861, ZN => n6496);
   U48276 : OAI22_X1 port map( A1 => n67869, A2 => n62923, B1 => n68161, B2 => 
                           n67861, ZN => n6497);
   U48277 : OAI22_X1 port map( A1 => n67869, A2 => n62922, B1 => n68164, B2 => 
                           n67861, ZN => n6498);
   U48278 : OAI22_X1 port map( A1 => n67869, A2 => n62921, B1 => n68167, B2 => 
                           n67862, ZN => n6499);
   U48279 : OAI22_X1 port map( A1 => n67869, A2 => n62920, B1 => n68170, B2 => 
                           n67862, ZN => n6500);
   U48280 : OAI22_X1 port map( A1 => n67870, A2 => n62919, B1 => n68173, B2 => 
                           n67862, ZN => n6501);
   U48281 : OAI22_X1 port map( A1 => n67870, A2 => n62918, B1 => n68176, B2 => 
                           n67862, ZN => n6502);
   U48282 : OAI22_X1 port map( A1 => n67870, A2 => n62917, B1 => n68179, B2 => 
                           n67862, ZN => n6503);
   U48283 : OAI22_X1 port map( A1 => n67870, A2 => n62916, B1 => n68182, B2 => 
                           n67862, ZN => n6504);
   U48284 : OAI22_X1 port map( A1 => n67870, A2 => n62915, B1 => n68185, B2 => 
                           n67862, ZN => n6505);
   U48285 : OAI22_X1 port map( A1 => n67870, A2 => n62914, B1 => n68188, B2 => 
                           n67862, ZN => n6506);
   U48286 : OAI22_X1 port map( A1 => n67870, A2 => n62913, B1 => n68191, B2 => 
                           n67862, ZN => n6507);
   U48287 : OAI22_X1 port map( A1 => n67870, A2 => n62912, B1 => n68194, B2 => 
                           n67862, ZN => n6508);
   U48288 : OAI22_X1 port map( A1 => n67870, A2 => n62911, B1 => n68197, B2 => 
                           n67862, ZN => n6509);
   U48289 : OAI22_X1 port map( A1 => n67870, A2 => n62910, B1 => n68200, B2 => 
                           n67862, ZN => n6510);
   U48290 : OAI22_X1 port map( A1 => n67870, A2 => n62909, B1 => n68203, B2 => 
                           n67863, ZN => n6511);
   U48291 : OAI22_X1 port map( A1 => n67870, A2 => n62908, B1 => n68206, B2 => 
                           n67863, ZN => n6512);
   U48292 : OAI22_X1 port map( A1 => n67870, A2 => n62907, B1 => n68209, B2 => 
                           n67863, ZN => n6513);
   U48293 : OAI22_X1 port map( A1 => n67871, A2 => n62906, B1 => n68212, B2 => 
                           n67863, ZN => n6514);
   U48294 : OAI22_X1 port map( A1 => n67871, A2 => n62905, B1 => n68215, B2 => 
                           n67863, ZN => n6515);
   U48295 : OAI22_X1 port map( A1 => n67871, A2 => n62904, B1 => n68218, B2 => 
                           n67863, ZN => n6516);
   U48296 : OAI22_X1 port map( A1 => n67871, A2 => n62903, B1 => n68221, B2 => 
                           n67863, ZN => n6517);
   U48297 : OAI22_X1 port map( A1 => n67871, A2 => n62902, B1 => n68224, B2 => 
                           n67863, ZN => n6518);
   U48298 : OAI22_X1 port map( A1 => n67871, A2 => n62901, B1 => n68227, B2 => 
                           n67863, ZN => n6519);
   U48299 : OAI22_X1 port map( A1 => n67871, A2 => n62900, B1 => n68230, B2 => 
                           n67863, ZN => n6520);
   U48300 : OAI22_X1 port map( A1 => n67871, A2 => n62899, B1 => n68233, B2 => 
                           n67863, ZN => n6521);
   U48301 : OAI22_X1 port map( A1 => n67871, A2 => n62898, B1 => n68236, B2 => 
                           n67863, ZN => n6522);
   U48302 : OAI22_X1 port map( A1 => n67918, A2 => n62761, B1 => n68058, B2 => 
                           n67910, ZN => n6719);
   U48303 : OAI22_X1 port map( A1 => n67918, A2 => n62760, B1 => n68061, B2 => 
                           n67910, ZN => n6720);
   U48304 : OAI22_X1 port map( A1 => n67918, A2 => n62759, B1 => n68064, B2 => 
                           n67910, ZN => n6721);
   U48305 : OAI22_X1 port map( A1 => n67918, A2 => n62758, B1 => n68067, B2 => 
                           n67910, ZN => n6722);
   U48306 : OAI22_X1 port map( A1 => n67918, A2 => n62757, B1 => n68070, B2 => 
                           n67910, ZN => n6723);
   U48307 : OAI22_X1 port map( A1 => n67918, A2 => n62756, B1 => n68073, B2 => 
                           n67910, ZN => n6724);
   U48308 : OAI22_X1 port map( A1 => n67918, A2 => n62755, B1 => n68076, B2 => 
                           n67910, ZN => n6725);
   U48309 : OAI22_X1 port map( A1 => n67918, A2 => n62754, B1 => n68079, B2 => 
                           n67910, ZN => n6726);
   U48310 : OAI22_X1 port map( A1 => n67918, A2 => n62753, B1 => n68082, B2 => 
                           n67910, ZN => n6727);
   U48311 : OAI22_X1 port map( A1 => n67918, A2 => n62752, B1 => n68085, B2 => 
                           n67910, ZN => n6728);
   U48312 : OAI22_X1 port map( A1 => n67918, A2 => n62751, B1 => n68088, B2 => 
                           n67910, ZN => n6729);
   U48313 : OAI22_X1 port map( A1 => n67918, A2 => n62750, B1 => n68091, B2 => 
                           n67910, ZN => n6730);
   U48314 : OAI22_X1 port map( A1 => n67919, A2 => n62749, B1 => n68094, B2 => 
                           n67911, ZN => n6731);
   U48315 : OAI22_X1 port map( A1 => n67919, A2 => n62748, B1 => n68097, B2 => 
                           n67911, ZN => n6732);
   U48316 : OAI22_X1 port map( A1 => n67919, A2 => n62747, B1 => n68100, B2 => 
                           n67911, ZN => n6733);
   U48317 : OAI22_X1 port map( A1 => n67919, A2 => n62746, B1 => n68103, B2 => 
                           n67911, ZN => n6734);
   U48318 : OAI22_X1 port map( A1 => n67919, A2 => n62745, B1 => n68106, B2 => 
                           n67911, ZN => n6735);
   U48319 : OAI22_X1 port map( A1 => n67919, A2 => n62744, B1 => n68109, B2 => 
                           n67911, ZN => n6736);
   U48320 : OAI22_X1 port map( A1 => n67919, A2 => n62743, B1 => n68112, B2 => 
                           n67911, ZN => n6737);
   U48321 : OAI22_X1 port map( A1 => n67919, A2 => n62742, B1 => n68115, B2 => 
                           n67911, ZN => n6738);
   U48322 : OAI22_X1 port map( A1 => n67919, A2 => n62741, B1 => n68118, B2 => 
                           n67911, ZN => n6739);
   U48323 : OAI22_X1 port map( A1 => n67919, A2 => n62740, B1 => n68121, B2 => 
                           n67911, ZN => n6740);
   U48324 : OAI22_X1 port map( A1 => n67919, A2 => n62739, B1 => n68124, B2 => 
                           n67911, ZN => n6741);
   U48325 : OAI22_X1 port map( A1 => n67919, A2 => n62738, B1 => n68127, B2 => 
                           n67911, ZN => n6742);
   U48326 : OAI22_X1 port map( A1 => n67919, A2 => n62737, B1 => n68130, B2 => 
                           n67912, ZN => n6743);
   U48327 : OAI22_X1 port map( A1 => n67920, A2 => n62736, B1 => n68133, B2 => 
                           n67912, ZN => n6744);
   U48328 : OAI22_X1 port map( A1 => n67920, A2 => n62735, B1 => n68136, B2 => 
                           n67912, ZN => n6745);
   U48329 : OAI22_X1 port map( A1 => n67920, A2 => n62734, B1 => n68139, B2 => 
                           n67912, ZN => n6746);
   U48330 : OAI22_X1 port map( A1 => n67920, A2 => n62733, B1 => n68142, B2 => 
                           n67912, ZN => n6747);
   U48331 : OAI22_X1 port map( A1 => n67920, A2 => n62732, B1 => n68145, B2 => 
                           n67912, ZN => n6748);
   U48332 : OAI22_X1 port map( A1 => n67920, A2 => n62731, B1 => n68148, B2 => 
                           n67912, ZN => n6749);
   U48333 : OAI22_X1 port map( A1 => n67920, A2 => n62730, B1 => n68151, B2 => 
                           n67912, ZN => n6750);
   U48334 : OAI22_X1 port map( A1 => n67920, A2 => n62729, B1 => n68154, B2 => 
                           n67912, ZN => n6751);
   U48335 : OAI22_X1 port map( A1 => n67920, A2 => n62728, B1 => n68157, B2 => 
                           n67912, ZN => n6752);
   U48336 : OAI22_X1 port map( A1 => n67920, A2 => n62727, B1 => n68160, B2 => 
                           n67912, ZN => n6753);
   U48337 : OAI22_X1 port map( A1 => n67920, A2 => n62726, B1 => n68163, B2 => 
                           n67912, ZN => n6754);
   U48338 : OAI22_X1 port map( A1 => n67920, A2 => n62725, B1 => n68166, B2 => 
                           n67913, ZN => n6755);
   U48339 : OAI22_X1 port map( A1 => n67920, A2 => n62724, B1 => n68169, B2 => 
                           n67913, ZN => n6756);
   U48340 : OAI22_X1 port map( A1 => n67921, A2 => n62723, B1 => n68172, B2 => 
                           n67913, ZN => n6757);
   U48341 : OAI22_X1 port map( A1 => n67921, A2 => n62722, B1 => n68175, B2 => 
                           n67913, ZN => n6758);
   U48342 : OAI22_X1 port map( A1 => n67921, A2 => n62721, B1 => n68178, B2 => 
                           n67913, ZN => n6759);
   U48343 : OAI22_X1 port map( A1 => n67921, A2 => n62720, B1 => n68181, B2 => 
                           n67913, ZN => n6760);
   U48344 : OAI22_X1 port map( A1 => n67921, A2 => n62719, B1 => n68184, B2 => 
                           n67913, ZN => n6761);
   U48345 : OAI22_X1 port map( A1 => n67921, A2 => n62718, B1 => n68187, B2 => 
                           n67913, ZN => n6762);
   U48346 : OAI22_X1 port map( A1 => n67921, A2 => n62717, B1 => n68190, B2 => 
                           n67913, ZN => n6763);
   U48347 : OAI22_X1 port map( A1 => n67921, A2 => n62716, B1 => n68193, B2 => 
                           n67913, ZN => n6764);
   U48348 : OAI22_X1 port map( A1 => n67921, A2 => n62715, B1 => n68196, B2 => 
                           n67913, ZN => n6765);
   U48349 : OAI22_X1 port map( A1 => n67921, A2 => n62714, B1 => n68199, B2 => 
                           n67913, ZN => n6766);
   U48350 : OAI22_X1 port map( A1 => n67921, A2 => n62713, B1 => n68202, B2 => 
                           n67914, ZN => n6767);
   U48351 : OAI22_X1 port map( A1 => n67921, A2 => n62712, B1 => n68205, B2 => 
                           n67914, ZN => n6768);
   U48352 : OAI22_X1 port map( A1 => n67921, A2 => n62711, B1 => n68208, B2 => 
                           n67914, ZN => n6769);
   U48353 : OAI22_X1 port map( A1 => n67922, A2 => n62710, B1 => n68211, B2 => 
                           n67914, ZN => n6770);
   U48354 : OAI22_X1 port map( A1 => n67922, A2 => n62709, B1 => n68214, B2 => 
                           n67914, ZN => n6771);
   U48355 : OAI22_X1 port map( A1 => n67922, A2 => n62708, B1 => n68217, B2 => 
                           n67914, ZN => n6772);
   U48356 : OAI22_X1 port map( A1 => n67922, A2 => n62707, B1 => n68220, B2 => 
                           n67914, ZN => n6773);
   U48357 : OAI22_X1 port map( A1 => n67922, A2 => n62706, B1 => n68223, B2 => 
                           n67914, ZN => n6774);
   U48358 : OAI22_X1 port map( A1 => n67922, A2 => n62705, B1 => n68226, B2 => 
                           n67914, ZN => n6775);
   U48359 : OAI22_X1 port map( A1 => n67922, A2 => n62704, B1 => n68229, B2 => 
                           n67914, ZN => n6776);
   U48360 : OAI22_X1 port map( A1 => n67922, A2 => n62703, B1 => n68232, B2 => 
                           n67914, ZN => n6777);
   U48361 : OAI22_X1 port map( A1 => n67922, A2 => n62702, B1 => n68235, B2 => 
                           n67914, ZN => n6778);
   U48362 : NAND2_X1 port map( A1 => n65076, A2 => n65086, ZN => n63807);
   U48363 : OAI21_X1 port map( B1 => n62156, B2 => n62489, A => n68052, ZN => 
                           n62493);
   U48364 : OAI21_X1 port map( B1 => n62156, B2 => n62223, A => n68052, ZN => 
                           n62224);
   U48365 : OAI21_X1 port map( B1 => n62156, B2 => n62356, A => n68052, ZN => 
                           n62357);
   U48366 : OAI21_X1 port map( B1 => n62088, B2 => n62356, A => n68052, ZN => 
                           n62290);
   U48367 : OAI21_X1 port map( B1 => n62088, B2 => n62223, A => n68052, ZN => 
                           n62157);
   U48368 : OAI21_X1 port map( B1 => n62088, B2 => n62489, A => n68052, ZN => 
                           n62423);
   U48369 : NAND2_X1 port map( A1 => n65087, A2 => n65074, ZN => n63785);
   U48370 : BUF_X1 port map( A => n62086, Z => n68060);
   U48371 : BUF_X1 port map( A => n62084, Z => n68063);
   U48372 : BUF_X1 port map( A => n62082, Z => n68066);
   U48373 : BUF_X1 port map( A => n62080, Z => n68069);
   U48374 : BUF_X1 port map( A => n62078, Z => n68072);
   U48375 : BUF_X1 port map( A => n62076, Z => n68075);
   U48376 : BUF_X1 port map( A => n62074, Z => n68078);
   U48377 : BUF_X1 port map( A => n62072, Z => n68081);
   U48378 : BUF_X1 port map( A => n62070, Z => n68084);
   U48379 : BUF_X1 port map( A => n62068, Z => n68087);
   U48380 : BUF_X1 port map( A => n62066, Z => n68090);
   U48381 : BUF_X1 port map( A => n62064, Z => n68093);
   U48382 : BUF_X1 port map( A => n62062, Z => n68096);
   U48383 : BUF_X1 port map( A => n62060, Z => n68099);
   U48384 : BUF_X1 port map( A => n62058, Z => n68102);
   U48385 : BUF_X1 port map( A => n62056, Z => n68105);
   U48386 : BUF_X1 port map( A => n62054, Z => n68108);
   U48387 : BUF_X1 port map( A => n62052, Z => n68111);
   U48388 : BUF_X1 port map( A => n62050, Z => n68114);
   U48389 : BUF_X1 port map( A => n62048, Z => n68117);
   U48390 : BUF_X1 port map( A => n62046, Z => n68120);
   U48391 : BUF_X1 port map( A => n62044, Z => n68123);
   U48392 : BUF_X1 port map( A => n62042, Z => n68126);
   U48393 : BUF_X1 port map( A => n62040, Z => n68129);
   U48394 : BUF_X1 port map( A => n62038, Z => n68132);
   U48395 : BUF_X1 port map( A => n62036, Z => n68135);
   U48396 : BUF_X1 port map( A => n62034, Z => n68138);
   U48397 : BUF_X1 port map( A => n62032, Z => n68141);
   U48398 : BUF_X1 port map( A => n62030, Z => n68144);
   U48399 : BUF_X1 port map( A => n62028, Z => n68147);
   U48400 : BUF_X1 port map( A => n62026, Z => n68150);
   U48401 : BUF_X1 port map( A => n62024, Z => n68153);
   U48402 : BUF_X1 port map( A => n62022, Z => n68156);
   U48403 : BUF_X1 port map( A => n62020, Z => n68159);
   U48404 : BUF_X1 port map( A => n62018, Z => n68162);
   U48405 : BUF_X1 port map( A => n62016, Z => n68165);
   U48406 : BUF_X1 port map( A => n62014, Z => n68168);
   U48407 : BUF_X1 port map( A => n62012, Z => n68171);
   U48408 : BUF_X1 port map( A => n62010, Z => n68174);
   U48409 : BUF_X1 port map( A => n62008, Z => n68177);
   U48410 : BUF_X1 port map( A => n62006, Z => n68180);
   U48411 : BUF_X1 port map( A => n62004, Z => n68183);
   U48412 : BUF_X1 port map( A => n62002, Z => n68186);
   U48413 : BUF_X1 port map( A => n62000, Z => n68189);
   U48414 : BUF_X1 port map( A => n61998, Z => n68192);
   U48415 : BUF_X1 port map( A => n61996, Z => n68195);
   U48416 : BUF_X1 port map( A => n61994, Z => n68198);
   U48417 : BUF_X1 port map( A => n61992, Z => n68201);
   U48418 : BUF_X1 port map( A => n61990, Z => n68204);
   U48419 : BUF_X1 port map( A => n61988, Z => n68207);
   U48420 : BUF_X1 port map( A => n61986, Z => n68210);
   U48421 : BUF_X1 port map( A => n61984, Z => n68213);
   U48422 : BUF_X1 port map( A => n61982, Z => n68216);
   U48423 : BUF_X1 port map( A => n61980, Z => n68219);
   U48424 : BUF_X1 port map( A => n61978, Z => n68222);
   U48425 : BUF_X1 port map( A => n61976, Z => n68225);
   U48426 : BUF_X1 port map( A => n61974, Z => n68228);
   U48427 : BUF_X1 port map( A => n61972, Z => n68231);
   U48428 : BUF_X1 port map( A => n61970, Z => n68234);
   U48429 : BUF_X1 port map( A => n61968, Z => n68237);
   U48430 : BUF_X1 port map( A => n61966, Z => n68240);
   U48431 : BUF_X1 port map( A => n61964, Z => n68243);
   U48432 : BUF_X1 port map( A => n61962, Z => n68246);
   U48433 : BUF_X1 port map( A => n61960, Z => n68249);
   U48434 : OAI21_X1 port map( B1 => n62489, B2 => n62625, A => n68053, ZN => 
                           n62826);
   U48435 : OAI21_X1 port map( B1 => n62356, B2 => n63495, A => n68053, ZN => 
                           n63632);
   U48436 : OAI21_X1 port map( B1 => n62089, B2 => n62692, A => n68052, ZN => 
                           n62626);
   U48437 : OAI21_X1 port map( B1 => n62089, B2 => n62625, A => n68052, ZN => 
                           n62559);
   U48438 : OAI21_X1 port map( B1 => n62356, B2 => n63025, A => n68053, ZN => 
                           n63161);
   U48439 : OAI21_X1 port map( B1 => n62089, B2 => n63495, A => n68054, ZN => 
                           n63429);
   U48440 : OAI21_X1 port map( B1 => n62489, B2 => n63495, A => n68053, ZN => 
                           n63764);
   U48441 : OAI21_X1 port map( B1 => n62489, B2 => n63025, A => n68054, ZN => 
                           n63229);
   U48442 : OAI21_X1 port map( B1 => n62223, B2 => n63495, A => n68054, ZN => 
                           n63500);
   U48443 : OAI21_X1 port map( B1 => n62089, B2 => n63092, A => n68053, ZN => 
                           n63026);
   U48444 : OAI21_X1 port map( B1 => n62089, B2 => n63428, A => n68054, ZN => 
                           n63362);
   U48445 : OAI21_X1 port map( B1 => n62223, B2 => n63092, A => n68053, ZN => 
                           n63095);
   U48446 : OAI21_X1 port map( B1 => n62489, B2 => n63428, A => n68054, ZN => 
                           n63698);
   U48447 : OAI21_X1 port map( B1 => n62489, B2 => n63092, A => n68054, ZN => 
                           n63296);
   U48448 : OAI21_X1 port map( B1 => n62356, B2 => n63428, A => n68054, ZN => 
                           n63566);
   U48449 : OAI21_X1 port map( B1 => n62489, B2 => n62692, A => n68053, ZN => 
                           n62892);
   U48450 : OAI21_X1 port map( B1 => n62356, B2 => n62692, A => n68053, ZN => 
                           n62764);
   U48451 : OAI21_X1 port map( B1 => n62223, B2 => n62692, A => n68052, ZN => 
                           n62696);
   U48452 : OAI21_X1 port map( B1 => n62089, B2 => n62156, A => n68052, ZN => 
                           n62090);
   U48453 : NAND2_X1 port map( A1 => n65075, A2 => n65082, ZN => n63780);
   U48454 : NAND2_X1 port map( A1 => n65074, A2 => n65081, ZN => n63809);
   U48455 : NAND2_X1 port map( A1 => n65075, A2 => n65073, ZN => n63791);
   U48456 : AND2_X1 port map( A1 => n66281, A2 => n66279, ZN => n65117);
   U48457 : AND2_X1 port map( A1 => n66281, A2 => n66287, ZN => n65146);
   U48458 : AND2_X1 port map( A1 => n65085, A2 => n65078, ZN => n63794);
   U48459 : AND2_X1 port map( A1 => n65080, A2 => n65086, ZN => n63795);
   U48460 : AND2_X1 port map( A1 => n65073, A2 => n65086, ZN => n63788);
   U48461 : AND2_X1 port map( A1 => n65082, A2 => n65078, ZN => n63811);
   U48462 : AND2_X1 port map( A1 => n65087, A2 => n65078, ZN => n63815);
   U48463 : AND2_X1 port map( A1 => n65087, A2 => n65086, ZN => n63816);
   U48464 : AND2_X1 port map( A1 => n66286, A2 => n66278, ZN => n65121);
   U48465 : AND2_X1 port map( A1 => n66289, A2 => n66278, ZN => n65126);
   U48466 : AND2_X1 port map( A1 => n66285, A2 => n66278, ZN => n65142);
   U48467 : AND2_X1 port map( A1 => n66285, A2 => n66281, ZN => n65122);
   U48468 : AND2_X1 port map( A1 => n66289, A2 => n66281, ZN => n65127);
   U48469 : AND2_X1 port map( A1 => n66280, A2 => n66277, ZN => n65116);
   U48470 : AND2_X1 port map( A1 => n66285, A2 => n66277, ZN => n65141);
   U48471 : AND2_X1 port map( A1 => n66286, A2 => n66277, ZN => n65147);
   U48472 : AND2_X1 port map( A1 => n65077, A2 => n65074, ZN => n63810);
   U48473 : AND2_X1 port map( A1 => n65073, A2 => n65074, ZN => n63778);
   U48474 : AND2_X1 port map( A1 => n65080, A2 => n65074, ZN => n63783);
   U48475 : AND2_X1 port map( A1 => n65074, A2 => n65076, ZN => n63784);
   U48476 : NOR3_X1 port map( A1 => n66297, A2 => ADD_RD2(3), A3 => n66291, ZN 
                           => n66290);
   U48477 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n65094,
                           ZN => n65081);
   U48478 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n66292,
                           ZN => n66279);
   U48479 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n66287);
   U48480 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n65095,
                           ZN => n65076);
   U48481 : NOR3_X1 port map( A1 => n65095, A2 => ADD_RD1(0), A3 => n65093, ZN 
                           => n65077);
   U48482 : NOR3_X1 port map( A1 => n65094, A2 => ADD_RD1(3), A3 => n65095, ZN 
                           => n65082);
   U48483 : NOR3_X1 port map( A1 => n66291, A2 => ADD_RD2(0), A3 => n66292, ZN 
                           => n66280);
   U48484 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n65093,
                           ZN => n65073);
   U48485 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n65087);
   U48486 : NOR3_X1 port map( A1 => n66297, A2 => ADD_RD2(4), A3 => n66292, ZN 
                           => n66289);
   U48487 : NOR3_X1 port map( A1 => n65094, A2 => ADD_RD1(4), A3 => n65093, ZN 
                           => n65080);
   U48488 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n66297,
                           ZN => n66286);
   U48489 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n66291,
                           ZN => n66285);
   U48490 : NOR4_X1 port map( A1 => n66271, A2 => n66272, A3 => n66273, A4 => 
                           n66274, ZN => n66270);
   U48491 : OAI221_X1 port map( B1 => n63631, B2 => n67380, C1 => n7489, C2 => 
                           n67374, A => n66288, ZN => n66271);
   U48492 : OAI221_X1 port map( B1 => n62488, B2 => n67404, C1 => n63697, C2 =>
                           n67398, A => n66284, ZN => n66272);
   U48493 : OAI221_X1 port map( B1 => n54670, B2 => n67428, C1 => n63565, C2 =>
                           n67422, A => n66282, ZN => n66273);
   U48494 : NOR4_X1 port map( A1 => n66253, A2 => n66254, A3 => n66255, A4 => 
                           n66256, ZN => n66252);
   U48495 : OAI221_X1 port map( B1 => n63630, B2 => n67380, C1 => n7505, C2 => 
                           n67374, A => n66260, ZN => n66253);
   U48496 : OAI221_X1 port map( B1 => n62487, B2 => n67404, C1 => n63696, C2 =>
                           n67398, A => n66259, ZN => n66254);
   U48497 : OAI221_X1 port map( B1 => n54669, B2 => n67428, C1 => n63564, C2 =>
                           n67422, A => n66258, ZN => n66255);
   U48498 : NOR4_X1 port map( A1 => n66235, A2 => n66236, A3 => n66237, A4 => 
                           n66238, ZN => n66234);
   U48499 : OAI221_X1 port map( B1 => n63629, B2 => n67380, C1 => n7521, C2 => 
                           n67374, A => n66242, ZN => n66235);
   U48500 : OAI221_X1 port map( B1 => n62486, B2 => n67404, C1 => n63695, C2 =>
                           n67398, A => n66241, ZN => n66236);
   U48501 : OAI221_X1 port map( B1 => n54668, B2 => n67428, C1 => n63563, C2 =>
                           n67422, A => n66240, ZN => n66237);
   U48502 : NOR4_X1 port map( A1 => n66217, A2 => n66218, A3 => n66219, A4 => 
                           n66220, ZN => n66216);
   U48503 : OAI221_X1 port map( B1 => n63628, B2 => n67380, C1 => n7537, C2 => 
                           n67374, A => n66224, ZN => n66217);
   U48504 : OAI221_X1 port map( B1 => n62485, B2 => n67404, C1 => n63694, C2 =>
                           n67398, A => n66223, ZN => n66218);
   U48505 : OAI221_X1 port map( B1 => n54667, B2 => n67428, C1 => n63562, C2 =>
                           n67422, A => n66222, ZN => n66219);
   U48506 : NOR4_X1 port map( A1 => n66199, A2 => n66200, A3 => n66201, A4 => 
                           n66202, ZN => n66198);
   U48507 : OAI221_X1 port map( B1 => n63627, B2 => n67380, C1 => n7553, C2 => 
                           n67374, A => n66206, ZN => n66199);
   U48508 : OAI221_X1 port map( B1 => n62484, B2 => n67404, C1 => n63693, C2 =>
                           n67398, A => n66205, ZN => n66200);
   U48509 : OAI221_X1 port map( B1 => n54666, B2 => n67428, C1 => n63561, C2 =>
                           n67422, A => n66204, ZN => n66201);
   U48510 : NOR4_X1 port map( A1 => n66181, A2 => n66182, A3 => n66183, A4 => 
                           n66184, ZN => n66180);
   U48511 : OAI221_X1 port map( B1 => n63626, B2 => n67380, C1 => n7569, C2 => 
                           n67374, A => n66188, ZN => n66181);
   U48512 : OAI221_X1 port map( B1 => n62483, B2 => n67404, C1 => n63692, C2 =>
                           n67398, A => n66187, ZN => n66182);
   U48513 : OAI221_X1 port map( B1 => n54665, B2 => n67428, C1 => n63560, C2 =>
                           n67422, A => n66186, ZN => n66183);
   U48514 : NOR4_X1 port map( A1 => n66163, A2 => n66164, A3 => n66165, A4 => 
                           n66166, ZN => n66162);
   U48515 : OAI221_X1 port map( B1 => n63625, B2 => n67380, C1 => n7585, C2 => 
                           n67374, A => n66170, ZN => n66163);
   U48516 : OAI221_X1 port map( B1 => n62482, B2 => n67404, C1 => n63691, C2 =>
                           n67398, A => n66169, ZN => n66164);
   U48517 : OAI221_X1 port map( B1 => n54664, B2 => n67428, C1 => n63559, C2 =>
                           n67422, A => n66168, ZN => n66165);
   U48518 : NOR4_X1 port map( A1 => n66145, A2 => n66146, A3 => n66147, A4 => 
                           n66148, ZN => n66144);
   U48519 : OAI221_X1 port map( B1 => n63624, B2 => n67380, C1 => n7601, C2 => 
                           n67374, A => n66152, ZN => n66145);
   U48520 : OAI221_X1 port map( B1 => n62481, B2 => n67404, C1 => n63690, C2 =>
                           n67398, A => n66151, ZN => n66146);
   U48521 : OAI221_X1 port map( B1 => n54663, B2 => n67428, C1 => n63558, C2 =>
                           n67422, A => n66150, ZN => n66147);
   U48522 : NOR4_X1 port map( A1 => n66127, A2 => n66128, A3 => n66129, A4 => 
                           n66130, ZN => n66126);
   U48523 : OAI221_X1 port map( B1 => n63623, B2 => n67380, C1 => n7617, C2 => 
                           n67374, A => n66134, ZN => n66127);
   U48524 : OAI221_X1 port map( B1 => n62480, B2 => n67404, C1 => n63689, C2 =>
                           n67398, A => n66133, ZN => n66128);
   U48525 : OAI221_X1 port map( B1 => n54662, B2 => n67428, C1 => n63557, C2 =>
                           n67422, A => n66132, ZN => n66129);
   U48526 : NOR4_X1 port map( A1 => n66109, A2 => n66110, A3 => n66111, A4 => 
                           n66112, ZN => n66108);
   U48527 : OAI221_X1 port map( B1 => n63622, B2 => n67380, C1 => n7633, C2 => 
                           n67374, A => n66116, ZN => n66109);
   U48528 : OAI221_X1 port map( B1 => n62479, B2 => n67404, C1 => n63688, C2 =>
                           n67398, A => n66115, ZN => n66110);
   U48529 : OAI221_X1 port map( B1 => n54661, B2 => n67428, C1 => n63556, C2 =>
                           n67422, A => n66114, ZN => n66111);
   U48530 : NOR4_X1 port map( A1 => n66091, A2 => n66092, A3 => n66093, A4 => 
                           n66094, ZN => n66090);
   U48531 : OAI221_X1 port map( B1 => n63621, B2 => n67380, C1 => n7649, C2 => 
                           n67374, A => n66098, ZN => n66091);
   U48532 : OAI221_X1 port map( B1 => n62478, B2 => n67404, C1 => n63687, C2 =>
                           n67398, A => n66097, ZN => n66092);
   U48533 : OAI221_X1 port map( B1 => n54660, B2 => n67428, C1 => n63555, C2 =>
                           n67422, A => n66096, ZN => n66093);
   U48534 : NOR4_X1 port map( A1 => n66073, A2 => n66074, A3 => n66075, A4 => 
                           n66076, ZN => n66072);
   U48535 : OAI221_X1 port map( B1 => n63620, B2 => n67380, C1 => n7665, C2 => 
                           n67374, A => n66080, ZN => n66073);
   U48536 : OAI221_X1 port map( B1 => n62477, B2 => n67404, C1 => n63686, C2 =>
                           n67398, A => n66079, ZN => n66074);
   U48537 : OAI221_X1 port map( B1 => n54659, B2 => n67428, C1 => n63554, C2 =>
                           n67422, A => n66078, ZN => n66075);
   U48538 : NOR4_X1 port map( A1 => n66055, A2 => n66056, A3 => n66057, A4 => 
                           n66058, ZN => n66054);
   U48539 : OAI221_X1 port map( B1 => n63619, B2 => n67381, C1 => n7681, C2 => 
                           n67375, A => n66062, ZN => n66055);
   U48540 : OAI221_X1 port map( B1 => n62476, B2 => n67405, C1 => n63685, C2 =>
                           n67399, A => n66061, ZN => n66056);
   U48541 : OAI221_X1 port map( B1 => n63415, B2 => n67453, C1 => n49244, C2 =>
                           n67447, A => n66059, ZN => n66058);
   U48542 : NOR4_X1 port map( A1 => n66037, A2 => n66038, A3 => n66039, A4 => 
                           n66040, ZN => n66036);
   U48543 : OAI221_X1 port map( B1 => n63618, B2 => n67381, C1 => n7697, C2 => 
                           n67375, A => n66044, ZN => n66037);
   U48544 : OAI221_X1 port map( B1 => n62475, B2 => n67405, C1 => n63684, C2 =>
                           n67399, A => n66043, ZN => n66038);
   U48545 : OAI221_X1 port map( B1 => n63414, B2 => n67453, C1 => n49245, C2 =>
                           n67447, A => n66041, ZN => n66040);
   U48546 : NOR4_X1 port map( A1 => n66019, A2 => n66020, A3 => n66021, A4 => 
                           n66022, ZN => n66018);
   U48547 : OAI221_X1 port map( B1 => n63617, B2 => n67381, C1 => n7713, C2 => 
                           n67375, A => n66026, ZN => n66019);
   U48548 : OAI221_X1 port map( B1 => n62474, B2 => n67405, C1 => n63683, C2 =>
                           n67399, A => n66025, ZN => n66020);
   U48549 : OAI221_X1 port map( B1 => n63413, B2 => n67453, C1 => n49246, C2 =>
                           n67447, A => n66023, ZN => n66022);
   U48550 : NOR4_X1 port map( A1 => n66001, A2 => n66002, A3 => n66003, A4 => 
                           n66004, ZN => n66000);
   U48551 : OAI221_X1 port map( B1 => n63616, B2 => n67381, C1 => n7729, C2 => 
                           n67375, A => n66008, ZN => n66001);
   U48552 : OAI221_X1 port map( B1 => n62473, B2 => n67405, C1 => n63682, C2 =>
                           n67399, A => n66007, ZN => n66002);
   U48553 : OAI221_X1 port map( B1 => n63412, B2 => n67453, C1 => n49247, C2 =>
                           n67447, A => n66005, ZN => n66004);
   U48554 : NOR4_X1 port map( A1 => n65983, A2 => n65984, A3 => n65985, A4 => 
                           n65986, ZN => n65982);
   U48555 : OAI221_X1 port map( B1 => n63615, B2 => n67381, C1 => n7745, C2 => 
                           n67375, A => n65990, ZN => n65983);
   U48556 : OAI221_X1 port map( B1 => n62472, B2 => n67405, C1 => n63681, C2 =>
                           n67399, A => n65989, ZN => n65984);
   U48557 : OAI221_X1 port map( B1 => n63411, B2 => n67453, C1 => n49248, C2 =>
                           n67447, A => n65987, ZN => n65986);
   U48558 : NOR4_X1 port map( A1 => n65965, A2 => n65966, A3 => n65967, A4 => 
                           n65968, ZN => n65964);
   U48559 : OAI221_X1 port map( B1 => n63614, B2 => n67381, C1 => n7761, C2 => 
                           n67375, A => n65972, ZN => n65965);
   U48560 : OAI221_X1 port map( B1 => n62471, B2 => n67405, C1 => n63680, C2 =>
                           n67399, A => n65971, ZN => n65966);
   U48561 : OAI221_X1 port map( B1 => n63410, B2 => n67453, C1 => n49249, C2 =>
                           n67447, A => n65969, ZN => n65968);
   U48562 : NOR4_X1 port map( A1 => n65947, A2 => n65948, A3 => n65949, A4 => 
                           n65950, ZN => n65946);
   U48563 : OAI221_X1 port map( B1 => n63613, B2 => n67381, C1 => n7777, C2 => 
                           n67375, A => n65954, ZN => n65947);
   U48564 : OAI221_X1 port map( B1 => n62470, B2 => n67405, C1 => n63679, C2 =>
                           n67399, A => n65953, ZN => n65948);
   U48565 : OAI221_X1 port map( B1 => n63409, B2 => n67453, C1 => n49250, C2 =>
                           n67447, A => n65951, ZN => n65950);
   U48566 : NOR4_X1 port map( A1 => n65929, A2 => n65930, A3 => n65931, A4 => 
                           n65932, ZN => n65928);
   U48567 : OAI221_X1 port map( B1 => n63612, B2 => n67381, C1 => n7793, C2 => 
                           n67375, A => n65936, ZN => n65929);
   U48568 : OAI221_X1 port map( B1 => n62469, B2 => n67405, C1 => n63678, C2 =>
                           n67399, A => n65935, ZN => n65930);
   U48569 : OAI221_X1 port map( B1 => n63408, B2 => n67453, C1 => n49251, C2 =>
                           n67447, A => n65933, ZN => n65932);
   U48570 : NOR4_X1 port map( A1 => n65911, A2 => n65912, A3 => n65913, A4 => 
                           n65914, ZN => n65910);
   U48571 : OAI221_X1 port map( B1 => n63611, B2 => n67381, C1 => n7809, C2 => 
                           n67375, A => n65918, ZN => n65911);
   U48572 : OAI221_X1 port map( B1 => n62468, B2 => n67405, C1 => n63677, C2 =>
                           n67399, A => n65917, ZN => n65912);
   U48573 : OAI221_X1 port map( B1 => n63407, B2 => n67453, C1 => n49252, C2 =>
                           n67447, A => n65915, ZN => n65914);
   U48574 : NOR4_X1 port map( A1 => n65893, A2 => n65894, A3 => n65895, A4 => 
                           n65896, ZN => n65892);
   U48575 : OAI221_X1 port map( B1 => n63610, B2 => n67381, C1 => n7825, C2 => 
                           n67375, A => n65900, ZN => n65893);
   U48576 : OAI221_X1 port map( B1 => n62467, B2 => n67405, C1 => n63676, C2 =>
                           n67399, A => n65899, ZN => n65894);
   U48577 : OAI221_X1 port map( B1 => n63406, B2 => n67453, C1 => n49253, C2 =>
                           n67447, A => n65897, ZN => n65896);
   U48578 : NOR4_X1 port map( A1 => n65875, A2 => n65876, A3 => n65877, A4 => 
                           n65878, ZN => n65874);
   U48579 : OAI221_X1 port map( B1 => n63609, B2 => n67381, C1 => n7841, C2 => 
                           n67375, A => n65882, ZN => n65875);
   U48580 : OAI221_X1 port map( B1 => n62466, B2 => n67405, C1 => n63675, C2 =>
                           n67399, A => n65881, ZN => n65876);
   U48581 : OAI221_X1 port map( B1 => n63405, B2 => n67453, C1 => n49254, C2 =>
                           n67447, A => n65879, ZN => n65878);
   U48582 : NOR4_X1 port map( A1 => n65857, A2 => n65858, A3 => n65859, A4 => 
                           n65860, ZN => n65856);
   U48583 : OAI221_X1 port map( B1 => n63608, B2 => n67381, C1 => n7857, C2 => 
                           n67375, A => n65864, ZN => n65857);
   U48584 : OAI221_X1 port map( B1 => n62465, B2 => n67405, C1 => n63674, C2 =>
                           n67399, A => n65863, ZN => n65858);
   U48585 : OAI221_X1 port map( B1 => n63404, B2 => n67453, C1 => n49255, C2 =>
                           n67447, A => n65861, ZN => n65860);
   U48586 : NOR4_X1 port map( A1 => n65839, A2 => n65840, A3 => n65841, A4 => 
                           n65842, ZN => n65838);
   U48587 : OAI221_X1 port map( B1 => n63607, B2 => n67382, C1 => n7873, C2 => 
                           n67376, A => n65846, ZN => n65839);
   U48588 : OAI221_X1 port map( B1 => n62464, B2 => n67406, C1 => n63673, C2 =>
                           n67400, A => n65845, ZN => n65840);
   U48589 : OAI221_X1 port map( B1 => n63403, B2 => n67454, C1 => n49256, C2 =>
                           n67448, A => n65843, ZN => n65842);
   U48590 : NOR4_X1 port map( A1 => n65821, A2 => n65822, A3 => n65823, A4 => 
                           n65824, ZN => n65820);
   U48591 : OAI221_X1 port map( B1 => n63606, B2 => n67382, C1 => n7889, C2 => 
                           n67376, A => n65828, ZN => n65821);
   U48592 : OAI221_X1 port map( B1 => n62463, B2 => n67406, C1 => n63672, C2 =>
                           n67400, A => n65827, ZN => n65822);
   U48593 : OAI221_X1 port map( B1 => n63402, B2 => n67454, C1 => n49257, C2 =>
                           n67448, A => n65825, ZN => n65824);
   U48594 : NOR4_X1 port map( A1 => n65803, A2 => n65804, A3 => n65805, A4 => 
                           n65806, ZN => n65802);
   U48595 : OAI221_X1 port map( B1 => n63605, B2 => n67382, C1 => n7905, C2 => 
                           n67376, A => n65810, ZN => n65803);
   U48596 : OAI221_X1 port map( B1 => n62462, B2 => n67406, C1 => n63671, C2 =>
                           n67400, A => n65809, ZN => n65804);
   U48597 : OAI221_X1 port map( B1 => n63401, B2 => n67454, C1 => n49258, C2 =>
                           n67448, A => n65807, ZN => n65806);
   U48598 : NOR4_X1 port map( A1 => n65785, A2 => n65786, A3 => n65787, A4 => 
                           n65788, ZN => n65784);
   U48599 : OAI221_X1 port map( B1 => n63604, B2 => n67382, C1 => n7921, C2 => 
                           n67376, A => n65792, ZN => n65785);
   U48600 : OAI221_X1 port map( B1 => n62461, B2 => n67406, C1 => n63670, C2 =>
                           n67400, A => n65791, ZN => n65786);
   U48601 : OAI221_X1 port map( B1 => n63400, B2 => n67454, C1 => n49259, C2 =>
                           n67448, A => n65789, ZN => n65788);
   U48602 : NOR4_X1 port map( A1 => n65767, A2 => n65768, A3 => n65769, A4 => 
                           n65770, ZN => n65766);
   U48603 : OAI221_X1 port map( B1 => n63603, B2 => n67382, C1 => n7937, C2 => 
                           n67376, A => n65774, ZN => n65767);
   U48604 : OAI221_X1 port map( B1 => n62460, B2 => n67406, C1 => n63669, C2 =>
                           n67400, A => n65773, ZN => n65768);
   U48605 : OAI221_X1 port map( B1 => n63399, B2 => n67454, C1 => n49260, C2 =>
                           n67448, A => n65771, ZN => n65770);
   U48606 : NOR4_X1 port map( A1 => n65749, A2 => n65750, A3 => n65751, A4 => 
                           n65752, ZN => n65748);
   U48607 : OAI221_X1 port map( B1 => n63602, B2 => n67382, C1 => n7953, C2 => 
                           n67376, A => n65756, ZN => n65749);
   U48608 : OAI221_X1 port map( B1 => n62459, B2 => n67406, C1 => n63668, C2 =>
                           n67400, A => n65755, ZN => n65750);
   U48609 : OAI221_X1 port map( B1 => n63398, B2 => n67454, C1 => n49261, C2 =>
                           n67448, A => n65753, ZN => n65752);
   U48610 : NOR4_X1 port map( A1 => n65731, A2 => n65732, A3 => n65733, A4 => 
                           n65734, ZN => n65730);
   U48611 : OAI221_X1 port map( B1 => n63601, B2 => n67382, C1 => n7969, C2 => 
                           n67376, A => n65738, ZN => n65731);
   U48612 : OAI221_X1 port map( B1 => n62458, B2 => n67406, C1 => n63667, C2 =>
                           n67400, A => n65737, ZN => n65732);
   U48613 : OAI221_X1 port map( B1 => n63397, B2 => n67454, C1 => n49262, C2 =>
                           n67448, A => n65735, ZN => n65734);
   U48614 : NOR4_X1 port map( A1 => n65713, A2 => n65714, A3 => n65715, A4 => 
                           n65716, ZN => n65712);
   U48615 : OAI221_X1 port map( B1 => n63600, B2 => n67382, C1 => n7985, C2 => 
                           n67376, A => n65720, ZN => n65713);
   U48616 : OAI221_X1 port map( B1 => n62457, B2 => n67406, C1 => n63666, C2 =>
                           n67400, A => n65719, ZN => n65714);
   U48617 : OAI221_X1 port map( B1 => n63396, B2 => n67454, C1 => n49263, C2 =>
                           n67448, A => n65717, ZN => n65716);
   U48618 : NOR4_X1 port map( A1 => n65695, A2 => n65696, A3 => n65697, A4 => 
                           n65698, ZN => n65694);
   U48619 : OAI221_X1 port map( B1 => n63599, B2 => n67382, C1 => n8001, C2 => 
                           n67376, A => n65702, ZN => n65695);
   U48620 : OAI221_X1 port map( B1 => n62456, B2 => n67406, C1 => n63665, C2 =>
                           n67400, A => n65701, ZN => n65696);
   U48621 : OAI221_X1 port map( B1 => n63395, B2 => n67454, C1 => n49264, C2 =>
                           n67448, A => n65699, ZN => n65698);
   U48622 : NOR4_X1 port map( A1 => n65677, A2 => n65678, A3 => n65679, A4 => 
                           n65680, ZN => n65676);
   U48623 : OAI221_X1 port map( B1 => n63598, B2 => n67382, C1 => n8017, C2 => 
                           n67376, A => n65684, ZN => n65677);
   U48624 : OAI221_X1 port map( B1 => n62455, B2 => n67406, C1 => n63664, C2 =>
                           n67400, A => n65683, ZN => n65678);
   U48625 : OAI221_X1 port map( B1 => n63394, B2 => n67454, C1 => n49265, C2 =>
                           n67448, A => n65681, ZN => n65680);
   U48626 : NOR4_X1 port map( A1 => n65659, A2 => n65660, A3 => n65661, A4 => 
                           n65662, ZN => n65658);
   U48627 : OAI221_X1 port map( B1 => n63597, B2 => n67382, C1 => n8033, C2 => 
                           n67376, A => n65666, ZN => n65659);
   U48628 : OAI221_X1 port map( B1 => n62454, B2 => n67406, C1 => n63663, C2 =>
                           n67400, A => n65665, ZN => n65660);
   U48629 : OAI221_X1 port map( B1 => n63393, B2 => n67454, C1 => n49266, C2 =>
                           n67448, A => n65663, ZN => n65662);
   U48630 : NOR4_X1 port map( A1 => n65641, A2 => n65642, A3 => n65643, A4 => 
                           n65644, ZN => n65640);
   U48631 : OAI221_X1 port map( B1 => n63596, B2 => n67382, C1 => n8049, C2 => 
                           n67376, A => n65648, ZN => n65641);
   U48632 : OAI221_X1 port map( B1 => n62453, B2 => n67406, C1 => n63662, C2 =>
                           n67400, A => n65647, ZN => n65642);
   U48633 : OAI221_X1 port map( B1 => n63392, B2 => n67454, C1 => n49267, C2 =>
                           n67448, A => n65645, ZN => n65644);
   U48634 : NOR4_X1 port map( A1 => n65623, A2 => n65624, A3 => n65625, A4 => 
                           n65626, ZN => n65622);
   U48635 : OAI221_X1 port map( B1 => n63595, B2 => n67383, C1 => n8065, C2 => 
                           n67377, A => n65630, ZN => n65623);
   U48636 : OAI221_X1 port map( B1 => n62452, B2 => n67407, C1 => n63661, C2 =>
                           n67401, A => n65629, ZN => n65624);
   U48637 : OAI221_X1 port map( B1 => n63391, B2 => n67455, C1 => n49268, C2 =>
                           n67449, A => n65627, ZN => n65626);
   U48638 : NOR4_X1 port map( A1 => n65605, A2 => n65606, A3 => n65607, A4 => 
                           n65608, ZN => n65604);
   U48639 : OAI221_X1 port map( B1 => n63594, B2 => n67383, C1 => n8081, C2 => 
                           n67377, A => n65612, ZN => n65605);
   U48640 : OAI221_X1 port map( B1 => n62451, B2 => n67407, C1 => n63660, C2 =>
                           n67401, A => n65611, ZN => n65606);
   U48641 : OAI221_X1 port map( B1 => n63390, B2 => n67455, C1 => n49269, C2 =>
                           n67449, A => n65609, ZN => n65608);
   U48642 : NOR4_X1 port map( A1 => n65587, A2 => n65588, A3 => n65589, A4 => 
                           n65590, ZN => n65586);
   U48643 : OAI221_X1 port map( B1 => n63593, B2 => n67383, C1 => n8097, C2 => 
                           n67377, A => n65594, ZN => n65587);
   U48644 : OAI221_X1 port map( B1 => n62450, B2 => n67407, C1 => n63659, C2 =>
                           n67401, A => n65593, ZN => n65588);
   U48645 : OAI221_X1 port map( B1 => n63389, B2 => n67455, C1 => n49270, C2 =>
                           n67449, A => n65591, ZN => n65590);
   U48646 : NOR4_X1 port map( A1 => n65569, A2 => n65570, A3 => n65571, A4 => 
                           n65572, ZN => n65568);
   U48647 : OAI221_X1 port map( B1 => n63592, B2 => n67383, C1 => n8113, C2 => 
                           n67377, A => n65576, ZN => n65569);
   U48648 : OAI221_X1 port map( B1 => n62449, B2 => n67407, C1 => n63658, C2 =>
                           n67401, A => n65575, ZN => n65570);
   U48649 : OAI221_X1 port map( B1 => n63388, B2 => n67455, C1 => n49271, C2 =>
                           n67449, A => n65573, ZN => n65572);
   U48650 : NOR4_X1 port map( A1 => n65551, A2 => n65552, A3 => n65553, A4 => 
                           n65554, ZN => n65550);
   U48651 : OAI221_X1 port map( B1 => n63591, B2 => n67383, C1 => n8129, C2 => 
                           n67377, A => n65558, ZN => n65551);
   U48652 : OAI221_X1 port map( B1 => n62448, B2 => n67407, C1 => n63657, C2 =>
                           n67401, A => n65557, ZN => n65552);
   U48653 : OAI221_X1 port map( B1 => n63387, B2 => n67455, C1 => n49272, C2 =>
                           n67449, A => n65555, ZN => n65554);
   U48654 : NOR4_X1 port map( A1 => n65533, A2 => n65534, A3 => n65535, A4 => 
                           n65536, ZN => n65532);
   U48655 : OAI221_X1 port map( B1 => n63590, B2 => n67383, C1 => n8145, C2 => 
                           n67377, A => n65540, ZN => n65533);
   U48656 : OAI221_X1 port map( B1 => n62447, B2 => n67407, C1 => n63656, C2 =>
                           n67401, A => n65539, ZN => n65534);
   U48657 : OAI221_X1 port map( B1 => n63386, B2 => n67455, C1 => n49273, C2 =>
                           n67449, A => n65537, ZN => n65536);
   U48658 : NOR4_X1 port map( A1 => n65515, A2 => n65516, A3 => n65517, A4 => 
                           n65518, ZN => n65514);
   U48659 : OAI221_X1 port map( B1 => n63589, B2 => n67383, C1 => n8161, C2 => 
                           n67377, A => n65522, ZN => n65515);
   U48660 : OAI221_X1 port map( B1 => n62446, B2 => n67407, C1 => n63655, C2 =>
                           n67401, A => n65521, ZN => n65516);
   U48661 : OAI221_X1 port map( B1 => n63385, B2 => n67455, C1 => n49274, C2 =>
                           n67449, A => n65519, ZN => n65518);
   U48662 : NOR4_X1 port map( A1 => n65497, A2 => n65498, A3 => n65499, A4 => 
                           n65500, ZN => n65496);
   U48663 : OAI221_X1 port map( B1 => n63588, B2 => n67383, C1 => n8177, C2 => 
                           n67377, A => n65504, ZN => n65497);
   U48664 : OAI221_X1 port map( B1 => n62445, B2 => n67407, C1 => n63654, C2 =>
                           n67401, A => n65503, ZN => n65498);
   U48665 : OAI221_X1 port map( B1 => n63384, B2 => n67455, C1 => n49275, C2 =>
                           n67449, A => n65501, ZN => n65500);
   U48666 : NOR4_X1 port map( A1 => n65479, A2 => n65480, A3 => n65481, A4 => 
                           n65482, ZN => n65478);
   U48667 : OAI221_X1 port map( B1 => n63587, B2 => n67383, C1 => n8193, C2 => 
                           n67377, A => n65486, ZN => n65479);
   U48668 : OAI221_X1 port map( B1 => n62444, B2 => n67407, C1 => n63653, C2 =>
                           n67401, A => n65485, ZN => n65480);
   U48669 : OAI221_X1 port map( B1 => n63383, B2 => n67455, C1 => n49276, C2 =>
                           n67449, A => n65483, ZN => n65482);
   U48670 : NOR4_X1 port map( A1 => n65461, A2 => n65462, A3 => n65463, A4 => 
                           n65464, ZN => n65460);
   U48671 : OAI221_X1 port map( B1 => n63586, B2 => n67383, C1 => n8209, C2 => 
                           n67377, A => n65468, ZN => n65461);
   U48672 : OAI221_X1 port map( B1 => n62443, B2 => n67407, C1 => n63652, C2 =>
                           n67401, A => n65467, ZN => n65462);
   U48673 : OAI221_X1 port map( B1 => n63382, B2 => n67455, C1 => n49277, C2 =>
                           n67449, A => n65465, ZN => n65464);
   U48674 : NOR4_X1 port map( A1 => n65443, A2 => n65444, A3 => n65445, A4 => 
                           n65446, ZN => n65442);
   U48675 : OAI221_X1 port map( B1 => n63585, B2 => n67383, C1 => n8225, C2 => 
                           n67377, A => n65450, ZN => n65443);
   U48676 : OAI221_X1 port map( B1 => n62442, B2 => n67407, C1 => n63651, C2 =>
                           n67401, A => n65449, ZN => n65444);
   U48677 : OAI221_X1 port map( B1 => n63381, B2 => n67455, C1 => n49278, C2 =>
                           n67449, A => n65447, ZN => n65446);
   U48678 : NOR4_X1 port map( A1 => n65425, A2 => n65426, A3 => n65427, A4 => 
                           n65428, ZN => n65424);
   U48679 : OAI221_X1 port map( B1 => n63584, B2 => n67383, C1 => n8241, C2 => 
                           n67377, A => n65432, ZN => n65425);
   U48680 : OAI221_X1 port map( B1 => n62441, B2 => n67407, C1 => n63650, C2 =>
                           n67401, A => n65431, ZN => n65426);
   U48681 : OAI221_X1 port map( B1 => n63380, B2 => n67455, C1 => n49279, C2 =>
                           n67449, A => n65429, ZN => n65428);
   U48682 : NOR4_X1 port map( A1 => n65407, A2 => n65408, A3 => n65409, A4 => 
                           n65410, ZN => n65406);
   U48683 : OAI221_X1 port map( B1 => n63583, B2 => n67384, C1 => n8257, C2 => 
                           n67378, A => n65414, ZN => n65407);
   U48684 : OAI221_X1 port map( B1 => n62440, B2 => n67408, C1 => n63649, C2 =>
                           n67402, A => n65413, ZN => n65408);
   U48685 : OAI221_X1 port map( B1 => n63379, B2 => n67456, C1 => n49280, C2 =>
                           n67450, A => n65411, ZN => n65410);
   U48686 : NOR4_X1 port map( A1 => n65389, A2 => n65390, A3 => n65391, A4 => 
                           n65392, ZN => n65388);
   U48687 : OAI221_X1 port map( B1 => n63582, B2 => n67384, C1 => n8273, C2 => 
                           n67378, A => n65396, ZN => n65389);
   U48688 : OAI221_X1 port map( B1 => n62439, B2 => n67408, C1 => n63648, C2 =>
                           n67402, A => n65395, ZN => n65390);
   U48689 : OAI221_X1 port map( B1 => n63378, B2 => n67456, C1 => n49281, C2 =>
                           n67450, A => n65393, ZN => n65392);
   U48690 : NOR4_X1 port map( A1 => n65371, A2 => n65372, A3 => n65373, A4 => 
                           n65374, ZN => n65370);
   U48691 : OAI221_X1 port map( B1 => n63581, B2 => n67384, C1 => n8289, C2 => 
                           n67378, A => n65378, ZN => n65371);
   U48692 : OAI221_X1 port map( B1 => n62438, B2 => n67408, C1 => n63647, C2 =>
                           n67402, A => n65377, ZN => n65372);
   U48693 : OAI221_X1 port map( B1 => n63377, B2 => n67456, C1 => n49282, C2 =>
                           n67450, A => n65375, ZN => n65374);
   U48694 : NOR4_X1 port map( A1 => n65353, A2 => n65354, A3 => n65355, A4 => 
                           n65356, ZN => n65352);
   U48695 : OAI221_X1 port map( B1 => n63580, B2 => n67384, C1 => n8305, C2 => 
                           n67378, A => n65360, ZN => n65353);
   U48696 : OAI221_X1 port map( B1 => n62437, B2 => n67408, C1 => n63646, C2 =>
                           n67402, A => n65359, ZN => n65354);
   U48697 : OAI221_X1 port map( B1 => n63376, B2 => n67456, C1 => n49283, C2 =>
                           n67450, A => n65357, ZN => n65356);
   U48698 : NOR4_X1 port map( A1 => n65335, A2 => n65336, A3 => n65337, A4 => 
                           n65338, ZN => n65334);
   U48699 : OAI221_X1 port map( B1 => n63579, B2 => n67384, C1 => n8321, C2 => 
                           n67378, A => n65342, ZN => n65335);
   U48700 : OAI221_X1 port map( B1 => n62436, B2 => n67408, C1 => n63645, C2 =>
                           n67402, A => n65341, ZN => n65336);
   U48701 : OAI221_X1 port map( B1 => n63375, B2 => n67456, C1 => n49284, C2 =>
                           n67450, A => n65339, ZN => n65338);
   U48702 : NOR4_X1 port map( A1 => n65317, A2 => n65318, A3 => n65319, A4 => 
                           n65320, ZN => n65316);
   U48703 : OAI221_X1 port map( B1 => n63578, B2 => n67384, C1 => n8337, C2 => 
                           n67378, A => n65324, ZN => n65317);
   U48704 : OAI221_X1 port map( B1 => n62435, B2 => n67408, C1 => n63644, C2 =>
                           n67402, A => n65323, ZN => n65318);
   U48705 : OAI221_X1 port map( B1 => n63374, B2 => n67456, C1 => n49285, C2 =>
                           n67450, A => n65321, ZN => n65320);
   U48706 : NOR4_X1 port map( A1 => n65299, A2 => n65300, A3 => n65301, A4 => 
                           n65302, ZN => n65298);
   U48707 : OAI221_X1 port map( B1 => n63577, B2 => n67384, C1 => n8353, C2 => 
                           n67378, A => n65306, ZN => n65299);
   U48708 : OAI221_X1 port map( B1 => n62434, B2 => n67408, C1 => n63643, C2 =>
                           n67402, A => n65305, ZN => n65300);
   U48709 : OAI221_X1 port map( B1 => n63373, B2 => n67456, C1 => n49286, C2 =>
                           n67450, A => n65303, ZN => n65302);
   U48710 : NOR4_X1 port map( A1 => n65281, A2 => n65282, A3 => n65283, A4 => 
                           n65284, ZN => n65280);
   U48711 : OAI221_X1 port map( B1 => n63576, B2 => n67384, C1 => n8369, C2 => 
                           n67378, A => n65288, ZN => n65281);
   U48712 : OAI221_X1 port map( B1 => n62433, B2 => n67408, C1 => n63642, C2 =>
                           n67402, A => n65287, ZN => n65282);
   U48713 : OAI221_X1 port map( B1 => n63372, B2 => n67456, C1 => n49287, C2 =>
                           n67450, A => n65285, ZN => n65284);
   U48714 : NOR4_X1 port map( A1 => n65263, A2 => n65264, A3 => n65265, A4 => 
                           n65266, ZN => n65262);
   U48715 : OAI221_X1 port map( B1 => n63575, B2 => n67384, C1 => n8385, C2 => 
                           n67378, A => n65270, ZN => n65263);
   U48716 : OAI221_X1 port map( B1 => n62432, B2 => n67408, C1 => n63641, C2 =>
                           n67402, A => n65269, ZN => n65264);
   U48717 : OAI221_X1 port map( B1 => n63371, B2 => n67456, C1 => n49288, C2 =>
                           n67450, A => n65267, ZN => n65266);
   U48718 : NOR4_X1 port map( A1 => n65245, A2 => n65246, A3 => n65247, A4 => 
                           n65248, ZN => n65244);
   U48719 : OAI221_X1 port map( B1 => n63574, B2 => n67384, C1 => n8401, C2 => 
                           n67378, A => n65252, ZN => n65245);
   U48720 : OAI221_X1 port map( B1 => n62431, B2 => n67408, C1 => n63640, C2 =>
                           n67402, A => n65251, ZN => n65246);
   U48721 : OAI221_X1 port map( B1 => n63370, B2 => n67456, C1 => n49289, C2 =>
                           n67450, A => n65249, ZN => n65248);
   U48722 : NOR4_X1 port map( A1 => n65227, A2 => n65228, A3 => n65229, A4 => 
                           n65230, ZN => n65226);
   U48723 : OAI221_X1 port map( B1 => n63573, B2 => n67384, C1 => n8417, C2 => 
                           n67378, A => n65234, ZN => n65227);
   U48724 : OAI221_X1 port map( B1 => n62430, B2 => n67408, C1 => n63639, C2 =>
                           n67402, A => n65233, ZN => n65228);
   U48725 : OAI221_X1 port map( B1 => n63369, B2 => n67456, C1 => n49290, C2 =>
                           n67450, A => n65231, ZN => n65230);
   U48726 : NOR4_X1 port map( A1 => n65209, A2 => n65210, A3 => n65211, A4 => 
                           n65212, ZN => n65208);
   U48727 : OAI221_X1 port map( B1 => n63572, B2 => n67384, C1 => n8433, C2 => 
                           n67378, A => n65216, ZN => n65209);
   U48728 : OAI221_X1 port map( B1 => n62429, B2 => n67408, C1 => n63638, C2 =>
                           n67402, A => n65215, ZN => n65210);
   U48729 : OAI221_X1 port map( B1 => n63368, B2 => n67456, C1 => n49291, C2 =>
                           n67450, A => n65213, ZN => n65212);
   U48730 : NOR4_X1 port map( A1 => n65068, A2 => n65069, A3 => n65070, A4 => 
                           n65071, ZN => n65067);
   U48731 : OAI221_X1 port map( B1 => n63160, B2 => n67626, C1 => n62289, C2 =>
                           n67620, A => n65079, ZN => n65070);
   U48732 : OAI221_X1 port map( B1 => n63427, B2 => n67648, C1 => n49420, C2 =>
                           n67642, A => n65072, ZN => n65071);
   U48733 : OAI221_X1 port map( B1 => n62488, B2 => n67602, C1 => n63565, C2 =>
                           n67596, A => n65083, ZN => n65069);
   U48734 : NOR4_X1 port map( A1 => n65048, A2 => n65049, A3 => n65050, A4 => 
                           n65051, ZN => n65047);
   U48735 : OAI221_X1 port map( B1 => n63159, B2 => n67626, C1 => n62288, C2 =>
                           n67620, A => n65053, ZN => n65050);
   U48736 : OAI221_X1 port map( B1 => n63426, B2 => n67648, C1 => n49421, C2 =>
                           n67642, A => n65052, ZN => n65051);
   U48737 : OAI221_X1 port map( B1 => n62487, B2 => n67602, C1 => n63564, C2 =>
                           n67596, A => n65054, ZN => n65049);
   U48738 : NOR4_X1 port map( A1 => n65028, A2 => n65029, A3 => n65030, A4 => 
                           n65031, ZN => n65027);
   U48739 : OAI221_X1 port map( B1 => n63158, B2 => n67626, C1 => n62287, C2 =>
                           n67620, A => n65033, ZN => n65030);
   U48740 : OAI221_X1 port map( B1 => n63425, B2 => n67648, C1 => n49422, C2 =>
                           n67642, A => n65032, ZN => n65031);
   U48741 : OAI221_X1 port map( B1 => n62486, B2 => n67602, C1 => n63563, C2 =>
                           n67596, A => n65034, ZN => n65029);
   U48742 : NOR4_X1 port map( A1 => n65008, A2 => n65009, A3 => n65010, A4 => 
                           n65011, ZN => n65007);
   U48743 : OAI221_X1 port map( B1 => n63157, B2 => n67626, C1 => n62286, C2 =>
                           n67620, A => n65013, ZN => n65010);
   U48744 : OAI221_X1 port map( B1 => n63424, B2 => n67648, C1 => n49423, C2 =>
                           n67642, A => n65012, ZN => n65011);
   U48745 : OAI221_X1 port map( B1 => n62485, B2 => n67602, C1 => n63562, C2 =>
                           n67596, A => n65014, ZN => n65009);
   U48746 : NOR4_X1 port map( A1 => n64988, A2 => n64989, A3 => n64990, A4 => 
                           n64991, ZN => n64987);
   U48747 : OAI221_X1 port map( B1 => n63156, B2 => n67626, C1 => n62285, C2 =>
                           n67620, A => n64993, ZN => n64990);
   U48748 : OAI221_X1 port map( B1 => n63423, B2 => n67648, C1 => n49424, C2 =>
                           n67642, A => n64992, ZN => n64991);
   U48749 : OAI221_X1 port map( B1 => n62484, B2 => n67602, C1 => n63561, C2 =>
                           n67596, A => n64994, ZN => n64989);
   U48750 : NOR4_X1 port map( A1 => n64968, A2 => n64969, A3 => n64970, A4 => 
                           n64971, ZN => n64967);
   U48751 : OAI221_X1 port map( B1 => n63155, B2 => n67626, C1 => n62284, C2 =>
                           n67620, A => n64973, ZN => n64970);
   U48752 : OAI221_X1 port map( B1 => n63422, B2 => n67648, C1 => n49425, C2 =>
                           n67642, A => n64972, ZN => n64971);
   U48753 : OAI221_X1 port map( B1 => n62483, B2 => n67602, C1 => n63560, C2 =>
                           n67596, A => n64974, ZN => n64969);
   U48754 : NOR4_X1 port map( A1 => n64948, A2 => n64949, A3 => n64950, A4 => 
                           n64951, ZN => n64947);
   U48755 : OAI221_X1 port map( B1 => n63154, B2 => n67626, C1 => n62283, C2 =>
                           n67620, A => n64953, ZN => n64950);
   U48756 : OAI221_X1 port map( B1 => n63421, B2 => n67648, C1 => n49426, C2 =>
                           n67642, A => n64952, ZN => n64951);
   U48757 : OAI221_X1 port map( B1 => n62482, B2 => n67602, C1 => n63559, C2 =>
                           n67596, A => n64954, ZN => n64949);
   U48758 : NOR4_X1 port map( A1 => n64928, A2 => n64929, A3 => n64930, A4 => 
                           n64931, ZN => n64927);
   U48759 : OAI221_X1 port map( B1 => n63153, B2 => n67626, C1 => n62282, C2 =>
                           n67620, A => n64933, ZN => n64930);
   U48760 : OAI221_X1 port map( B1 => n63420, B2 => n67648, C1 => n49427, C2 =>
                           n67642, A => n64932, ZN => n64931);
   U48761 : OAI221_X1 port map( B1 => n62481, B2 => n67602, C1 => n63558, C2 =>
                           n67596, A => n64934, ZN => n64929);
   U48762 : NOR4_X1 port map( A1 => n64908, A2 => n64909, A3 => n64910, A4 => 
                           n64911, ZN => n64907);
   U48763 : OAI221_X1 port map( B1 => n63152, B2 => n67626, C1 => n62281, C2 =>
                           n67620, A => n64913, ZN => n64910);
   U48764 : OAI221_X1 port map( B1 => n63419, B2 => n67648, C1 => n49428, C2 =>
                           n67642, A => n64912, ZN => n64911);
   U48765 : OAI221_X1 port map( B1 => n62480, B2 => n67602, C1 => n63557, C2 =>
                           n67596, A => n64914, ZN => n64909);
   U48766 : NOR4_X1 port map( A1 => n64888, A2 => n64889, A3 => n64890, A4 => 
                           n64891, ZN => n64887);
   U48767 : OAI221_X1 port map( B1 => n63151, B2 => n67626, C1 => n62280, C2 =>
                           n67620, A => n64893, ZN => n64890);
   U48768 : OAI221_X1 port map( B1 => n63418, B2 => n67648, C1 => n49429, C2 =>
                           n67642, A => n64892, ZN => n64891);
   U48769 : OAI221_X1 port map( B1 => n62479, B2 => n67602, C1 => n63556, C2 =>
                           n67596, A => n64894, ZN => n64889);
   U48770 : NOR4_X1 port map( A1 => n64868, A2 => n64869, A3 => n64870, A4 => 
                           n64871, ZN => n64867);
   U48771 : OAI221_X1 port map( B1 => n63150, B2 => n67626, C1 => n62279, C2 =>
                           n67620, A => n64873, ZN => n64870);
   U48772 : OAI221_X1 port map( B1 => n63417, B2 => n67648, C1 => n49430, C2 =>
                           n67642, A => n64872, ZN => n64871);
   U48773 : OAI221_X1 port map( B1 => n62478, B2 => n67602, C1 => n63555, C2 =>
                           n67596, A => n64874, ZN => n64869);
   U48774 : NOR4_X1 port map( A1 => n64848, A2 => n64849, A3 => n64850, A4 => 
                           n64851, ZN => n64847);
   U48775 : OAI221_X1 port map( B1 => n63149, B2 => n67626, C1 => n62278, C2 =>
                           n67620, A => n64853, ZN => n64850);
   U48776 : OAI221_X1 port map( B1 => n63416, B2 => n67648, C1 => n49431, C2 =>
                           n67642, A => n64852, ZN => n64851);
   U48777 : OAI221_X1 port map( B1 => n62477, B2 => n67602, C1 => n63554, C2 =>
                           n67596, A => n64854, ZN => n64849);
   U48778 : NOR4_X1 port map( A1 => n64828, A2 => n64829, A3 => n64830, A4 => 
                           n64831, ZN => n64827);
   U48779 : OAI221_X1 port map( B1 => n63148, B2 => n67627, C1 => n62277, C2 =>
                           n67621, A => n64833, ZN => n64830);
   U48780 : OAI221_X1 port map( B1 => n62476, B2 => n67603, C1 => n63553, C2 =>
                           n67597, A => n64834, ZN => n64829);
   U48781 : OAI221_X1 port map( B1 => n54234, B2 => n67579, C1 => n63619, C2 =>
                           n67573, A => n64836, ZN => n64828);
   U48782 : NOR4_X1 port map( A1 => n64808, A2 => n64809, A3 => n64810, A4 => 
                           n64811, ZN => n64807);
   U48783 : OAI221_X1 port map( B1 => n63147, B2 => n67627, C1 => n62276, C2 =>
                           n67621, A => n64813, ZN => n64810);
   U48784 : OAI221_X1 port map( B1 => n62475, B2 => n67603, C1 => n63552, C2 =>
                           n67597, A => n64814, ZN => n64809);
   U48785 : OAI221_X1 port map( B1 => n54233, B2 => n67579, C1 => n63618, C2 =>
                           n67573, A => n64816, ZN => n64808);
   U48786 : NOR4_X1 port map( A1 => n64788, A2 => n64789, A3 => n64790, A4 => 
                           n64791, ZN => n64787);
   U48787 : OAI221_X1 port map( B1 => n63146, B2 => n67627, C1 => n62275, C2 =>
                           n67621, A => n64793, ZN => n64790);
   U48788 : OAI221_X1 port map( B1 => n62474, B2 => n67603, C1 => n63551, C2 =>
                           n67597, A => n64794, ZN => n64789);
   U48789 : OAI221_X1 port map( B1 => n54232, B2 => n67579, C1 => n63617, C2 =>
                           n67573, A => n64796, ZN => n64788);
   U48790 : NOR4_X1 port map( A1 => n64768, A2 => n64769, A3 => n64770, A4 => 
                           n64771, ZN => n64767);
   U48791 : OAI221_X1 port map( B1 => n63145, B2 => n67627, C1 => n62274, C2 =>
                           n67621, A => n64773, ZN => n64770);
   U48792 : OAI221_X1 port map( B1 => n62473, B2 => n67603, C1 => n63550, C2 =>
                           n67597, A => n64774, ZN => n64769);
   U48793 : OAI221_X1 port map( B1 => n54231, B2 => n67579, C1 => n63616, C2 =>
                           n67573, A => n64776, ZN => n64768);
   U48794 : NOR4_X1 port map( A1 => n64748, A2 => n64749, A3 => n64750, A4 => 
                           n64751, ZN => n64747);
   U48795 : OAI221_X1 port map( B1 => n63144, B2 => n67627, C1 => n62273, C2 =>
                           n67621, A => n64753, ZN => n64750);
   U48796 : OAI221_X1 port map( B1 => n62472, B2 => n67603, C1 => n63549, C2 =>
                           n67597, A => n64754, ZN => n64749);
   U48797 : OAI221_X1 port map( B1 => n54230, B2 => n67579, C1 => n63615, C2 =>
                           n67573, A => n64756, ZN => n64748);
   U48798 : NOR4_X1 port map( A1 => n64728, A2 => n64729, A3 => n64730, A4 => 
                           n64731, ZN => n64727);
   U48799 : OAI221_X1 port map( B1 => n63143, B2 => n67627, C1 => n62272, C2 =>
                           n67621, A => n64733, ZN => n64730);
   U48800 : OAI221_X1 port map( B1 => n62471, B2 => n67603, C1 => n63548, C2 =>
                           n67597, A => n64734, ZN => n64729);
   U48801 : OAI221_X1 port map( B1 => n54229, B2 => n67579, C1 => n63614, C2 =>
                           n67573, A => n64736, ZN => n64728);
   U48802 : NOR4_X1 port map( A1 => n64708, A2 => n64709, A3 => n64710, A4 => 
                           n64711, ZN => n64707);
   U48803 : OAI221_X1 port map( B1 => n63142, B2 => n67627, C1 => n62271, C2 =>
                           n67621, A => n64713, ZN => n64710);
   U48804 : OAI221_X1 port map( B1 => n62470, B2 => n67603, C1 => n63547, C2 =>
                           n67597, A => n64714, ZN => n64709);
   U48805 : OAI221_X1 port map( B1 => n54228, B2 => n67579, C1 => n63613, C2 =>
                           n67573, A => n64716, ZN => n64708);
   U48806 : NOR4_X1 port map( A1 => n64688, A2 => n64689, A3 => n64690, A4 => 
                           n64691, ZN => n64687);
   U48807 : OAI221_X1 port map( B1 => n63141, B2 => n67627, C1 => n62270, C2 =>
                           n67621, A => n64693, ZN => n64690);
   U48808 : OAI221_X1 port map( B1 => n62469, B2 => n67603, C1 => n63546, C2 =>
                           n67597, A => n64694, ZN => n64689);
   U48809 : OAI221_X1 port map( B1 => n54227, B2 => n67579, C1 => n63612, C2 =>
                           n67573, A => n64696, ZN => n64688);
   U48810 : NOR4_X1 port map( A1 => n64668, A2 => n64669, A3 => n64670, A4 => 
                           n64671, ZN => n64667);
   U48811 : OAI221_X1 port map( B1 => n63140, B2 => n67627, C1 => n62269, C2 =>
                           n67621, A => n64673, ZN => n64670);
   U48812 : OAI221_X1 port map( B1 => n62468, B2 => n67603, C1 => n63545, C2 =>
                           n67597, A => n64674, ZN => n64669);
   U48813 : OAI221_X1 port map( B1 => n54226, B2 => n67579, C1 => n63611, C2 =>
                           n67573, A => n64676, ZN => n64668);
   U48814 : NOR4_X1 port map( A1 => n64648, A2 => n64649, A3 => n64650, A4 => 
                           n64651, ZN => n64647);
   U48815 : OAI221_X1 port map( B1 => n63139, B2 => n67627, C1 => n62268, C2 =>
                           n67621, A => n64653, ZN => n64650);
   U48816 : OAI221_X1 port map( B1 => n62467, B2 => n67603, C1 => n63544, C2 =>
                           n67597, A => n64654, ZN => n64649);
   U48817 : OAI221_X1 port map( B1 => n54225, B2 => n67579, C1 => n63610, C2 =>
                           n67573, A => n64656, ZN => n64648);
   U48818 : NOR4_X1 port map( A1 => n64628, A2 => n64629, A3 => n64630, A4 => 
                           n64631, ZN => n64627);
   U48819 : OAI221_X1 port map( B1 => n63138, B2 => n67627, C1 => n62267, C2 =>
                           n67621, A => n64633, ZN => n64630);
   U48820 : OAI221_X1 port map( B1 => n62466, B2 => n67603, C1 => n63543, C2 =>
                           n67597, A => n64634, ZN => n64629);
   U48821 : OAI221_X1 port map( B1 => n54224, B2 => n67579, C1 => n63609, C2 =>
                           n67573, A => n64636, ZN => n64628);
   U48822 : NOR4_X1 port map( A1 => n64608, A2 => n64609, A3 => n64610, A4 => 
                           n64611, ZN => n64607);
   U48823 : OAI221_X1 port map( B1 => n63137, B2 => n67627, C1 => n62266, C2 =>
                           n67621, A => n64613, ZN => n64610);
   U48824 : OAI221_X1 port map( B1 => n62465, B2 => n67603, C1 => n63542, C2 =>
                           n67597, A => n64614, ZN => n64609);
   U48825 : OAI221_X1 port map( B1 => n54223, B2 => n67579, C1 => n63608, C2 =>
                           n67573, A => n64616, ZN => n64608);
   U48826 : NOR4_X1 port map( A1 => n64588, A2 => n64589, A3 => n64590, A4 => 
                           n64591, ZN => n64587);
   U48827 : OAI221_X1 port map( B1 => n63136, B2 => n67628, C1 => n62265, C2 =>
                           n67622, A => n64593, ZN => n64590);
   U48828 : OAI221_X1 port map( B1 => n62464, B2 => n67604, C1 => n63541, C2 =>
                           n67598, A => n64594, ZN => n64589);
   U48829 : OAI221_X1 port map( B1 => n54222, B2 => n67580, C1 => n63607, C2 =>
                           n67574, A => n64596, ZN => n64588);
   U48830 : NOR4_X1 port map( A1 => n64568, A2 => n64569, A3 => n64570, A4 => 
                           n64571, ZN => n64567);
   U48831 : OAI221_X1 port map( B1 => n63135, B2 => n67628, C1 => n62264, C2 =>
                           n67622, A => n64573, ZN => n64570);
   U48832 : OAI221_X1 port map( B1 => n62463, B2 => n67604, C1 => n63540, C2 =>
                           n67598, A => n64574, ZN => n64569);
   U48833 : OAI221_X1 port map( B1 => n54221, B2 => n67580, C1 => n63606, C2 =>
                           n67574, A => n64576, ZN => n64568);
   U48834 : NOR4_X1 port map( A1 => n64548, A2 => n64549, A3 => n64550, A4 => 
                           n64551, ZN => n64547);
   U48835 : OAI221_X1 port map( B1 => n63134, B2 => n67628, C1 => n62263, C2 =>
                           n67622, A => n64553, ZN => n64550);
   U48836 : OAI221_X1 port map( B1 => n62462, B2 => n67604, C1 => n63539, C2 =>
                           n67598, A => n64554, ZN => n64549);
   U48837 : OAI221_X1 port map( B1 => n54220, B2 => n67580, C1 => n63605, C2 =>
                           n67574, A => n64556, ZN => n64548);
   U48838 : NOR4_X1 port map( A1 => n64528, A2 => n64529, A3 => n64530, A4 => 
                           n64531, ZN => n64527);
   U48839 : OAI221_X1 port map( B1 => n63133, B2 => n67628, C1 => n62262, C2 =>
                           n67622, A => n64533, ZN => n64530);
   U48840 : OAI221_X1 port map( B1 => n62461, B2 => n67604, C1 => n63538, C2 =>
                           n67598, A => n64534, ZN => n64529);
   U48841 : OAI221_X1 port map( B1 => n54219, B2 => n67580, C1 => n63604, C2 =>
                           n67574, A => n64536, ZN => n64528);
   U48842 : NOR4_X1 port map( A1 => n64508, A2 => n64509, A3 => n64510, A4 => 
                           n64511, ZN => n64507);
   U48843 : OAI221_X1 port map( B1 => n63132, B2 => n67628, C1 => n62261, C2 =>
                           n67622, A => n64513, ZN => n64510);
   U48844 : OAI221_X1 port map( B1 => n62460, B2 => n67604, C1 => n63537, C2 =>
                           n67598, A => n64514, ZN => n64509);
   U48845 : OAI221_X1 port map( B1 => n54218, B2 => n67580, C1 => n63603, C2 =>
                           n67574, A => n64516, ZN => n64508);
   U48846 : NOR4_X1 port map( A1 => n64488, A2 => n64489, A3 => n64490, A4 => 
                           n64491, ZN => n64487);
   U48847 : OAI221_X1 port map( B1 => n63131, B2 => n67628, C1 => n62260, C2 =>
                           n67622, A => n64493, ZN => n64490);
   U48848 : OAI221_X1 port map( B1 => n62459, B2 => n67604, C1 => n63536, C2 =>
                           n67598, A => n64494, ZN => n64489);
   U48849 : OAI221_X1 port map( B1 => n54217, B2 => n67580, C1 => n63602, C2 =>
                           n67574, A => n64496, ZN => n64488);
   U48850 : NOR4_X1 port map( A1 => n64468, A2 => n64469, A3 => n64470, A4 => 
                           n64471, ZN => n64467);
   U48851 : OAI221_X1 port map( B1 => n63130, B2 => n67628, C1 => n62259, C2 =>
                           n67622, A => n64473, ZN => n64470);
   U48852 : OAI221_X1 port map( B1 => n62458, B2 => n67604, C1 => n63535, C2 =>
                           n67598, A => n64474, ZN => n64469);
   U48853 : OAI221_X1 port map( B1 => n54216, B2 => n67580, C1 => n63601, C2 =>
                           n67574, A => n64476, ZN => n64468);
   U48854 : NOR4_X1 port map( A1 => n64448, A2 => n64449, A3 => n64450, A4 => 
                           n64451, ZN => n64447);
   U48855 : OAI221_X1 port map( B1 => n63129, B2 => n67628, C1 => n62258, C2 =>
                           n67622, A => n64453, ZN => n64450);
   U48856 : OAI221_X1 port map( B1 => n62457, B2 => n67604, C1 => n63534, C2 =>
                           n67598, A => n64454, ZN => n64449);
   U48857 : OAI221_X1 port map( B1 => n54215, B2 => n67580, C1 => n63600, C2 =>
                           n67574, A => n64456, ZN => n64448);
   U48858 : NOR4_X1 port map( A1 => n64428, A2 => n64429, A3 => n64430, A4 => 
                           n64431, ZN => n64427);
   U48859 : OAI221_X1 port map( B1 => n63128, B2 => n67628, C1 => n62257, C2 =>
                           n67622, A => n64433, ZN => n64430);
   U48860 : OAI221_X1 port map( B1 => n62456, B2 => n67604, C1 => n63533, C2 =>
                           n67598, A => n64434, ZN => n64429);
   U48861 : OAI221_X1 port map( B1 => n54214, B2 => n67580, C1 => n63599, C2 =>
                           n67574, A => n64436, ZN => n64428);
   U48862 : NOR4_X1 port map( A1 => n64408, A2 => n64409, A3 => n64410, A4 => 
                           n64411, ZN => n64407);
   U48863 : OAI221_X1 port map( B1 => n63127, B2 => n67628, C1 => n62256, C2 =>
                           n67622, A => n64413, ZN => n64410);
   U48864 : OAI221_X1 port map( B1 => n62455, B2 => n67604, C1 => n63532, C2 =>
                           n67598, A => n64414, ZN => n64409);
   U48865 : OAI221_X1 port map( B1 => n54213, B2 => n67580, C1 => n63598, C2 =>
                           n67574, A => n64416, ZN => n64408);
   U48866 : NOR4_X1 port map( A1 => n64388, A2 => n64389, A3 => n64390, A4 => 
                           n64391, ZN => n64387);
   U48867 : OAI221_X1 port map( B1 => n63126, B2 => n67628, C1 => n62255, C2 =>
                           n67622, A => n64393, ZN => n64390);
   U48868 : OAI221_X1 port map( B1 => n62454, B2 => n67604, C1 => n63531, C2 =>
                           n67598, A => n64394, ZN => n64389);
   U48869 : OAI221_X1 port map( B1 => n54212, B2 => n67580, C1 => n63597, C2 =>
                           n67574, A => n64396, ZN => n64388);
   U48870 : NOR4_X1 port map( A1 => n64368, A2 => n64369, A3 => n64370, A4 => 
                           n64371, ZN => n64367);
   U48871 : OAI221_X1 port map( B1 => n63125, B2 => n67628, C1 => n62254, C2 =>
                           n67622, A => n64373, ZN => n64370);
   U48872 : OAI221_X1 port map( B1 => n62453, B2 => n67604, C1 => n63530, C2 =>
                           n67598, A => n64374, ZN => n64369);
   U48873 : OAI221_X1 port map( B1 => n54211, B2 => n67580, C1 => n63596, C2 =>
                           n67574, A => n64376, ZN => n64368);
   U48874 : NOR4_X1 port map( A1 => n64348, A2 => n64349, A3 => n64350, A4 => 
                           n64351, ZN => n64347);
   U48875 : OAI221_X1 port map( B1 => n63124, B2 => n67629, C1 => n62253, C2 =>
                           n67623, A => n64353, ZN => n64350);
   U48876 : OAI221_X1 port map( B1 => n62452, B2 => n67605, C1 => n63529, C2 =>
                           n67599, A => n64354, ZN => n64349);
   U48877 : OAI221_X1 port map( B1 => n54210, B2 => n67581, C1 => n63595, C2 =>
                           n67575, A => n64356, ZN => n64348);
   U48878 : NOR4_X1 port map( A1 => n64328, A2 => n64329, A3 => n64330, A4 => 
                           n64331, ZN => n64327);
   U48879 : OAI221_X1 port map( B1 => n63123, B2 => n67629, C1 => n62252, C2 =>
                           n67623, A => n64333, ZN => n64330);
   U48880 : OAI221_X1 port map( B1 => n62451, B2 => n67605, C1 => n63528, C2 =>
                           n67599, A => n64334, ZN => n64329);
   U48881 : OAI221_X1 port map( B1 => n54209, B2 => n67581, C1 => n63594, C2 =>
                           n67575, A => n64336, ZN => n64328);
   U48882 : NOR4_X1 port map( A1 => n64308, A2 => n64309, A3 => n64310, A4 => 
                           n64311, ZN => n64307);
   U48883 : OAI221_X1 port map( B1 => n63122, B2 => n67629, C1 => n62251, C2 =>
                           n67623, A => n64313, ZN => n64310);
   U48884 : OAI221_X1 port map( B1 => n62450, B2 => n67605, C1 => n63527, C2 =>
                           n67599, A => n64314, ZN => n64309);
   U48885 : OAI221_X1 port map( B1 => n54208, B2 => n67581, C1 => n63593, C2 =>
                           n67575, A => n64316, ZN => n64308);
   U48886 : NOR4_X1 port map( A1 => n64288, A2 => n64289, A3 => n64290, A4 => 
                           n64291, ZN => n64287);
   U48887 : OAI221_X1 port map( B1 => n63121, B2 => n67629, C1 => n62250, C2 =>
                           n67623, A => n64293, ZN => n64290);
   U48888 : OAI221_X1 port map( B1 => n62449, B2 => n67605, C1 => n63526, C2 =>
                           n67599, A => n64294, ZN => n64289);
   U48889 : OAI221_X1 port map( B1 => n54207, B2 => n67581, C1 => n63592, C2 =>
                           n67575, A => n64296, ZN => n64288);
   U48890 : NOR4_X1 port map( A1 => n64268, A2 => n64269, A3 => n64270, A4 => 
                           n64271, ZN => n64267);
   U48891 : OAI221_X1 port map( B1 => n63120, B2 => n67629, C1 => n62249, C2 =>
                           n67623, A => n64273, ZN => n64270);
   U48892 : OAI221_X1 port map( B1 => n62448, B2 => n67605, C1 => n63525, C2 =>
                           n67599, A => n64274, ZN => n64269);
   U48893 : OAI221_X1 port map( B1 => n54206, B2 => n67581, C1 => n63591, C2 =>
                           n67575, A => n64276, ZN => n64268);
   U48894 : NOR4_X1 port map( A1 => n64248, A2 => n64249, A3 => n64250, A4 => 
                           n64251, ZN => n64247);
   U48895 : OAI221_X1 port map( B1 => n63119, B2 => n67629, C1 => n62248, C2 =>
                           n67623, A => n64253, ZN => n64250);
   U48896 : OAI221_X1 port map( B1 => n62447, B2 => n67605, C1 => n63524, C2 =>
                           n67599, A => n64254, ZN => n64249);
   U48897 : OAI221_X1 port map( B1 => n54205, B2 => n67581, C1 => n63590, C2 =>
                           n67575, A => n64256, ZN => n64248);
   U48898 : NOR4_X1 port map( A1 => n64228, A2 => n64229, A3 => n64230, A4 => 
                           n64231, ZN => n64227);
   U48899 : OAI221_X1 port map( B1 => n63118, B2 => n67629, C1 => n62247, C2 =>
                           n67623, A => n64233, ZN => n64230);
   U48900 : OAI221_X1 port map( B1 => n62446, B2 => n67605, C1 => n63523, C2 =>
                           n67599, A => n64234, ZN => n64229);
   U48901 : OAI221_X1 port map( B1 => n54204, B2 => n67581, C1 => n63589, C2 =>
                           n67575, A => n64236, ZN => n64228);
   U48902 : NOR4_X1 port map( A1 => n64208, A2 => n64209, A3 => n64210, A4 => 
                           n64211, ZN => n64207);
   U48903 : OAI221_X1 port map( B1 => n63117, B2 => n67629, C1 => n62246, C2 =>
                           n67623, A => n64213, ZN => n64210);
   U48904 : OAI221_X1 port map( B1 => n62445, B2 => n67605, C1 => n63522, C2 =>
                           n67599, A => n64214, ZN => n64209);
   U48905 : OAI221_X1 port map( B1 => n54203, B2 => n67581, C1 => n63588, C2 =>
                           n67575, A => n64216, ZN => n64208);
   U48906 : NOR4_X1 port map( A1 => n64188, A2 => n64189, A3 => n64190, A4 => 
                           n64191, ZN => n64187);
   U48907 : OAI221_X1 port map( B1 => n63116, B2 => n67629, C1 => n62245, C2 =>
                           n67623, A => n64193, ZN => n64190);
   U48908 : OAI221_X1 port map( B1 => n62444, B2 => n67605, C1 => n63521, C2 =>
                           n67599, A => n64194, ZN => n64189);
   U48909 : OAI221_X1 port map( B1 => n54202, B2 => n67581, C1 => n63587, C2 =>
                           n67575, A => n64196, ZN => n64188);
   U48910 : NOR4_X1 port map( A1 => n64168, A2 => n64169, A3 => n64170, A4 => 
                           n64171, ZN => n64167);
   U48911 : OAI221_X1 port map( B1 => n63115, B2 => n67629, C1 => n62244, C2 =>
                           n67623, A => n64173, ZN => n64170);
   U48912 : OAI221_X1 port map( B1 => n62443, B2 => n67605, C1 => n63520, C2 =>
                           n67599, A => n64174, ZN => n64169);
   U48913 : OAI221_X1 port map( B1 => n54201, B2 => n67581, C1 => n63586, C2 =>
                           n67575, A => n64176, ZN => n64168);
   U48914 : NOR4_X1 port map( A1 => n64148, A2 => n64149, A3 => n64150, A4 => 
                           n64151, ZN => n64147);
   U48915 : OAI221_X1 port map( B1 => n63114, B2 => n67629, C1 => n62243, C2 =>
                           n67623, A => n64153, ZN => n64150);
   U48916 : OAI221_X1 port map( B1 => n62442, B2 => n67605, C1 => n63519, C2 =>
                           n67599, A => n64154, ZN => n64149);
   U48917 : OAI221_X1 port map( B1 => n54200, B2 => n67581, C1 => n63585, C2 =>
                           n67575, A => n64156, ZN => n64148);
   U48918 : NOR4_X1 port map( A1 => n64128, A2 => n64129, A3 => n64130, A4 => 
                           n64131, ZN => n64127);
   U48919 : OAI221_X1 port map( B1 => n63113, B2 => n67629, C1 => n62242, C2 =>
                           n67623, A => n64133, ZN => n64130);
   U48920 : OAI221_X1 port map( B1 => n62441, B2 => n67605, C1 => n63518, C2 =>
                           n67599, A => n64134, ZN => n64129);
   U48921 : OAI221_X1 port map( B1 => n54199, B2 => n67581, C1 => n63584, C2 =>
                           n67575, A => n64136, ZN => n64128);
   U48922 : NOR4_X1 port map( A1 => n64108, A2 => n64109, A3 => n64110, A4 => 
                           n64111, ZN => n64107);
   U48923 : OAI221_X1 port map( B1 => n63112, B2 => n67630, C1 => n62241, C2 =>
                           n67624, A => n64113, ZN => n64110);
   U48924 : OAI221_X1 port map( B1 => n62440, B2 => n67606, C1 => n63517, C2 =>
                           n67600, A => n64114, ZN => n64109);
   U48925 : OAI221_X1 port map( B1 => n54198, B2 => n67582, C1 => n63583, C2 =>
                           n67576, A => n64116, ZN => n64108);
   U48926 : NOR4_X1 port map( A1 => n64088, A2 => n64089, A3 => n64090, A4 => 
                           n64091, ZN => n64087);
   U48927 : OAI221_X1 port map( B1 => n63111, B2 => n67630, C1 => n62240, C2 =>
                           n67624, A => n64093, ZN => n64090);
   U48928 : OAI221_X1 port map( B1 => n62439, B2 => n67606, C1 => n63516, C2 =>
                           n67600, A => n64094, ZN => n64089);
   U48929 : OAI221_X1 port map( B1 => n54197, B2 => n67582, C1 => n63582, C2 =>
                           n67576, A => n64096, ZN => n64088);
   U48930 : NOR4_X1 port map( A1 => n64068, A2 => n64069, A3 => n64070, A4 => 
                           n64071, ZN => n64067);
   U48931 : OAI221_X1 port map( B1 => n63110, B2 => n67630, C1 => n62239, C2 =>
                           n67624, A => n64073, ZN => n64070);
   U48932 : OAI221_X1 port map( B1 => n62438, B2 => n67606, C1 => n63515, C2 =>
                           n67600, A => n64074, ZN => n64069);
   U48933 : OAI221_X1 port map( B1 => n54196, B2 => n67582, C1 => n63581, C2 =>
                           n67576, A => n64076, ZN => n64068);
   U48934 : NOR4_X1 port map( A1 => n64048, A2 => n64049, A3 => n64050, A4 => 
                           n64051, ZN => n64047);
   U48935 : OAI221_X1 port map( B1 => n63109, B2 => n67630, C1 => n62238, C2 =>
                           n67624, A => n64053, ZN => n64050);
   U48936 : OAI221_X1 port map( B1 => n62437, B2 => n67606, C1 => n63514, C2 =>
                           n67600, A => n64054, ZN => n64049);
   U48937 : OAI221_X1 port map( B1 => n54195, B2 => n67582, C1 => n63580, C2 =>
                           n67576, A => n64056, ZN => n64048);
   U48938 : NOR4_X1 port map( A1 => n64028, A2 => n64029, A3 => n64030, A4 => 
                           n64031, ZN => n64027);
   U48939 : OAI221_X1 port map( B1 => n63108, B2 => n67630, C1 => n62237, C2 =>
                           n67624, A => n64033, ZN => n64030);
   U48940 : OAI221_X1 port map( B1 => n62436, B2 => n67606, C1 => n63513, C2 =>
                           n67600, A => n64034, ZN => n64029);
   U48941 : OAI221_X1 port map( B1 => n54194, B2 => n67582, C1 => n63579, C2 =>
                           n67576, A => n64036, ZN => n64028);
   U48942 : NOR4_X1 port map( A1 => n64008, A2 => n64009, A3 => n64010, A4 => 
                           n64011, ZN => n64007);
   U48943 : OAI221_X1 port map( B1 => n63107, B2 => n67630, C1 => n62236, C2 =>
                           n67624, A => n64013, ZN => n64010);
   U48944 : OAI221_X1 port map( B1 => n62435, B2 => n67606, C1 => n63512, C2 =>
                           n67600, A => n64014, ZN => n64009);
   U48945 : OAI221_X1 port map( B1 => n54193, B2 => n67582, C1 => n63578, C2 =>
                           n67576, A => n64016, ZN => n64008);
   U48946 : NOR4_X1 port map( A1 => n63988, A2 => n63989, A3 => n63990, A4 => 
                           n63991, ZN => n63987);
   U48947 : OAI221_X1 port map( B1 => n63106, B2 => n67630, C1 => n62235, C2 =>
                           n67624, A => n63993, ZN => n63990);
   U48948 : OAI221_X1 port map( B1 => n62434, B2 => n67606, C1 => n63511, C2 =>
                           n67600, A => n63994, ZN => n63989);
   U48949 : OAI221_X1 port map( B1 => n54192, B2 => n67582, C1 => n63577, C2 =>
                           n67576, A => n63996, ZN => n63988);
   U48950 : NOR4_X1 port map( A1 => n63968, A2 => n63969, A3 => n63970, A4 => 
                           n63971, ZN => n63967);
   U48951 : OAI221_X1 port map( B1 => n63105, B2 => n67630, C1 => n62234, C2 =>
                           n67624, A => n63973, ZN => n63970);
   U48952 : OAI221_X1 port map( B1 => n62433, B2 => n67606, C1 => n63510, C2 =>
                           n67600, A => n63974, ZN => n63969);
   U48953 : OAI221_X1 port map( B1 => n54191, B2 => n67582, C1 => n63576, C2 =>
                           n67576, A => n63976, ZN => n63968);
   U48954 : NOR4_X1 port map( A1 => n63948, A2 => n63949, A3 => n63950, A4 => 
                           n63951, ZN => n63947);
   U48955 : OAI221_X1 port map( B1 => n63104, B2 => n67630, C1 => n62233, C2 =>
                           n67624, A => n63953, ZN => n63950);
   U48956 : OAI221_X1 port map( B1 => n62432, B2 => n67606, C1 => n63509, C2 =>
                           n67600, A => n63954, ZN => n63949);
   U48957 : OAI221_X1 port map( B1 => n54190, B2 => n67582, C1 => n63575, C2 =>
                           n67576, A => n63956, ZN => n63948);
   U48958 : NOR4_X1 port map( A1 => n63928, A2 => n63929, A3 => n63930, A4 => 
                           n63931, ZN => n63927);
   U48959 : OAI221_X1 port map( B1 => n63103, B2 => n67630, C1 => n62232, C2 =>
                           n67624, A => n63933, ZN => n63930);
   U48960 : OAI221_X1 port map( B1 => n62431, B2 => n67606, C1 => n63508, C2 =>
                           n67600, A => n63934, ZN => n63929);
   U48961 : OAI221_X1 port map( B1 => n54189, B2 => n67582, C1 => n63574, C2 =>
                           n67576, A => n63936, ZN => n63928);
   U48962 : NOR4_X1 port map( A1 => n63908, A2 => n63909, A3 => n63910, A4 => 
                           n63911, ZN => n63907);
   U48963 : OAI221_X1 port map( B1 => n63102, B2 => n67630, C1 => n62231, C2 =>
                           n67624, A => n63913, ZN => n63910);
   U48964 : OAI221_X1 port map( B1 => n62430, B2 => n67606, C1 => n63507, C2 =>
                           n67600, A => n63914, ZN => n63909);
   U48965 : OAI221_X1 port map( B1 => n54188, B2 => n67582, C1 => n63573, C2 =>
                           n67576, A => n63916, ZN => n63908);
   U48966 : NOR4_X1 port map( A1 => n63888, A2 => n63889, A3 => n63890, A4 => 
                           n63891, ZN => n63887);
   U48967 : OAI221_X1 port map( B1 => n63101, B2 => n67630, C1 => n62230, C2 =>
                           n67624, A => n63893, ZN => n63890);
   U48968 : OAI221_X1 port map( B1 => n62429, B2 => n67606, C1 => n63506, C2 =>
                           n67600, A => n63894, ZN => n63889);
   U48969 : OAI221_X1 port map( B1 => n54187, B2 => n67582, C1 => n63572, C2 =>
                           n67576, A => n63896, ZN => n63888);
   U48970 : NOR4_X1 port map( A1 => n63877, A2 => n63878, A3 => n63879, A4 => 
                           n63880, ZN => n63865);
   U48971 : OAI222_X1 port map( A1 => n63166, A2 => n67523, B1 => n62095, B2 =>
                           n67517, C1 => n62498, C2 => n67511, ZN => n63877);
   U48972 : OAI22_X1 port map( A1 => n8449, A2 => n67547, B1 => n62362, B2 => 
                           n67541, ZN => n63879);
   U48973 : OAI22_X1 port map( A1 => n62631, A2 => n67559, B1 => n54610, B2 => 
                           n67553, ZN => n63880);
   U48974 : NOR4_X1 port map( A1 => n63856, A2 => n63857, A3 => n63858, A4 => 
                           n63859, ZN => n63844);
   U48975 : OAI222_X1 port map( A1 => n63165, A2 => n67523, B1 => n62094, B2 =>
                           n67517, C1 => n62497, C2 => n67511, ZN => n63856);
   U48976 : OAI22_X1 port map( A1 => n8465, A2 => n67547, B1 => n62361, B2 => 
                           n67541, ZN => n63858);
   U48977 : OAI22_X1 port map( A1 => n62630, A2 => n67559, B1 => n54609, B2 => 
                           n67553, ZN => n63859);
   U48978 : NOR4_X1 port map( A1 => n63835, A2 => n63836, A3 => n63837, A4 => 
                           n63838, ZN => n63823);
   U48979 : OAI222_X1 port map( A1 => n63164, A2 => n67523, B1 => n62093, B2 =>
                           n67517, C1 => n62496, C2 => n67511, ZN => n63835);
   U48980 : OAI22_X1 port map( A1 => n8481, A2 => n67547, B1 => n62360, B2 => 
                           n67541, ZN => n63837);
   U48981 : OAI22_X1 port map( A1 => n62629, A2 => n67559, B1 => n54608, B2 => 
                           n67553, ZN => n63838);
   U48982 : NOR4_X1 port map( A1 => n63797, A2 => n63798, A3 => n63799, A4 => 
                           n63800, ZN => n63769);
   U48983 : OAI222_X1 port map( A1 => n63162, A2 => n67523, B1 => n62091, B2 =>
                           n67517, C1 => n62494, C2 => n67511, ZN => n63797);
   U48984 : OAI22_X1 port map( A1 => n8497, A2 => n67547, B1 => n62358, B2 => 
                           n67541, ZN => n63799);
   U48985 : OAI22_X1 port map( A1 => n62627, A2 => n67559, B1 => n54606, B2 => 
                           n67553, ZN => n63800);
   U48986 : AOI221_X1 port map( B1 => n67307, B2 => n58717, C1 => n67301, C2 =>
                           n58299, A => n65167, ZN => n65152);
   U48987 : OAI22_X1 port map( A1 => n62093, A2 => n67295, B1 => n62160, B2 => 
                           n67289, ZN => n65167);
   U48988 : AOI221_X1 port map( B1 => n67307, B2 => n58718, C1 => n67301, C2 =>
                           n58301, A => n65143, ZN => n65101);
   U48989 : OAI22_X1 port map( A1 => n62091, A2 => n67295, B1 => n62158, B2 => 
                           n67289, ZN => n65143);
   U48990 : AOI221_X1 port map( B1 => n67307, B2 => n58715, C1 => n67301, C2 =>
                           n58295, A => n65203, ZN => n65188);
   U48991 : OAI22_X1 port map( A1 => n62095, A2 => n67295, B1 => n62162, B2 => 
                           n67289, ZN => n65203);
   U48992 : AOI221_X1 port map( B1 => n67307, B2 => n58716, C1 => n67301, C2 =>
                           n58297, A => n65185, ZN => n65170);
   U48993 : OAI22_X1 port map( A1 => n62094, A2 => n67295, B1 => n62161, B2 => 
                           n67289, ZN => n65185);
   U48994 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), ZN => n62489);
   U48995 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => n63497, ZN => n62356);
   U48996 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n63496, ZN => n62223);
   U48997 : AND3_X1 port map( A1 => n66494, A2 => n65099, A3 => ADD_RD1(1), ZN 
                           => n65075);
   U48998 : OAI221_X1 port map( B1 => n63415, B2 => n67649, C1 => n49432, C2 =>
                           n67643, A => n64832, ZN => n64831);
   U48999 : AOI22_X1 port map( A1 => n67637, A2 => n57725, B1 => n67633, B2 => 
                           OUT1_12_port, ZN => n64832);
   U49000 : OAI221_X1 port map( B1 => n63414, B2 => n67649, C1 => n49433, C2 =>
                           n67643, A => n64812, ZN => n64811);
   U49001 : AOI22_X1 port map( A1 => n67637, A2 => n57701, B1 => n67635, B2 => 
                           OUT1_13_port, ZN => n64812);
   U49002 : OAI221_X1 port map( B1 => n63413, B2 => n67649, C1 => n49434, C2 =>
                           n67643, A => n64792, ZN => n64791);
   U49003 : AOI22_X1 port map( A1 => n67637, A2 => n57677, B1 => n67634, B2 => 
                           OUT1_14_port, ZN => n64792);
   U49004 : OAI221_X1 port map( B1 => n63412, B2 => n67649, C1 => n49435, C2 =>
                           n67643, A => n64772, ZN => n64771);
   U49005 : AOI22_X1 port map( A1 => n67637, A2 => n57653, B1 => n67633, B2 => 
                           OUT1_15_port, ZN => n64772);
   U49006 : OAI221_X1 port map( B1 => n63411, B2 => n67649, C1 => n49436, C2 =>
                           n67643, A => n64752, ZN => n64751);
   U49007 : AOI22_X1 port map( A1 => n67637, A2 => n57629, B1 => n67635, B2 => 
                           OUT1_16_port, ZN => n64752);
   U49008 : OAI221_X1 port map( B1 => n63410, B2 => n67649, C1 => n49437, C2 =>
                           n67643, A => n64732, ZN => n64731);
   U49009 : AOI22_X1 port map( A1 => n67637, A2 => n57605, B1 => n67634, B2 => 
                           OUT1_17_port, ZN => n64732);
   U49010 : OAI221_X1 port map( B1 => n63409, B2 => n67649, C1 => n49438, C2 =>
                           n67643, A => n64712, ZN => n64711);
   U49011 : AOI22_X1 port map( A1 => n67637, A2 => n57581, B1 => n67633, B2 => 
                           OUT1_18_port, ZN => n64712);
   U49012 : OAI221_X1 port map( B1 => n63408, B2 => n67649, C1 => n49439, C2 =>
                           n67643, A => n64692, ZN => n64691);
   U49013 : AOI22_X1 port map( A1 => n67637, A2 => n57557, B1 => n67635, B2 => 
                           OUT1_19_port, ZN => n64692);
   U49014 : OAI221_X1 port map( B1 => n63407, B2 => n67649, C1 => n49440, C2 =>
                           n67643, A => n64672, ZN => n64671);
   U49015 : AOI22_X1 port map( A1 => n67637, A2 => n57533, B1 => n67634, B2 => 
                           OUT1_20_port, ZN => n64672);
   U49016 : OAI221_X1 port map( B1 => n63406, B2 => n67649, C1 => n49441, C2 =>
                           n67643, A => n64652, ZN => n64651);
   U49017 : AOI22_X1 port map( A1 => n67637, A2 => n57509, B1 => n67633, B2 => 
                           OUT1_21_port, ZN => n64652);
   U49018 : OAI221_X1 port map( B1 => n63405, B2 => n67649, C1 => n49442, C2 =>
                           n67643, A => n64632, ZN => n64631);
   U49019 : AOI22_X1 port map( A1 => n67637, A2 => n57485, B1 => n67634, B2 => 
                           OUT1_22_port, ZN => n64632);
   U49020 : OAI221_X1 port map( B1 => n63404, B2 => n67649, C1 => n49443, C2 =>
                           n67643, A => n64612, ZN => n64611);
   U49021 : AOI22_X1 port map( A1 => n67637, A2 => n57461, B1 => n67633, B2 => 
                           OUT1_23_port, ZN => n64612);
   U49022 : OAI221_X1 port map( B1 => n63403, B2 => n67650, C1 => n49444, C2 =>
                           n67644, A => n64592, ZN => n64591);
   U49023 : AOI22_X1 port map( A1 => n67638, A2 => n57437, B1 => n67633, B2 => 
                           OUT1_24_port, ZN => n64592);
   U49024 : OAI221_X1 port map( B1 => n63402, B2 => n67650, C1 => n49445, C2 =>
                           n67644, A => n64572, ZN => n64571);
   U49025 : AOI22_X1 port map( A1 => n67638, A2 => n57413, B1 => n67633, B2 => 
                           OUT1_25_port, ZN => n64572);
   U49026 : OAI221_X1 port map( B1 => n63401, B2 => n67650, C1 => n49446, C2 =>
                           n67644, A => n64552, ZN => n64551);
   U49027 : AOI22_X1 port map( A1 => n67638, A2 => n57389, B1 => n67633, B2 => 
                           OUT1_26_port, ZN => n64552);
   U49028 : OAI221_X1 port map( B1 => n63400, B2 => n67650, C1 => n49447, C2 =>
                           n67644, A => n64532, ZN => n64531);
   U49029 : AOI22_X1 port map( A1 => n67638, A2 => n57365, B1 => n67633, B2 => 
                           OUT1_27_port, ZN => n64532);
   U49030 : OAI221_X1 port map( B1 => n63399, B2 => n67650, C1 => n49448, C2 =>
                           n67644, A => n64512, ZN => n64511);
   U49031 : AOI22_X1 port map( A1 => n67638, A2 => n57341, B1 => n67633, B2 => 
                           OUT1_28_port, ZN => n64512);
   U49032 : OAI221_X1 port map( B1 => n63398, B2 => n67650, C1 => n49449, C2 =>
                           n67644, A => n64492, ZN => n64491);
   U49033 : AOI22_X1 port map( A1 => n67638, A2 => n57317, B1 => n67633, B2 => 
                           OUT1_29_port, ZN => n64492);
   U49034 : OAI221_X1 port map( B1 => n63397, B2 => n67650, C1 => n49450, C2 =>
                           n67644, A => n64472, ZN => n64471);
   U49035 : AOI22_X1 port map( A1 => n67638, A2 => n57293, B1 => n67633, B2 => 
                           OUT1_30_port, ZN => n64472);
   U49036 : OAI221_X1 port map( B1 => n63396, B2 => n67650, C1 => n49451, C2 =>
                           n67644, A => n64452, ZN => n64451);
   U49037 : AOI22_X1 port map( A1 => n67638, A2 => n57269, B1 => n67633, B2 => 
                           OUT1_31_port, ZN => n64452);
   U49038 : OAI221_X1 port map( B1 => n63395, B2 => n67650, C1 => n49452, C2 =>
                           n67644, A => n64432, ZN => n64431);
   U49039 : AOI22_X1 port map( A1 => n67638, A2 => n57245, B1 => n67633, B2 => 
                           OUT1_32_port, ZN => n64432);
   U49040 : OAI221_X1 port map( B1 => n63394, B2 => n67650, C1 => n49453, C2 =>
                           n67644, A => n64412, ZN => n64411);
   U49041 : AOI22_X1 port map( A1 => n67638, A2 => n57221, B1 => n67633, B2 => 
                           OUT1_33_port, ZN => n64412);
   U49042 : OAI221_X1 port map( B1 => n63393, B2 => n67650, C1 => n49454, C2 =>
                           n67644, A => n64392, ZN => n64391);
   U49043 : AOI22_X1 port map( A1 => n67638, A2 => n57197, B1 => n67633, B2 => 
                           OUT1_34_port, ZN => n64392);
   U49044 : OAI221_X1 port map( B1 => n63392, B2 => n67650, C1 => n49455, C2 =>
                           n67644, A => n64372, ZN => n64371);
   U49045 : AOI22_X1 port map( A1 => n67638, A2 => n57173, B1 => n67633, B2 => 
                           OUT1_35_port, ZN => n64372);
   U49046 : OAI221_X1 port map( B1 => n63391, B2 => n67651, C1 => n49456, C2 =>
                           n67645, A => n64352, ZN => n64351);
   U49047 : AOI22_X1 port map( A1 => n67639, A2 => n57149, B1 => n67633, B2 => 
                           OUT1_36_port, ZN => n64352);
   U49048 : OAI221_X1 port map( B1 => n63390, B2 => n67651, C1 => n49457, C2 =>
                           n67645, A => n64332, ZN => n64331);
   U49049 : AOI22_X1 port map( A1 => n67639, A2 => n57125, B1 => n67634, B2 => 
                           OUT1_37_port, ZN => n64332);
   U49050 : OAI221_X1 port map( B1 => n63389, B2 => n67651, C1 => n49458, C2 =>
                           n67645, A => n64312, ZN => n64311);
   U49051 : AOI22_X1 port map( A1 => n67639, A2 => n57101, B1 => n67634, B2 => 
                           OUT1_38_port, ZN => n64312);
   U49052 : OAI221_X1 port map( B1 => n63388, B2 => n67651, C1 => n49459, C2 =>
                           n67645, A => n64292, ZN => n64291);
   U49053 : AOI22_X1 port map( A1 => n67639, A2 => n57077, B1 => n67634, B2 => 
                           OUT1_39_port, ZN => n64292);
   U49054 : OAI221_X1 port map( B1 => n63387, B2 => n67651, C1 => n49460, C2 =>
                           n67645, A => n64272, ZN => n64271);
   U49055 : AOI22_X1 port map( A1 => n67639, A2 => n57053, B1 => n67634, B2 => 
                           OUT1_40_port, ZN => n64272);
   U49056 : OAI221_X1 port map( B1 => n63386, B2 => n67651, C1 => n49461, C2 =>
                           n67645, A => n64252, ZN => n64251);
   U49057 : AOI22_X1 port map( A1 => n67639, A2 => n57029, B1 => n67634, B2 => 
                           OUT1_41_port, ZN => n64252);
   U49058 : OAI221_X1 port map( B1 => n63385, B2 => n67651, C1 => n49462, C2 =>
                           n67645, A => n64232, ZN => n64231);
   U49059 : AOI22_X1 port map( A1 => n67639, A2 => n57005, B1 => n67634, B2 => 
                           OUT1_42_port, ZN => n64232);
   U49060 : OAI221_X1 port map( B1 => n63384, B2 => n67651, C1 => n49463, C2 =>
                           n67645, A => n64212, ZN => n64211);
   U49061 : AOI22_X1 port map( A1 => n67639, A2 => n56981, B1 => n67634, B2 => 
                           OUT1_43_port, ZN => n64212);
   U49062 : OAI221_X1 port map( B1 => n63383, B2 => n67651, C1 => n49464, C2 =>
                           n67645, A => n64192, ZN => n64191);
   U49063 : AOI22_X1 port map( A1 => n67639, A2 => n56957, B1 => n67634, B2 => 
                           OUT1_44_port, ZN => n64192);
   U49064 : OAI221_X1 port map( B1 => n63382, B2 => n67651, C1 => n49465, C2 =>
                           n67645, A => n64172, ZN => n64171);
   U49065 : AOI22_X1 port map( A1 => n67639, A2 => n56933, B1 => n67634, B2 => 
                           OUT1_45_port, ZN => n64172);
   U49066 : OAI221_X1 port map( B1 => n63381, B2 => n67651, C1 => n49466, C2 =>
                           n67645, A => n64152, ZN => n64151);
   U49067 : AOI22_X1 port map( A1 => n67639, A2 => n56909, B1 => n67634, B2 => 
                           OUT1_46_port, ZN => n64152);
   U49068 : OAI221_X1 port map( B1 => n63380, B2 => n67651, C1 => n49467, C2 =>
                           n67645, A => n64132, ZN => n64131);
   U49069 : AOI22_X1 port map( A1 => n67639, A2 => n56885, B1 => n67634, B2 => 
                           OUT1_47_port, ZN => n64132);
   U49070 : OAI221_X1 port map( B1 => n63379, B2 => n67652, C1 => n49468, C2 =>
                           n67646, A => n64112, ZN => n64111);
   U49071 : AOI22_X1 port map( A1 => n67640, A2 => n56861, B1 => n67634, B2 => 
                           OUT1_48_port, ZN => n64112);
   U49072 : OAI221_X1 port map( B1 => n63378, B2 => n67652, C1 => n49469, C2 =>
                           n67646, A => n64092, ZN => n64091);
   U49073 : AOI22_X1 port map( A1 => n67640, A2 => n56837, B1 => n67634, B2 => 
                           OUT1_49_port, ZN => n64092);
   U49074 : OAI221_X1 port map( B1 => n63377, B2 => n67652, C1 => n49470, C2 =>
                           n67646, A => n64072, ZN => n64071);
   U49075 : AOI22_X1 port map( A1 => n67640, A2 => n56813, B1 => n67635, B2 => 
                           OUT1_50_port, ZN => n64072);
   U49076 : OAI221_X1 port map( B1 => n63376, B2 => n67652, C1 => n49471, C2 =>
                           n67646, A => n64052, ZN => n64051);
   U49077 : AOI22_X1 port map( A1 => n67640, A2 => n56789, B1 => n67635, B2 => 
                           OUT1_51_port, ZN => n64052);
   U49078 : OAI221_X1 port map( B1 => n63375, B2 => n67652, C1 => n49472, C2 =>
                           n67646, A => n64032, ZN => n64031);
   U49079 : AOI22_X1 port map( A1 => n67640, A2 => n56765, B1 => n67635, B2 => 
                           OUT1_52_port, ZN => n64032);
   U49080 : OAI221_X1 port map( B1 => n63374, B2 => n67652, C1 => n49473, C2 =>
                           n67646, A => n64012, ZN => n64011);
   U49081 : AOI22_X1 port map( A1 => n67640, A2 => n56741, B1 => n67635, B2 => 
                           OUT1_53_port, ZN => n64012);
   U49082 : OAI221_X1 port map( B1 => n63373, B2 => n67652, C1 => n49474, C2 =>
                           n67646, A => n63992, ZN => n63991);
   U49083 : AOI22_X1 port map( A1 => n67640, A2 => n56717, B1 => n67635, B2 => 
                           OUT1_54_port, ZN => n63992);
   U49084 : OAI221_X1 port map( B1 => n63372, B2 => n67652, C1 => n49475, C2 =>
                           n67646, A => n63972, ZN => n63971);
   U49085 : AOI22_X1 port map( A1 => n67640, A2 => n56693, B1 => n67635, B2 => 
                           OUT1_55_port, ZN => n63972);
   U49086 : OAI221_X1 port map( B1 => n63371, B2 => n67652, C1 => n49476, C2 =>
                           n67646, A => n63952, ZN => n63951);
   U49087 : AOI22_X1 port map( A1 => n67640, A2 => n56669, B1 => n67635, B2 => 
                           OUT1_56_port, ZN => n63952);
   U49088 : OAI221_X1 port map( B1 => n63370, B2 => n67652, C1 => n49477, C2 =>
                           n67646, A => n63932, ZN => n63931);
   U49089 : AOI22_X1 port map( A1 => n67640, A2 => n56645, B1 => n67635, B2 => 
                           OUT1_57_port, ZN => n63932);
   U49090 : OAI221_X1 port map( B1 => n63369, B2 => n67652, C1 => n49478, C2 =>
                           n67646, A => n63912, ZN => n63911);
   U49091 : AOI22_X1 port map( A1 => n67640, A2 => n56621, B1 => n67635, B2 => 
                           OUT1_58_port, ZN => n63912);
   U49092 : OAI221_X1 port map( B1 => n63368, B2 => n67652, C1 => n49479, C2 =>
                           n67646, A => n63892, ZN => n63891);
   U49093 : AOI22_X1 port map( A1 => n67640, A2 => n56597, B1 => n67635, B2 => 
                           OUT1_59_port, ZN => n63892);
   U49094 : OAI221_X1 port map( B1 => n63365, B2 => n67457, C1 => n49231, C2 =>
                           n67451, A => n65159, ZN => n65158);
   U49095 : AOI22_X1 port map( A1 => n67445, A2 => n58377, B1 => n67439, B2 => 
                           OUT2_62_port, ZN => n65159);
   U49096 : OAI221_X1 port map( B1 => n63363, B2 => n67457, C1 => n49228, C2 =>
                           n67451, A => n65110, ZN => n65107);
   U49097 : AOI22_X1 port map( A1 => n67445, A2 => n58378, B1 => n67439, B2 => 
                           OUT2_63_port, ZN => n65110);
   U49098 : OAI221_X1 port map( B1 => n63367, B2 => n67457, C1 => n49229, C2 =>
                           n67451, A => n65195, ZN => n65194);
   U49099 : AOI22_X1 port map( A1 => n67445, A2 => n58375, B1 => n67438, B2 => 
                           OUT2_60_port, ZN => n65195);
   U49100 : OAI221_X1 port map( B1 => n63366, B2 => n67457, C1 => n49230, C2 =>
                           n67451, A => n65177, ZN => n65176);
   U49101 : AOI22_X1 port map( A1 => n67445, A2 => n58376, B1 => n67439, B2 => 
                           OUT2_61_port, ZN => n65177);
   U49102 : OAI221_X1 port map( B1 => n63367, B2 => n67653, C1 => n49480, C2 =>
                           n67647, A => n63871, ZN => n63870);
   U49103 : AOI22_X1 port map( A1 => n67641, A2 => n58784, B1 => n67635, B2 => 
                           OUT1_60_port, ZN => n63871);
   U49104 : OAI221_X1 port map( B1 => n63366, B2 => n67653, C1 => n49481, C2 =>
                           n67647, A => n63850, ZN => n63849);
   U49105 : AOI22_X1 port map( A1 => n67641, A2 => n58785, B1 => n67635, B2 => 
                           OUT1_61_port, ZN => n63850);
   U49106 : OAI221_X1 port map( B1 => n63365, B2 => n67653, C1 => n49482, C2 =>
                           n67647, A => n63829, ZN => n63828);
   U49107 : AOI22_X1 port map( A1 => n67641, A2 => n58786, B1 => n67635, B2 => 
                           OUT1_62_port, ZN => n63829);
   U49108 : OAI221_X1 port map( B1 => n63363, B2 => n67653, C1 => n49483, C2 =>
                           n67647, A => n63777, ZN => n63774);
   U49109 : AOI22_X1 port map( A1 => n67641, A2 => n58783, B1 => n67635, B2 => 
                           OUT1_63_port, ZN => n63777);
   U49110 : OAI221_X1 port map( B1 => n54658, B2 => n67429, C1 => n63553, C2 =>
                           n67423, A => n66060, ZN => n66057);
   U49111 : AOI22_X1 port map( A1 => n67417, A2 => n66325, B1 => n67411, B2 => 
                           n58319, ZN => n66060);
   U49112 : OAI221_X1 port map( B1 => n54657, B2 => n67429, C1 => n63552, C2 =>
                           n67423, A => n66042, ZN => n66039);
   U49113 : AOI22_X1 port map( A1 => n67417, A2 => n66326, B1 => n67411, B2 => 
                           n58320, ZN => n66042);
   U49114 : OAI221_X1 port map( B1 => n54656, B2 => n67429, C1 => n63551, C2 =>
                           n67423, A => n66024, ZN => n66021);
   U49115 : AOI22_X1 port map( A1 => n67417, A2 => n66327, B1 => n67411, B2 => 
                           n58321, ZN => n66024);
   U49116 : OAI221_X1 port map( B1 => n54655, B2 => n67429, C1 => n63550, C2 =>
                           n67423, A => n66006, ZN => n66003);
   U49117 : AOI22_X1 port map( A1 => n67417, A2 => n66328, B1 => n67411, B2 => 
                           n58322, ZN => n66006);
   U49118 : OAI221_X1 port map( B1 => n54654, B2 => n67429, C1 => n63549, C2 =>
                           n67423, A => n65988, ZN => n65985);
   U49119 : AOI22_X1 port map( A1 => n67417, A2 => n66329, B1 => n67411, B2 => 
                           n58323, ZN => n65988);
   U49120 : OAI221_X1 port map( B1 => n54653, B2 => n67429, C1 => n63548, C2 =>
                           n67423, A => n65970, ZN => n65967);
   U49121 : AOI22_X1 port map( A1 => n67417, A2 => n66330, B1 => n67411, B2 => 
                           n58324, ZN => n65970);
   U49122 : OAI221_X1 port map( B1 => n54652, B2 => n67429, C1 => n63547, C2 =>
                           n67423, A => n65952, ZN => n65949);
   U49123 : AOI22_X1 port map( A1 => n67417, A2 => n66331, B1 => n67411, B2 => 
                           n58325, ZN => n65952);
   U49124 : OAI221_X1 port map( B1 => n54651, B2 => n67429, C1 => n63546, C2 =>
                           n67423, A => n65934, ZN => n65931);
   U49125 : AOI22_X1 port map( A1 => n67417, A2 => n66332, B1 => n67411, B2 => 
                           n58326, ZN => n65934);
   U49126 : OAI221_X1 port map( B1 => n54650, B2 => n67429, C1 => n63545, C2 =>
                           n67423, A => n65916, ZN => n65913);
   U49127 : AOI22_X1 port map( A1 => n67417, A2 => n66333, B1 => n67411, B2 => 
                           n58327, ZN => n65916);
   U49128 : OAI221_X1 port map( B1 => n54649, B2 => n67429, C1 => n63544, C2 =>
                           n67423, A => n65898, ZN => n65895);
   U49129 : AOI22_X1 port map( A1 => n67417, A2 => n66334, B1 => n67411, B2 => 
                           n58328, ZN => n65898);
   U49130 : OAI221_X1 port map( B1 => n54648, B2 => n67429, C1 => n63543, C2 =>
                           n67423, A => n65880, ZN => n65877);
   U49131 : AOI22_X1 port map( A1 => n67417, A2 => n66335, B1 => n67411, B2 => 
                           n58329, ZN => n65880);
   U49132 : OAI221_X1 port map( B1 => n54647, B2 => n67429, C1 => n63542, C2 =>
                           n67423, A => n65862, ZN => n65859);
   U49133 : AOI22_X1 port map( A1 => n67417, A2 => n66336, B1 => n67411, B2 => 
                           n58330, ZN => n65862);
   U49134 : OAI221_X1 port map( B1 => n54646, B2 => n67430, C1 => n63541, C2 =>
                           n67424, A => n65844, ZN => n65841);
   U49135 : AOI22_X1 port map( A1 => n67418, A2 => n66337, B1 => n67412, B2 => 
                           n58331, ZN => n65844);
   U49136 : OAI221_X1 port map( B1 => n54645, B2 => n67430, C1 => n63540, C2 =>
                           n67424, A => n65826, ZN => n65823);
   U49137 : AOI22_X1 port map( A1 => n67418, A2 => n66338, B1 => n67412, B2 => 
                           n58332, ZN => n65826);
   U49138 : OAI221_X1 port map( B1 => n54644, B2 => n67430, C1 => n63539, C2 =>
                           n67424, A => n65808, ZN => n65805);
   U49139 : AOI22_X1 port map( A1 => n67418, A2 => n66339, B1 => n67412, B2 => 
                           n58333, ZN => n65808);
   U49140 : OAI221_X1 port map( B1 => n54643, B2 => n67430, C1 => n63538, C2 =>
                           n67424, A => n65790, ZN => n65787);
   U49141 : AOI22_X1 port map( A1 => n67418, A2 => n66340, B1 => n67412, B2 => 
                           n58334, ZN => n65790);
   U49142 : OAI221_X1 port map( B1 => n54642, B2 => n67430, C1 => n63537, C2 =>
                           n67424, A => n65772, ZN => n65769);
   U49143 : AOI22_X1 port map( A1 => n67418, A2 => n66341, B1 => n67412, B2 => 
                           n58335, ZN => n65772);
   U49144 : OAI221_X1 port map( B1 => n54641, B2 => n67430, C1 => n63536, C2 =>
                           n67424, A => n65754, ZN => n65751);
   U49145 : AOI22_X1 port map( A1 => n67418, A2 => n66342, B1 => n67412, B2 => 
                           n58336, ZN => n65754);
   U49146 : OAI221_X1 port map( B1 => n54640, B2 => n67430, C1 => n63535, C2 =>
                           n67424, A => n65736, ZN => n65733);
   U49147 : AOI22_X1 port map( A1 => n67418, A2 => n66343, B1 => n67412, B2 => 
                           n58337, ZN => n65736);
   U49148 : OAI221_X1 port map( B1 => n54639, B2 => n67430, C1 => n63534, C2 =>
                           n67424, A => n65718, ZN => n65715);
   U49149 : AOI22_X1 port map( A1 => n67418, A2 => n66344, B1 => n67412, B2 => 
                           n58338, ZN => n65718);
   U49150 : OAI221_X1 port map( B1 => n54638, B2 => n67430, C1 => n63533, C2 =>
                           n67424, A => n65700, ZN => n65697);
   U49151 : AOI22_X1 port map( A1 => n67418, A2 => n66345, B1 => n67412, B2 => 
                           n58339, ZN => n65700);
   U49152 : OAI221_X1 port map( B1 => n54637, B2 => n67430, C1 => n63532, C2 =>
                           n67424, A => n65682, ZN => n65679);
   U49153 : AOI22_X1 port map( A1 => n67418, A2 => n66346, B1 => n67412, B2 => 
                           n58340, ZN => n65682);
   U49154 : OAI221_X1 port map( B1 => n54636, B2 => n67430, C1 => n63531, C2 =>
                           n67424, A => n65664, ZN => n65661);
   U49155 : AOI22_X1 port map( A1 => n67418, A2 => n66347, B1 => n67412, B2 => 
                           n58341, ZN => n65664);
   U49156 : OAI221_X1 port map( B1 => n54635, B2 => n67430, C1 => n63530, C2 =>
                           n67424, A => n65646, ZN => n65643);
   U49157 : AOI22_X1 port map( A1 => n67418, A2 => n66348, B1 => n67412, B2 => 
                           n58342, ZN => n65646);
   U49158 : OAI221_X1 port map( B1 => n54634, B2 => n67431, C1 => n63529, C2 =>
                           n67425, A => n65628, ZN => n65625);
   U49159 : AOI22_X1 port map( A1 => n67419, A2 => n66349, B1 => n67413, B2 => 
                           n58343, ZN => n65628);
   U49160 : OAI221_X1 port map( B1 => n54633, B2 => n67431, C1 => n63528, C2 =>
                           n67425, A => n65610, ZN => n65607);
   U49161 : AOI22_X1 port map( A1 => n67419, A2 => n66350, B1 => n67413, B2 => 
                           n58344, ZN => n65610);
   U49162 : OAI221_X1 port map( B1 => n54632, B2 => n67431, C1 => n63527, C2 =>
                           n67425, A => n65592, ZN => n65589);
   U49163 : AOI22_X1 port map( A1 => n67419, A2 => n66351, B1 => n67413, B2 => 
                           n58345, ZN => n65592);
   U49164 : OAI221_X1 port map( B1 => n54631, B2 => n67431, C1 => n63526, C2 =>
                           n67425, A => n65574, ZN => n65571);
   U49165 : AOI22_X1 port map( A1 => n67419, A2 => n66352, B1 => n67413, B2 => 
                           n58346, ZN => n65574);
   U49166 : OAI221_X1 port map( B1 => n54630, B2 => n67431, C1 => n63525, C2 =>
                           n67425, A => n65556, ZN => n65553);
   U49167 : AOI22_X1 port map( A1 => n67419, A2 => n66353, B1 => n67413, B2 => 
                           n58347, ZN => n65556);
   U49168 : OAI221_X1 port map( B1 => n54629, B2 => n67431, C1 => n63524, C2 =>
                           n67425, A => n65538, ZN => n65535);
   U49169 : AOI22_X1 port map( A1 => n67419, A2 => n66354, B1 => n67413, B2 => 
                           n58348, ZN => n65538);
   U49170 : OAI221_X1 port map( B1 => n54628, B2 => n67431, C1 => n63523, C2 =>
                           n67425, A => n65520, ZN => n65517);
   U49171 : AOI22_X1 port map( A1 => n67419, A2 => n66355, B1 => n67413, B2 => 
                           n58349, ZN => n65520);
   U49172 : OAI221_X1 port map( B1 => n54627, B2 => n67431, C1 => n63522, C2 =>
                           n67425, A => n65502, ZN => n65499);
   U49173 : AOI22_X1 port map( A1 => n67419, A2 => n66356, B1 => n67413, B2 => 
                           n58350, ZN => n65502);
   U49174 : OAI221_X1 port map( B1 => n54626, B2 => n67431, C1 => n63521, C2 =>
                           n67425, A => n65484, ZN => n65481);
   U49175 : AOI22_X1 port map( A1 => n67419, A2 => n66357, B1 => n67413, B2 => 
                           n58351, ZN => n65484);
   U49176 : OAI221_X1 port map( B1 => n54625, B2 => n67431, C1 => n63520, C2 =>
                           n67425, A => n65466, ZN => n65463);
   U49177 : AOI22_X1 port map( A1 => n67419, A2 => n66358, B1 => n67413, B2 => 
                           n58352, ZN => n65466);
   U49178 : OAI221_X1 port map( B1 => n54624, B2 => n67431, C1 => n63519, C2 =>
                           n67425, A => n65448, ZN => n65445);
   U49179 : AOI22_X1 port map( A1 => n67419, A2 => n66359, B1 => n67413, B2 => 
                           n58353, ZN => n65448);
   U49180 : OAI221_X1 port map( B1 => n54623, B2 => n67431, C1 => n63518, C2 =>
                           n67425, A => n65430, ZN => n65427);
   U49181 : AOI22_X1 port map( A1 => n67419, A2 => n66360, B1 => n67413, B2 => 
                           n58354, ZN => n65430);
   U49182 : OAI221_X1 port map( B1 => n54622, B2 => n67432, C1 => n63517, C2 =>
                           n67426, A => n65412, ZN => n65409);
   U49183 : AOI22_X1 port map( A1 => n67420, A2 => n66361, B1 => n67414, B2 => 
                           n58355, ZN => n65412);
   U49184 : OAI221_X1 port map( B1 => n54621, B2 => n67432, C1 => n63516, C2 =>
                           n67426, A => n65394, ZN => n65391);
   U49185 : AOI22_X1 port map( A1 => n67420, A2 => n66362, B1 => n67414, B2 => 
                           n58356, ZN => n65394);
   U49186 : OAI221_X1 port map( B1 => n54620, B2 => n67432, C1 => n63515, C2 =>
                           n67426, A => n65376, ZN => n65373);
   U49187 : AOI22_X1 port map( A1 => n67420, A2 => n66363, B1 => n67414, B2 => 
                           n58357, ZN => n65376);
   U49188 : OAI221_X1 port map( B1 => n54619, B2 => n67432, C1 => n63514, C2 =>
                           n67426, A => n65358, ZN => n65355);
   U49189 : AOI22_X1 port map( A1 => n67420, A2 => n66364, B1 => n67414, B2 => 
                           n58358, ZN => n65358);
   U49190 : OAI221_X1 port map( B1 => n54618, B2 => n67432, C1 => n63513, C2 =>
                           n67426, A => n65340, ZN => n65337);
   U49191 : AOI22_X1 port map( A1 => n67420, A2 => n66365, B1 => n67414, B2 => 
                           n58359, ZN => n65340);
   U49192 : OAI221_X1 port map( B1 => n54617, B2 => n67432, C1 => n63512, C2 =>
                           n67426, A => n65322, ZN => n65319);
   U49193 : AOI22_X1 port map( A1 => n67420, A2 => n66366, B1 => n67414, B2 => 
                           n58360, ZN => n65322);
   U49194 : OAI221_X1 port map( B1 => n54616, B2 => n67432, C1 => n63511, C2 =>
                           n67426, A => n65304, ZN => n65301);
   U49195 : AOI22_X1 port map( A1 => n67420, A2 => n66367, B1 => n67414, B2 => 
                           n58361, ZN => n65304);
   U49196 : OAI221_X1 port map( B1 => n54615, B2 => n67432, C1 => n63510, C2 =>
                           n67426, A => n65286, ZN => n65283);
   U49197 : AOI22_X1 port map( A1 => n67420, A2 => n66368, B1 => n67414, B2 => 
                           n58362, ZN => n65286);
   U49198 : OAI221_X1 port map( B1 => n54614, B2 => n67432, C1 => n63509, C2 =>
                           n67426, A => n65268, ZN => n65265);
   U49199 : AOI22_X1 port map( A1 => n67420, A2 => n66369, B1 => n67414, B2 => 
                           n58363, ZN => n65268);
   U49200 : OAI221_X1 port map( B1 => n54613, B2 => n67432, C1 => n63508, C2 =>
                           n67426, A => n65250, ZN => n65247);
   U49201 : AOI22_X1 port map( A1 => n67420, A2 => n66370, B1 => n67414, B2 => 
                           n58364, ZN => n65250);
   U49202 : OAI221_X1 port map( B1 => n54612, B2 => n67432, C1 => n63507, C2 =>
                           n67426, A => n65232, ZN => n65229);
   U49203 : AOI22_X1 port map( A1 => n67420, A2 => n66371, B1 => n67414, B2 => 
                           n58365, ZN => n65232);
   U49204 : OAI221_X1 port map( B1 => n54611, B2 => n67432, C1 => n63506, C2 =>
                           n67426, A => n65214, ZN => n65211);
   U49205 : AOI22_X1 port map( A1 => n67420, A2 => n66372, B1 => n67414, B2 => 
                           n58366, ZN => n65214);
   U49206 : OAI221_X1 port map( B1 => n54608, B2 => n67433, C1 => n63503, C2 =>
                           n67427, A => n65160, ZN => n65157);
   U49207 : AOI22_X1 port map( A1 => n67421, A2 => n66307, B1 => n67415, B2 => 
                           n58306, ZN => n65160);
   U49208 : OAI221_X1 port map( B1 => n54606, B2 => n67433, C1 => n63501, C2 =>
                           n67427, A => n65115, ZN => n65106);
   U49209 : AOI22_X1 port map( A1 => n67421, A2 => n66308, B1 => n67415, B2 => 
                           n58303, ZN => n65115);
   U49210 : OAI221_X1 port map( B1 => n54610, B2 => n67433, C1 => n63505, C2 =>
                           n67427, A => n65196, ZN => n65193);
   U49211 : AOI22_X1 port map( A1 => n67421, A2 => n66305, B1 => n67415, B2 => 
                           n58304, ZN => n65196);
   U49212 : OAI221_X1 port map( B1 => n54609, B2 => n67433, C1 => n63504, C2 =>
                           n67427, A => n65178, ZN => n65175);
   U49213 : AOI22_X1 port map( A1 => n67421, A2 => n66306, B1 => n67415, B2 => 
                           n58305, ZN => n65178);
   U49214 : OAI221_X1 port map( B1 => n62426, B2 => n67409, C1 => n63635, C2 =>
                           n67403, A => n65161, ZN => n65156);
   U49215 : AOI22_X1 port map( A1 => n67397, A2 => n58781, B1 => n67391, B2 => 
                           n58369, ZN => n65161);
   U49216 : OAI221_X1 port map( B1 => n62424, B2 => n67409, C1 => n63633, C2 =>
                           n67403, A => n65120, ZN => n65105);
   U49217 : AOI22_X1 port map( A1 => n67397, A2 => n58782, B1 => n67391, B2 => 
                           n58370, ZN => n65120);
   U49218 : OAI221_X1 port map( B1 => n62428, B2 => n67409, C1 => n63637, C2 =>
                           n67403, A => n65197, ZN => n65192);
   U49219 : AOI22_X1 port map( A1 => n67397, A2 => n58779, B1 => n67391, B2 => 
                           n58367, ZN => n65197);
   U49220 : OAI221_X1 port map( B1 => n62427, B2 => n67409, C1 => n63636, C2 =>
                           n67403, A => n65179, ZN => n65174);
   U49221 : AOI22_X1 port map( A1 => n67397, A2 => n58780, B1 => n67391, B2 => 
                           n58368, ZN => n65179);
   U49222 : OAI221_X1 port map( B1 => n62428, B2 => n67607, C1 => n63505, C2 =>
                           n67601, A => n63873, ZN => n63868);
   U49223 : AOI22_X1 port map( A1 => n67595, A2 => n66499, B1 => n58375, B2 => 
                           n67589, ZN => n63873);
   U49224 : OAI221_X1 port map( B1 => n62427, B2 => n67607, C1 => n63504, C2 =>
                           n67601, A => n63852, ZN => n63847);
   U49225 : AOI22_X1 port map( A1 => n67595, A2 => n66500, B1 => n58376, B2 => 
                           n67589, ZN => n63852);
   U49226 : OAI221_X1 port map( B1 => n62426, B2 => n67607, C1 => n63503, C2 =>
                           n67601, A => n63831, ZN => n63826);
   U49227 : AOI22_X1 port map( A1 => n67595, A2 => n66501, B1 => n58377, B2 => 
                           n67589, ZN => n63831);
   U49228 : OAI221_X1 port map( B1 => n63569, B2 => n67385, C1 => n8481, C2 => 
                           n67379, A => n65162, ZN => n65155);
   U49229 : AOI22_X1 port map( A1 => n67373, A2 => n66497, B1 => n67367, B2 => 
                           n8896, ZN => n65162);
   U49230 : OAI221_X1 port map( B1 => n63567, B2 => n67385, C1 => n8497, C2 => 
                           n67379, A => n65125, ZN => n65104);
   U49231 : AOI22_X1 port map( A1 => n67373, A2 => n66498, B1 => n67367, B2 => 
                           n8895, ZN => n65125);
   U49232 : OAI221_X1 port map( B1 => n63571, B2 => n67385, C1 => n8449, C2 => 
                           n67379, A => n65198, ZN => n65191);
   U49233 : AOI22_X1 port map( A1 => n67373, A2 => n66495, B1 => n67367, B2 => 
                           n8898, ZN => n65198);
   U49234 : OAI221_X1 port map( B1 => n63570, B2 => n67385, C1 => n8465, C2 => 
                           n67379, A => n65180, ZN => n65173);
   U49235 : AOI22_X1 port map( A1 => n67373, A2 => n66496, B1 => n67367, B2 => 
                           n8897, ZN => n65180);
   U49236 : OAI221_X1 port map( B1 => n54186, B2 => n67583, C1 => n63571, C2 =>
                           n67577, A => n63875, ZN => n63867);
   U49237 : AOI22_X1 port map( A1 => n67571, A2 => n8965, B1 => n67565, B2 => 
                           n66495, ZN => n63875);
   U49238 : OAI221_X1 port map( B1 => n54185, B2 => n67583, C1 => n63570, C2 =>
                           n67577, A => n63854, ZN => n63846);
   U49239 : AOI22_X1 port map( A1 => n67571, A2 => n8963, B1 => n67565, B2 => 
                           n66496, ZN => n63854);
   U49240 : OAI221_X1 port map( B1 => n54184, B2 => n67583, C1 => n63569, C2 =>
                           n67577, A => n63833, ZN => n63825);
   U49241 : AOI22_X1 port map( A1 => n67571, A2 => n8961, B1 => n67565, B2 => 
                           n66497, ZN => n63833);
   U49242 : OAI221_X1 port map( B1 => n62694, B2 => n67583, C1 => n63567, C2 =>
                           n67577, A => n63793, ZN => n63771);
   U49243 : AOI22_X1 port map( A1 => n67571, A2 => n8959, B1 => n67565, B2 => 
                           n66498, ZN => n63793);
   U49244 : OAI221_X1 port map( B1 => n54246, B2 => n67578, C1 => n63631, C2 =>
                           n67572, A => n65088, ZN => n65068);
   U49245 : AOI22_X1 port map( A1 => n67566, A2 => n9085, B1 => n67560, B2 => 
                           n58036, ZN => n65088);
   U49246 : OAI221_X1 port map( B1 => n54245, B2 => n67578, C1 => n63630, C2 =>
                           n67572, A => n65056, ZN => n65048);
   U49247 : AOI22_X1 port map( A1 => n67566, A2 => n9083, B1 => n67560, B2 => 
                           n58001, ZN => n65056);
   U49248 : OAI221_X1 port map( B1 => n54244, B2 => n67578, C1 => n63629, C2 =>
                           n67572, A => n65036, ZN => n65028);
   U49249 : AOI22_X1 port map( A1 => n67566, A2 => n9081, B1 => n67560, B2 => 
                           n57977, ZN => n65036);
   U49250 : OAI221_X1 port map( B1 => n54243, B2 => n67578, C1 => n63628, C2 =>
                           n67572, A => n65016, ZN => n65008);
   U49251 : AOI22_X1 port map( A1 => n67566, A2 => n9079, B1 => n67560, B2 => 
                           n57953, ZN => n65016);
   U49252 : OAI221_X1 port map( B1 => n54242, B2 => n67578, C1 => n63627, C2 =>
                           n67572, A => n64996, ZN => n64988);
   U49253 : AOI22_X1 port map( A1 => n67566, A2 => n9077, B1 => n67560, B2 => 
                           n57929, ZN => n64996);
   U49254 : OAI221_X1 port map( B1 => n54241, B2 => n67578, C1 => n63626, C2 =>
                           n67572, A => n64976, ZN => n64968);
   U49255 : AOI22_X1 port map( A1 => n67566, A2 => n9075, B1 => n67560, B2 => 
                           n57905, ZN => n64976);
   U49256 : OAI221_X1 port map( B1 => n54240, B2 => n67578, C1 => n63625, C2 =>
                           n67572, A => n64956, ZN => n64948);
   U49257 : AOI22_X1 port map( A1 => n67566, A2 => n9073, B1 => n67560, B2 => 
                           n57881, ZN => n64956);
   U49258 : OAI221_X1 port map( B1 => n54239, B2 => n67578, C1 => n63624, C2 =>
                           n67572, A => n64936, ZN => n64928);
   U49259 : AOI22_X1 port map( A1 => n67566, A2 => n9071, B1 => n67560, B2 => 
                           n57857, ZN => n64936);
   U49260 : OAI221_X1 port map( B1 => n54238, B2 => n67578, C1 => n63623, C2 =>
                           n67572, A => n64916, ZN => n64908);
   U49261 : AOI22_X1 port map( A1 => n67566, A2 => n9069, B1 => n67560, B2 => 
                           n57833, ZN => n64916);
   U49262 : OAI221_X1 port map( B1 => n54237, B2 => n67578, C1 => n63622, C2 =>
                           n67572, A => n64896, ZN => n64888);
   U49263 : AOI22_X1 port map( A1 => n67566, A2 => n9067, B1 => n67560, B2 => 
                           n57809, ZN => n64896);
   U49264 : OAI221_X1 port map( B1 => n54236, B2 => n67578, C1 => n63621, C2 =>
                           n67572, A => n64876, ZN => n64868);
   U49265 : AOI22_X1 port map( A1 => n67566, A2 => n9065, B1 => n67560, B2 => 
                           n57785, ZN => n64876);
   U49266 : OAI221_X1 port map( B1 => n54235, B2 => n67578, C1 => n63620, C2 =>
                           n67572, A => n64856, ZN => n64848);
   U49267 : AOI22_X1 port map( A1 => n67566, A2 => n9063, B1 => n67560, B2 => 
                           n57761, ZN => n64856);
   U49268 : OAI22_X1 port map( A1 => n54184, A2 => n67361, B1 => n49482, B2 => 
                           n67355, ZN => n65166);
   U49269 : OAI22_X1 port map( A1 => n62694, A2 => n67361, B1 => n49483, B2 => 
                           n67355, ZN => n65131);
   U49270 : OAI22_X1 port map( A1 => n54186, A2 => n67361, B1 => n49480, B2 => 
                           n67355, ZN => n65202);
   U49271 : OAI22_X1 port map( A1 => n54185, A2 => n67361, B1 => n49481, B2 => 
                           n67355, ZN => n65184);
   U49272 : OAI22_X1 port map( A1 => n62691, A2 => n67554, B1 => n54670, B2 => 
                           n67548, ZN => n65092);
   U49273 : OAI22_X1 port map( A1 => n62690, A2 => n67554, B1 => n54669, B2 => 
                           n67548, ZN => n65060);
   U49274 : OAI22_X1 port map( A1 => n62689, A2 => n67554, B1 => n54668, B2 => 
                           n67548, ZN => n65040);
   U49275 : OAI22_X1 port map( A1 => n62688, A2 => n67554, B1 => n54667, B2 => 
                           n67548, ZN => n65020);
   U49276 : OAI22_X1 port map( A1 => n62687, A2 => n67554, B1 => n54666, B2 => 
                           n67548, ZN => n65000);
   U49277 : OAI22_X1 port map( A1 => n62686, A2 => n67554, B1 => n54665, B2 => 
                           n67548, ZN => n64980);
   U49278 : OAI22_X1 port map( A1 => n62685, A2 => n67554, B1 => n54664, B2 => 
                           n67548, ZN => n64960);
   U49279 : OAI22_X1 port map( A1 => n62684, A2 => n67554, B1 => n54663, B2 => 
                           n67548, ZN => n64940);
   U49280 : OAI22_X1 port map( A1 => n62683, A2 => n67554, B1 => n54662, B2 => 
                           n67548, ZN => n64920);
   U49281 : OAI22_X1 port map( A1 => n62682, A2 => n67554, B1 => n54661, B2 => 
                           n67548, ZN => n64900);
   U49282 : OAI22_X1 port map( A1 => n62681, A2 => n67554, B1 => n54660, B2 => 
                           n67548, ZN => n64880);
   U49283 : OAI22_X1 port map( A1 => n62680, A2 => n67554, B1 => n54659, B2 => 
                           n67548, ZN => n64860);
   U49284 : OAI22_X1 port map( A1 => n62679, A2 => n67555, B1 => n54658, B2 => 
                           n67549, ZN => n64840);
   U49285 : OAI22_X1 port map( A1 => n62678, A2 => n67555, B1 => n54657, B2 => 
                           n67549, ZN => n64820);
   U49286 : OAI22_X1 port map( A1 => n62677, A2 => n67555, B1 => n54656, B2 => 
                           n67549, ZN => n64800);
   U49287 : OAI22_X1 port map( A1 => n62676, A2 => n67555, B1 => n54655, B2 => 
                           n67549, ZN => n64780);
   U49288 : OAI22_X1 port map( A1 => n62675, A2 => n67555, B1 => n54654, B2 => 
                           n67549, ZN => n64760);
   U49289 : OAI22_X1 port map( A1 => n62674, A2 => n67555, B1 => n54653, B2 => 
                           n67549, ZN => n64740);
   U49290 : OAI22_X1 port map( A1 => n62673, A2 => n67555, B1 => n54652, B2 => 
                           n67549, ZN => n64720);
   U49291 : OAI22_X1 port map( A1 => n62672, A2 => n67555, B1 => n54651, B2 => 
                           n67549, ZN => n64700);
   U49292 : OAI22_X1 port map( A1 => n62671, A2 => n67555, B1 => n54650, B2 => 
                           n67549, ZN => n64680);
   U49293 : OAI22_X1 port map( A1 => n62670, A2 => n67555, B1 => n54649, B2 => 
                           n67549, ZN => n64660);
   U49294 : OAI22_X1 port map( A1 => n62669, A2 => n67555, B1 => n54648, B2 => 
                           n67549, ZN => n64640);
   U49295 : OAI22_X1 port map( A1 => n62668, A2 => n67555, B1 => n54647, B2 => 
                           n67549, ZN => n64620);
   U49296 : OAI22_X1 port map( A1 => n62667, A2 => n67556, B1 => n54646, B2 => 
                           n67550, ZN => n64600);
   U49297 : OAI22_X1 port map( A1 => n62666, A2 => n67556, B1 => n54645, B2 => 
                           n67550, ZN => n64580);
   U49298 : OAI22_X1 port map( A1 => n62665, A2 => n67556, B1 => n54644, B2 => 
                           n67550, ZN => n64560);
   U49299 : OAI22_X1 port map( A1 => n62664, A2 => n67556, B1 => n54643, B2 => 
                           n67550, ZN => n64540);
   U49300 : OAI22_X1 port map( A1 => n62663, A2 => n67556, B1 => n54642, B2 => 
                           n67550, ZN => n64520);
   U49301 : OAI22_X1 port map( A1 => n62662, A2 => n67556, B1 => n54641, B2 => 
                           n67550, ZN => n64500);
   U49302 : OAI22_X1 port map( A1 => n62661, A2 => n67556, B1 => n54640, B2 => 
                           n67550, ZN => n64480);
   U49303 : OAI22_X1 port map( A1 => n62660, A2 => n67556, B1 => n54639, B2 => 
                           n67550, ZN => n64460);
   U49304 : OAI22_X1 port map( A1 => n62659, A2 => n67556, B1 => n54638, B2 => 
                           n67550, ZN => n64440);
   U49305 : OAI22_X1 port map( A1 => n62658, A2 => n67556, B1 => n54637, B2 => 
                           n67550, ZN => n64420);
   U49306 : OAI22_X1 port map( A1 => n62657, A2 => n67556, B1 => n54636, B2 => 
                           n67550, ZN => n64400);
   U49307 : OAI22_X1 port map( A1 => n62656, A2 => n67556, B1 => n54635, B2 => 
                           n67550, ZN => n64380);
   U49308 : OAI22_X1 port map( A1 => n62655, A2 => n67557, B1 => n54634, B2 => 
                           n67551, ZN => n64360);
   U49309 : OAI22_X1 port map( A1 => n62654, A2 => n67557, B1 => n54633, B2 => 
                           n67551, ZN => n64340);
   U49310 : OAI22_X1 port map( A1 => n62653, A2 => n67557, B1 => n54632, B2 => 
                           n67551, ZN => n64320);
   U49311 : OAI22_X1 port map( A1 => n62652, A2 => n67557, B1 => n54631, B2 => 
                           n67551, ZN => n64300);
   U49312 : OAI22_X1 port map( A1 => n62651, A2 => n67557, B1 => n54630, B2 => 
                           n67551, ZN => n64280);
   U49313 : OAI22_X1 port map( A1 => n62650, A2 => n67557, B1 => n54629, B2 => 
                           n67551, ZN => n64260);
   U49314 : OAI22_X1 port map( A1 => n62649, A2 => n67557, B1 => n54628, B2 => 
                           n67551, ZN => n64240);
   U49315 : OAI22_X1 port map( A1 => n62648, A2 => n67557, B1 => n54627, B2 => 
                           n67551, ZN => n64220);
   U49316 : OAI22_X1 port map( A1 => n62647, A2 => n67557, B1 => n54626, B2 => 
                           n67551, ZN => n64200);
   U49317 : OAI22_X1 port map( A1 => n62646, A2 => n67557, B1 => n54625, B2 => 
                           n67551, ZN => n64180);
   U49318 : OAI22_X1 port map( A1 => n62645, A2 => n67557, B1 => n54624, B2 => 
                           n67551, ZN => n64160);
   U49319 : OAI22_X1 port map( A1 => n62644, A2 => n67557, B1 => n54623, B2 => 
                           n67551, ZN => n64140);
   U49320 : OAI22_X1 port map( A1 => n62643, A2 => n67558, B1 => n54622, B2 => 
                           n67552, ZN => n64120);
   U49321 : OAI22_X1 port map( A1 => n62642, A2 => n67558, B1 => n54621, B2 => 
                           n67552, ZN => n64100);
   U49322 : OAI22_X1 port map( A1 => n62641, A2 => n67558, B1 => n54620, B2 => 
                           n67552, ZN => n64080);
   U49323 : OAI22_X1 port map( A1 => n62640, A2 => n67558, B1 => n54619, B2 => 
                           n67552, ZN => n64060);
   U49324 : OAI22_X1 port map( A1 => n62639, A2 => n67558, B1 => n54618, B2 => 
                           n67552, ZN => n64040);
   U49325 : OAI22_X1 port map( A1 => n62638, A2 => n67558, B1 => n54617, B2 => 
                           n67552, ZN => n64020);
   U49326 : OAI22_X1 port map( A1 => n62637, A2 => n67558, B1 => n54616, B2 => 
                           n67552, ZN => n64000);
   U49327 : OAI22_X1 port map( A1 => n62636, A2 => n67558, B1 => n54615, B2 => 
                           n67552, ZN => n63980);
   U49328 : OAI22_X1 port map( A1 => n62635, A2 => n67558, B1 => n54614, B2 => 
                           n67552, ZN => n63960);
   U49329 : OAI22_X1 port map( A1 => n62634, A2 => n67558, B1 => n54613, B2 => 
                           n67552, ZN => n63940);
   U49330 : OAI22_X1 port map( A1 => n62633, A2 => n67558, B1 => n54612, B2 => 
                           n67552, ZN => n63920);
   U49331 : OAI22_X1 port map( A1 => n62632, A2 => n67558, B1 => n54611, B2 => 
                           n67552, ZN => n63900);
   U49332 : OAI22_X1 port map( A1 => n54246, A2 => n67356, B1 => n49420, B2 => 
                           n67350, ZN => n66296);
   U49333 : OAI22_X1 port map( A1 => n54245, A2 => n67356, B1 => n49421, B2 => 
                           n67350, ZN => n66264);
   U49334 : OAI22_X1 port map( A1 => n54244, A2 => n67356, B1 => n49422, B2 => 
                           n67350, ZN => n66246);
   U49335 : OAI22_X1 port map( A1 => n54243, A2 => n67356, B1 => n49423, B2 => 
                           n67350, ZN => n66228);
   U49336 : OAI22_X1 port map( A1 => n54242, A2 => n67356, B1 => n49424, B2 => 
                           n67350, ZN => n66210);
   U49337 : OAI22_X1 port map( A1 => n54241, A2 => n67356, B1 => n49425, B2 => 
                           n67350, ZN => n66192);
   U49338 : OAI22_X1 port map( A1 => n54240, A2 => n67356, B1 => n49426, B2 => 
                           n67350, ZN => n66174);
   U49339 : OAI22_X1 port map( A1 => n54239, A2 => n67356, B1 => n49427, B2 => 
                           n67350, ZN => n66156);
   U49340 : OAI22_X1 port map( A1 => n54238, A2 => n67356, B1 => n49428, B2 => 
                           n67350, ZN => n66138);
   U49341 : OAI22_X1 port map( A1 => n54237, A2 => n67356, B1 => n49429, B2 => 
                           n67350, ZN => n66120);
   U49342 : OAI22_X1 port map( A1 => n54236, A2 => n67356, B1 => n49430, B2 => 
                           n67350, ZN => n66102);
   U49343 : OAI22_X1 port map( A1 => n54235, A2 => n67356, B1 => n49431, B2 => 
                           n67350, ZN => n66084);
   U49344 : OAI22_X1 port map( A1 => n54234, A2 => n67357, B1 => n49432, B2 => 
                           n67351, ZN => n66066);
   U49345 : OAI22_X1 port map( A1 => n54233, A2 => n67357, B1 => n49433, B2 => 
                           n67351, ZN => n66048);
   U49346 : OAI22_X1 port map( A1 => n54232, A2 => n67357, B1 => n49434, B2 => 
                           n67351, ZN => n66030);
   U49347 : OAI22_X1 port map( A1 => n54231, A2 => n67357, B1 => n49435, B2 => 
                           n67351, ZN => n66012);
   U49348 : OAI22_X1 port map( A1 => n54230, A2 => n67357, B1 => n49436, B2 => 
                           n67351, ZN => n65994);
   U49349 : OAI22_X1 port map( A1 => n54229, A2 => n67357, B1 => n49437, B2 => 
                           n67351, ZN => n65976);
   U49350 : OAI22_X1 port map( A1 => n54228, A2 => n67357, B1 => n49438, B2 => 
                           n67351, ZN => n65958);
   U49351 : OAI22_X1 port map( A1 => n54227, A2 => n67357, B1 => n49439, B2 => 
                           n67351, ZN => n65940);
   U49352 : OAI22_X1 port map( A1 => n54226, A2 => n67357, B1 => n49440, B2 => 
                           n67351, ZN => n65922);
   U49353 : OAI22_X1 port map( A1 => n54225, A2 => n67357, B1 => n49441, B2 => 
                           n67351, ZN => n65904);
   U49354 : OAI22_X1 port map( A1 => n54224, A2 => n67357, B1 => n49442, B2 => 
                           n67351, ZN => n65886);
   U49355 : OAI22_X1 port map( A1 => n54223, A2 => n67357, B1 => n49443, B2 => 
                           n67351, ZN => n65868);
   U49356 : OAI22_X1 port map( A1 => n54222, A2 => n67358, B1 => n49444, B2 => 
                           n67352, ZN => n65850);
   U49357 : OAI22_X1 port map( A1 => n54221, A2 => n67358, B1 => n49445, B2 => 
                           n67352, ZN => n65832);
   U49358 : OAI22_X1 port map( A1 => n54220, A2 => n67358, B1 => n49446, B2 => 
                           n67352, ZN => n65814);
   U49359 : OAI22_X1 port map( A1 => n54219, A2 => n67358, B1 => n49447, B2 => 
                           n67352, ZN => n65796);
   U49360 : OAI22_X1 port map( A1 => n54218, A2 => n67358, B1 => n49448, B2 => 
                           n67352, ZN => n65778);
   U49361 : OAI22_X1 port map( A1 => n54217, A2 => n67358, B1 => n49449, B2 => 
                           n67352, ZN => n65760);
   U49362 : OAI22_X1 port map( A1 => n54216, A2 => n67358, B1 => n49450, B2 => 
                           n67352, ZN => n65742);
   U49363 : OAI22_X1 port map( A1 => n54215, A2 => n67358, B1 => n49451, B2 => 
                           n67352, ZN => n65724);
   U49364 : OAI22_X1 port map( A1 => n54214, A2 => n67358, B1 => n49452, B2 => 
                           n67352, ZN => n65706);
   U49365 : OAI22_X1 port map( A1 => n54213, A2 => n67358, B1 => n49453, B2 => 
                           n67352, ZN => n65688);
   U49366 : OAI22_X1 port map( A1 => n54212, A2 => n67358, B1 => n49454, B2 => 
                           n67352, ZN => n65670);
   U49367 : OAI22_X1 port map( A1 => n54211, A2 => n67358, B1 => n49455, B2 => 
                           n67352, ZN => n65652);
   U49368 : OAI22_X1 port map( A1 => n54210, A2 => n67359, B1 => n49456, B2 => 
                           n67353, ZN => n65634);
   U49369 : OAI22_X1 port map( A1 => n54209, A2 => n67359, B1 => n49457, B2 => 
                           n67353, ZN => n65616);
   U49370 : OAI22_X1 port map( A1 => n54208, A2 => n67359, B1 => n49458, B2 => 
                           n67353, ZN => n65598);
   U49371 : OAI22_X1 port map( A1 => n54207, A2 => n67359, B1 => n49459, B2 => 
                           n67353, ZN => n65580);
   U49372 : OAI22_X1 port map( A1 => n54206, A2 => n67359, B1 => n49460, B2 => 
                           n67353, ZN => n65562);
   U49373 : OAI22_X1 port map( A1 => n54205, A2 => n67359, B1 => n49461, B2 => 
                           n67353, ZN => n65544);
   U49374 : OAI22_X1 port map( A1 => n54204, A2 => n67359, B1 => n49462, B2 => 
                           n67353, ZN => n65526);
   U49375 : OAI22_X1 port map( A1 => n54203, A2 => n67359, B1 => n49463, B2 => 
                           n67353, ZN => n65508);
   U49376 : OAI22_X1 port map( A1 => n54202, A2 => n67359, B1 => n49464, B2 => 
                           n67353, ZN => n65490);
   U49377 : OAI22_X1 port map( A1 => n54201, A2 => n67359, B1 => n49465, B2 => 
                           n67353, ZN => n65472);
   U49378 : OAI22_X1 port map( A1 => n54200, A2 => n67359, B1 => n49466, B2 => 
                           n67353, ZN => n65454);
   U49379 : OAI22_X1 port map( A1 => n54199, A2 => n67359, B1 => n49467, B2 => 
                           n67353, ZN => n65436);
   U49380 : OAI22_X1 port map( A1 => n54198, A2 => n67360, B1 => n49468, B2 => 
                           n67354, ZN => n65418);
   U49381 : OAI22_X1 port map( A1 => n54197, A2 => n67360, B1 => n49469, B2 => 
                           n67354, ZN => n65400);
   U49382 : OAI22_X1 port map( A1 => n54196, A2 => n67360, B1 => n49470, B2 => 
                           n67354, ZN => n65382);
   U49383 : OAI22_X1 port map( A1 => n54195, A2 => n67360, B1 => n49471, B2 => 
                           n67354, ZN => n65364);
   U49384 : OAI22_X1 port map( A1 => n54194, A2 => n67360, B1 => n49472, B2 => 
                           n67354, ZN => n65346);
   U49385 : OAI22_X1 port map( A1 => n54193, A2 => n67360, B1 => n49473, B2 => 
                           n67354, ZN => n65328);
   U49386 : OAI22_X1 port map( A1 => n54192, A2 => n67360, B1 => n49474, B2 => 
                           n67354, ZN => n65310);
   U49387 : OAI22_X1 port map( A1 => n54191, A2 => n67360, B1 => n49475, B2 => 
                           n67354, ZN => n65292);
   U49388 : OAI22_X1 port map( A1 => n54190, A2 => n67360, B1 => n49476, B2 => 
                           n67354, ZN => n65274);
   U49389 : OAI22_X1 port map( A1 => n54189, A2 => n67360, B1 => n49477, B2 => 
                           n67354, ZN => n65256);
   U49390 : OAI22_X1 port map( A1 => n54188, A2 => n67360, B1 => n49478, B2 => 
                           n67354, ZN => n65238);
   U49391 : OAI22_X1 port map( A1 => n54187, A2 => n67360, B1 => n49479, B2 => 
                           n67354, ZN => n65220);
   U49392 : OAI22_X1 port map( A1 => n7489, A2 => n67542, B1 => n62422, B2 => 
                           n67536, ZN => n65091);
   U49393 : OAI22_X1 port map( A1 => n7505, A2 => n67542, B1 => n62421, B2 => 
                           n67536, ZN => n65059);
   U49394 : OAI22_X1 port map( A1 => n7521, A2 => n67542, B1 => n62420, B2 => 
                           n67536, ZN => n65039);
   U49395 : OAI22_X1 port map( A1 => n7537, A2 => n67542, B1 => n62419, B2 => 
                           n67536, ZN => n65019);
   U49396 : OAI22_X1 port map( A1 => n7553, A2 => n67542, B1 => n62418, B2 => 
                           n67536, ZN => n64999);
   U49397 : OAI22_X1 port map( A1 => n7569, A2 => n67542, B1 => n62417, B2 => 
                           n67536, ZN => n64979);
   U49398 : OAI22_X1 port map( A1 => n7585, A2 => n67542, B1 => n62416, B2 => 
                           n67536, ZN => n64959);
   U49399 : OAI22_X1 port map( A1 => n7601, A2 => n67542, B1 => n62415, B2 => 
                           n67536, ZN => n64939);
   U49400 : OAI22_X1 port map( A1 => n7617, A2 => n67542, B1 => n62414, B2 => 
                           n67536, ZN => n64919);
   U49401 : OAI22_X1 port map( A1 => n7633, A2 => n67542, B1 => n62413, B2 => 
                           n67536, ZN => n64899);
   U49402 : OAI22_X1 port map( A1 => n7649, A2 => n67542, B1 => n62412, B2 => 
                           n67536, ZN => n64879);
   U49403 : OAI22_X1 port map( A1 => n7665, A2 => n67542, B1 => n62411, B2 => 
                           n67536, ZN => n64859);
   U49404 : OAI22_X1 port map( A1 => n7681, A2 => n67543, B1 => n62410, B2 => 
                           n67537, ZN => n64839);
   U49405 : OAI22_X1 port map( A1 => n7697, A2 => n67543, B1 => n62409, B2 => 
                           n67537, ZN => n64819);
   U49406 : OAI22_X1 port map( A1 => n7713, A2 => n67543, B1 => n62408, B2 => 
                           n67537, ZN => n64799);
   U49407 : OAI22_X1 port map( A1 => n7729, A2 => n67543, B1 => n62407, B2 => 
                           n67537, ZN => n64779);
   U49408 : OAI22_X1 port map( A1 => n7745, A2 => n67543, B1 => n62406, B2 => 
                           n67537, ZN => n64759);
   U49409 : OAI22_X1 port map( A1 => n7761, A2 => n67543, B1 => n62405, B2 => 
                           n67537, ZN => n64739);
   U49410 : OAI22_X1 port map( A1 => n7777, A2 => n67543, B1 => n62404, B2 => 
                           n67537, ZN => n64719);
   U49411 : OAI22_X1 port map( A1 => n7793, A2 => n67543, B1 => n62403, B2 => 
                           n67537, ZN => n64699);
   U49412 : OAI22_X1 port map( A1 => n7809, A2 => n67543, B1 => n62402, B2 => 
                           n67537, ZN => n64679);
   U49413 : OAI22_X1 port map( A1 => n7825, A2 => n67543, B1 => n62401, B2 => 
                           n67537, ZN => n64659);
   U49414 : OAI22_X1 port map( A1 => n7841, A2 => n67543, B1 => n62400, B2 => 
                           n67537, ZN => n64639);
   U49415 : OAI22_X1 port map( A1 => n7857, A2 => n67543, B1 => n62399, B2 => 
                           n67537, ZN => n64619);
   U49416 : OAI22_X1 port map( A1 => n7873, A2 => n67544, B1 => n62398, B2 => 
                           n67538, ZN => n64599);
   U49417 : OAI22_X1 port map( A1 => n7889, A2 => n67544, B1 => n62397, B2 => 
                           n67538, ZN => n64579);
   U49418 : OAI22_X1 port map( A1 => n7905, A2 => n67544, B1 => n62396, B2 => 
                           n67538, ZN => n64559);
   U49419 : OAI22_X1 port map( A1 => n7921, A2 => n67544, B1 => n62395, B2 => 
                           n67538, ZN => n64539);
   U49420 : OAI22_X1 port map( A1 => n7937, A2 => n67544, B1 => n62394, B2 => 
                           n67538, ZN => n64519);
   U49421 : OAI22_X1 port map( A1 => n7953, A2 => n67544, B1 => n62393, B2 => 
                           n67538, ZN => n64499);
   U49422 : OAI22_X1 port map( A1 => n7969, A2 => n67544, B1 => n62392, B2 => 
                           n67538, ZN => n64479);
   U49423 : OAI22_X1 port map( A1 => n7985, A2 => n67544, B1 => n62391, B2 => 
                           n67538, ZN => n64459);
   U49424 : OAI22_X1 port map( A1 => n8001, A2 => n67544, B1 => n62390, B2 => 
                           n67538, ZN => n64439);
   U49425 : OAI22_X1 port map( A1 => n8017, A2 => n67544, B1 => n62389, B2 => 
                           n67538, ZN => n64419);
   U49426 : OAI22_X1 port map( A1 => n8033, A2 => n67544, B1 => n62388, B2 => 
                           n67538, ZN => n64399);
   U49427 : OAI22_X1 port map( A1 => n8049, A2 => n67544, B1 => n62387, B2 => 
                           n67538, ZN => n64379);
   U49428 : OAI22_X1 port map( A1 => n8065, A2 => n67545, B1 => n62386, B2 => 
                           n67539, ZN => n64359);
   U49429 : OAI22_X1 port map( A1 => n8081, A2 => n67545, B1 => n62385, B2 => 
                           n67539, ZN => n64339);
   U49430 : OAI22_X1 port map( A1 => n8097, A2 => n67545, B1 => n62384, B2 => 
                           n67539, ZN => n64319);
   U49431 : OAI22_X1 port map( A1 => n8113, A2 => n67545, B1 => n62383, B2 => 
                           n67539, ZN => n64299);
   U49432 : OAI22_X1 port map( A1 => n8129, A2 => n67545, B1 => n62382, B2 => 
                           n67539, ZN => n64279);
   U49433 : OAI22_X1 port map( A1 => n8145, A2 => n67545, B1 => n62381, B2 => 
                           n67539, ZN => n64259);
   U49434 : OAI22_X1 port map( A1 => n8161, A2 => n67545, B1 => n62380, B2 => 
                           n67539, ZN => n64239);
   U49435 : OAI22_X1 port map( A1 => n8177, A2 => n67545, B1 => n62379, B2 => 
                           n67539, ZN => n64219);
   U49436 : OAI22_X1 port map( A1 => n8193, A2 => n67545, B1 => n62378, B2 => 
                           n67539, ZN => n64199);
   U49437 : OAI22_X1 port map( A1 => n8209, A2 => n67545, B1 => n62377, B2 => 
                           n67539, ZN => n64179);
   U49438 : OAI22_X1 port map( A1 => n8225, A2 => n67545, B1 => n62376, B2 => 
                           n67539, ZN => n64159);
   U49439 : OAI22_X1 port map( A1 => n8241, A2 => n67545, B1 => n62375, B2 => 
                           n67539, ZN => n64139);
   U49440 : OAI22_X1 port map( A1 => n8257, A2 => n67546, B1 => n62374, B2 => 
                           n67540, ZN => n64119);
   U49441 : OAI22_X1 port map( A1 => n8273, A2 => n67546, B1 => n62373, B2 => 
                           n67540, ZN => n64099);
   U49442 : OAI22_X1 port map( A1 => n8289, A2 => n67546, B1 => n62372, B2 => 
                           n67540, ZN => n64079);
   U49443 : OAI22_X1 port map( A1 => n8305, A2 => n67546, B1 => n62371, B2 => 
                           n67540, ZN => n64059);
   U49444 : OAI22_X1 port map( A1 => n8321, A2 => n67546, B1 => n62370, B2 => 
                           n67540, ZN => n64039);
   U49445 : OAI22_X1 port map( A1 => n8337, A2 => n67546, B1 => n62369, B2 => 
                           n67540, ZN => n64019);
   U49446 : OAI22_X1 port map( A1 => n8353, A2 => n67546, B1 => n62368, B2 => 
                           n67540, ZN => n63999);
   U49447 : OAI22_X1 port map( A1 => n8369, A2 => n67546, B1 => n62367, B2 => 
                           n67540, ZN => n63979);
   U49448 : OAI22_X1 port map( A1 => n8385, A2 => n67546, B1 => n62366, B2 => 
                           n67540, ZN => n63959);
   U49449 : OAI22_X1 port map( A1 => n8401, A2 => n67546, B1 => n62365, B2 => 
                           n67540, ZN => n63939);
   U49450 : OAI22_X1 port map( A1 => n8417, A2 => n67546, B1 => n62364, B2 => 
                           n67540, ZN => n63919);
   U49451 : OAI22_X1 port map( A1 => n8433, A2 => n67546, B1 => n62363, B2 => 
                           n67540, ZN => n63899);
   U49452 : AND3_X1 port map( A1 => ADD_RD1(2), A2 => n66494, A3 => ADD_RD1(1),
                           ZN => n65074);
   U49453 : OAI22_X1 port map( A1 => n68259, A2 => n62061, B1 => n68251, B2 => 
                           n68094, ZN => n7435);
   U49454 : OAI22_X1 port map( A1 => n68259, A2 => n62059, B1 => n68251, B2 => 
                           n68097, ZN => n7436);
   U49455 : OAI22_X1 port map( A1 => n68259, A2 => n62057, B1 => n68251, B2 => 
                           n68100, ZN => n7437);
   U49456 : OAI22_X1 port map( A1 => n68259, A2 => n62055, B1 => n68251, B2 => 
                           n68103, ZN => n7438);
   U49457 : OAI22_X1 port map( A1 => n68259, A2 => n62053, B1 => n68251, B2 => 
                           n68106, ZN => n7439);
   U49458 : OAI22_X1 port map( A1 => n68259, A2 => n62051, B1 => n68251, B2 => 
                           n68109, ZN => n7440);
   U49459 : OAI22_X1 port map( A1 => n68259, A2 => n62049, B1 => n68251, B2 => 
                           n68112, ZN => n7441);
   U49460 : OAI22_X1 port map( A1 => n68259, A2 => n62047, B1 => n68251, B2 => 
                           n68115, ZN => n7442);
   U49461 : OAI22_X1 port map( A1 => n68259, A2 => n62045, B1 => n68251, B2 => 
                           n68118, ZN => n7443);
   U49462 : OAI22_X1 port map( A1 => n68259, A2 => n62043, B1 => n68251, B2 => 
                           n68121, ZN => n7444);
   U49463 : OAI22_X1 port map( A1 => n68259, A2 => n62041, B1 => n68251, B2 => 
                           n68124, ZN => n7445);
   U49464 : OAI22_X1 port map( A1 => n68259, A2 => n62039, B1 => n68251, B2 => 
                           n68127, ZN => n7446);
   U49465 : OAI22_X1 port map( A1 => n68259, A2 => n62037, B1 => n68252, B2 => 
                           n68130, ZN => n7447);
   U49466 : OAI22_X1 port map( A1 => n68260, A2 => n62035, B1 => n68252, B2 => 
                           n68133, ZN => n7448);
   U49467 : OAI22_X1 port map( A1 => n68260, A2 => n62033, B1 => n68252, B2 => 
                           n68136, ZN => n7449);
   U49468 : OAI22_X1 port map( A1 => n68260, A2 => n62031, B1 => n68252, B2 => 
                           n68139, ZN => n7450);
   U49469 : OAI22_X1 port map( A1 => n68260, A2 => n62029, B1 => n68252, B2 => 
                           n68142, ZN => n7451);
   U49470 : OAI22_X1 port map( A1 => n68260, A2 => n62027, B1 => n68252, B2 => 
                           n68145, ZN => n7452);
   U49471 : OAI22_X1 port map( A1 => n68260, A2 => n62025, B1 => n68252, B2 => 
                           n68148, ZN => n7453);
   U49472 : OAI22_X1 port map( A1 => n68260, A2 => n62023, B1 => n68252, B2 => 
                           n68151, ZN => n7454);
   U49473 : OAI22_X1 port map( A1 => n68260, A2 => n62021, B1 => n68252, B2 => 
                           n68154, ZN => n7455);
   U49474 : OAI22_X1 port map( A1 => n68260, A2 => n62019, B1 => n68252, B2 => 
                           n68157, ZN => n7456);
   U49475 : OAI22_X1 port map( A1 => n68260, A2 => n62017, B1 => n68252, B2 => 
                           n68160, ZN => n7457);
   U49476 : OAI22_X1 port map( A1 => n68260, A2 => n62015, B1 => n68252, B2 => 
                           n68163, ZN => n7458);
   U49477 : OAI22_X1 port map( A1 => n68260, A2 => n62013, B1 => n68253, B2 => 
                           n68166, ZN => n7459);
   U49478 : OAI22_X1 port map( A1 => n68260, A2 => n62011, B1 => n68253, B2 => 
                           n68169, ZN => n7460);
   U49479 : OAI22_X1 port map( A1 => n68261, A2 => n62009, B1 => n68253, B2 => 
                           n68172, ZN => n7461);
   U49480 : OAI22_X1 port map( A1 => n68261, A2 => n62007, B1 => n68253, B2 => 
                           n68175, ZN => n7462);
   U49481 : OAI22_X1 port map( A1 => n68261, A2 => n62005, B1 => n68253, B2 => 
                           n68178, ZN => n7463);
   U49482 : OAI22_X1 port map( A1 => n68261, A2 => n62003, B1 => n68253, B2 => 
                           n68181, ZN => n7464);
   U49483 : OAI22_X1 port map( A1 => n68261, A2 => n62001, B1 => n68253, B2 => 
                           n68184, ZN => n7465);
   U49484 : OAI22_X1 port map( A1 => n68261, A2 => n61999, B1 => n68253, B2 => 
                           n68187, ZN => n7466);
   U49485 : OAI22_X1 port map( A1 => n68261, A2 => n61997, B1 => n68253, B2 => 
                           n68190, ZN => n7467);
   U49486 : OAI22_X1 port map( A1 => n68261, A2 => n61995, B1 => n68253, B2 => 
                           n68193, ZN => n7468);
   U49487 : OAI22_X1 port map( A1 => n68261, A2 => n61993, B1 => n68253, B2 => 
                           n68196, ZN => n7469);
   U49488 : OAI22_X1 port map( A1 => n68261, A2 => n61991, B1 => n68253, B2 => 
                           n68199, ZN => n7470);
   U49489 : OAI22_X1 port map( A1 => n68261, A2 => n61989, B1 => n68254, B2 => 
                           n68202, ZN => n7471);
   U49490 : OAI22_X1 port map( A1 => n68261, A2 => n61987, B1 => n68254, B2 => 
                           n68205, ZN => n7472);
   U49491 : OAI22_X1 port map( A1 => n68261, A2 => n61985, B1 => n68254, B2 => 
                           n68208, ZN => n7473);
   U49492 : OAI22_X1 port map( A1 => n68262, A2 => n61983, B1 => n68254, B2 => 
                           n68211, ZN => n7474);
   U49493 : OAI22_X1 port map( A1 => n68262, A2 => n61981, B1 => n68254, B2 => 
                           n68214, ZN => n7475);
   U49494 : OAI22_X1 port map( A1 => n68262, A2 => n61979, B1 => n68254, B2 => 
                           n68217, ZN => n7476);
   U49495 : OAI22_X1 port map( A1 => n68262, A2 => n61977, B1 => n68254, B2 => 
                           n68220, ZN => n7477);
   U49496 : OAI22_X1 port map( A1 => n68262, A2 => n61975, B1 => n68254, B2 => 
                           n68223, ZN => n7478);
   U49497 : OAI22_X1 port map( A1 => n68262, A2 => n61973, B1 => n68254, B2 => 
                           n68226, ZN => n7479);
   U49498 : OAI22_X1 port map( A1 => n68262, A2 => n61971, B1 => n68254, B2 => 
                           n68229, ZN => n7480);
   U49499 : OAI22_X1 port map( A1 => n68262, A2 => n61969, B1 => n68254, B2 => 
                           n68232, ZN => n7481);
   U49500 : OAI22_X1 port map( A1 => n68262, A2 => n61967, B1 => n68254, B2 => 
                           n68235, ZN => n7482);
   U49501 : OAI22_X1 port map( A1 => n68262, A2 => n61965, B1 => n68255, B2 => 
                           n68238, ZN => n7483);
   U49502 : OAI22_X1 port map( A1 => n68262, A2 => n61963, B1 => n68255, B2 => 
                           n68241, ZN => n7484);
   U49503 : OAI22_X1 port map( A1 => n68262, A2 => n61961, B1 => n68255, B2 => 
                           n68244, ZN => n7485);
   U49504 : OAI22_X1 port map( A1 => n68262, A2 => n61958, B1 => n68255, B2 => 
                           n68247, ZN => n7486);
   U49505 : AOI22_X1 port map( A1 => n67594, A2 => n66502, B1 => n58427, B2 => 
                           n67588, ZN => n64114);
   U49506 : AOI22_X1 port map( A1 => n67594, A2 => n66503, B1 => n58428, B2 => 
                           n67588, ZN => n64094);
   U49507 : AOI22_X1 port map( A1 => n67594, A2 => n66504, B1 => n58429, B2 => 
                           n67588, ZN => n64074);
   U49508 : AOI22_X1 port map( A1 => n67594, A2 => n66505, B1 => n58430, B2 => 
                           n67588, ZN => n64054);
   U49509 : AOI22_X1 port map( A1 => n67594, A2 => n66506, B1 => n58431, B2 => 
                           n67588, ZN => n64034);
   U49510 : AOI22_X1 port map( A1 => n67594, A2 => n66507, B1 => n58432, B2 => 
                           n67588, ZN => n64014);
   U49511 : AOI22_X1 port map( A1 => n67594, A2 => n66508, B1 => n58433, B2 => 
                           n67588, ZN => n63994);
   U49512 : AOI22_X1 port map( A1 => n67594, A2 => n66509, B1 => n58434, B2 => 
                           n67588, ZN => n63974);
   U49513 : AOI22_X1 port map( A1 => n67594, A2 => n66510, B1 => n58435, B2 => 
                           n67588, ZN => n63954);
   U49514 : AOI22_X1 port map( A1 => n67594, A2 => n66511, B1 => n58436, B2 => 
                           n67588, ZN => n63934);
   U49515 : AOI22_X1 port map( A1 => n67594, A2 => n66512, B1 => n58437, B2 => 
                           n67588, ZN => n63914);
   U49516 : AOI22_X1 port map( A1 => n67594, A2 => n66513, B1 => n58438, B2 => 
                           n67588, ZN => n63894);
   U49517 : OAI22_X1 port map( A1 => n54186, A2 => n67934, B1 => n68238, B2 => 
                           n67928, ZN => n6843);
   U49518 : OAI22_X1 port map( A1 => n54185, A2 => n67934, B1 => n68241, B2 => 
                           n67928, ZN => n6844);
   U49519 : OAI22_X1 port map( A1 => n54184, A2 => n67934, B1 => n68244, B2 => 
                           n67928, ZN => n6845);
   U49520 : OAI22_X1 port map( A1 => n54610, A2 => n67730, B1 => n68240, B2 => 
                           n67724, ZN => n5819);
   U49521 : OAI22_X1 port map( A1 => n54609, A2 => n67730, B1 => n68243, B2 => 
                           n67724, ZN => n5820);
   U49522 : OAI22_X1 port map( A1 => n54608, A2 => n67730, B1 => n68246, B2 => 
                           n67724, ZN => n5821);
   U49523 : OAI22_X1 port map( A1 => n54606, A2 => n67730, B1 => n68249, B2 => 
                           n67724, ZN => n5822);
   U49524 : OAI22_X1 port map( A1 => n67666, A2 => n63862, B1 => n68240, B2 => 
                           n67659, ZN => n5496);
   U49525 : OAI22_X1 port map( A1 => n67666, A2 => n63841, B1 => n68243, B2 => 
                           n67659, ZN => n5498);
   U49526 : OAI22_X1 port map( A1 => n67666, A2 => n63820, B1 => n68246, B2 => 
                           n67659, ZN => n5500);
   U49527 : OAI22_X1 port map( A1 => n67666, A2 => n63765, B1 => n68249, B2 => 
                           n67659, ZN => n5502);
   U49528 : OAI22_X1 port map( A1 => n49229, A2 => n67909, B1 => n68239, B2 => 
                           n67903, ZN => n6715);
   U49529 : OAI22_X1 port map( A1 => n49230, A2 => n67909, B1 => n68242, B2 => 
                           n67903, ZN => n6716);
   U49530 : OAI22_X1 port map( A1 => n49231, A2 => n67909, B1 => n68245, B2 => 
                           n67903, ZN => n6717);
   U49531 : OAI22_X1 port map( A1 => n49228, A2 => n67909, B1 => n68248, B2 => 
                           n67903, ZN => n6718);
   U49532 : OAI22_X1 port map( A1 => n67679, A2 => n63703, B1 => n68240, B2 => 
                           n67672, ZN => n5563);
   U49533 : OAI22_X1 port map( A1 => n67679, A2 => n63702, B1 => n68243, B2 => 
                           n67672, ZN => n5564);
   U49534 : OAI22_X1 port map( A1 => n67679, A2 => n63701, B1 => n68246, B2 => 
                           n67672, ZN => n5565);
   U49535 : OAI22_X1 port map( A1 => n67679, A2 => n63699, B1 => n68249, B2 => 
                           n67672, ZN => n5566);
   U49536 : OAI22_X1 port map( A1 => n8461, A2 => n67893, B1 => n68239, B2 => 
                           n67890, ZN => n6651);
   U49537 : OAI22_X1 port map( A1 => n8477, A2 => n67893, B1 => n68242, B2 => 
                           n67890, ZN => n6652);
   U49538 : OAI22_X1 port map( A1 => n8493, A2 => n67893, B1 => n68245, B2 => 
                           n67890, ZN => n6653);
   U49539 : OAI22_X1 port map( A1 => n8509, A2 => n67893, B1 => n68248, B2 => 
                           n67890, ZN => n6654);
   U49540 : OAI22_X1 port map( A1 => n49480, A2 => n67832, B1 => n68239, B2 => 
                           n67826, ZN => n6331);
   U49541 : OAI22_X1 port map( A1 => n49481, A2 => n67832, B1 => n68242, B2 => 
                           n67826, ZN => n6332);
   U49542 : OAI22_X1 port map( A1 => n49482, A2 => n67832, B1 => n68245, B2 => 
                           n67826, ZN => n6333);
   U49543 : OAI22_X1 port map( A1 => n49483, A2 => n67832, B1 => n68248, B2 => 
                           n67826, ZN => n6334);
   U49544 : OAI22_X1 port map( A1 => n67782, A2 => n63234, B1 => n68239, B2 => 
                           n67775, ZN => n6075);
   U49545 : OAI22_X1 port map( A1 => n67782, A2 => n63233, B1 => n68242, B2 => 
                           n67775, ZN => n6076);
   U49546 : OAI22_X1 port map( A1 => n67782, A2 => n63232, B1 => n68245, B2 => 
                           n67775, ZN => n6077);
   U49547 : OAI22_X1 port map( A1 => n67782, A2 => n63230, B1 => n68248, B2 => 
                           n67775, ZN => n6078);
   U49548 : OAI22_X1 port map( A1 => n8449, A2 => n67794, B1 => n68239, B2 => 
                           n67788, ZN => n6139);
   U49549 : OAI22_X1 port map( A1 => n8465, A2 => n67794, B1 => n68242, B2 => 
                           n67788, ZN => n6140);
   U49550 : OAI22_X1 port map( A1 => n8481, A2 => n67794, B1 => n68245, B2 => 
                           n67788, ZN => n6141);
   U49551 : OAI22_X1 port map( A1 => n8497, A2 => n67794, B1 => n68248, B2 => 
                           n67788, ZN => n6142);
   U49552 : AOI22_X1 port map( A1 => n67416, A2 => n66313, B1 => n67410, B2 => 
                           n58307, ZN => n66282);
   U49553 : AOI22_X1 port map( A1 => n67392, A2 => n58787, B1 => n67386, B2 => 
                           n58439, ZN => n66284);
   U49554 : AOI22_X1 port map( A1 => n67368, A2 => n58036, B1 => n67362, B2 => 
                           n8958, ZN => n66288);
   U49555 : AOI22_X1 port map( A1 => n67416, A2 => n66314, B1 => n67410, B2 => 
                           n58308, ZN => n66258);
   U49556 : AOI22_X1 port map( A1 => n67392, A2 => n58788, B1 => n67386, B2 => 
                           n58440, ZN => n66259);
   U49557 : AOI22_X1 port map( A1 => n67368, A2 => n58001, B1 => n67362, B2 => 
                           n8957, ZN => n66260);
   U49558 : AOI22_X1 port map( A1 => n67416, A2 => n66315, B1 => n67410, B2 => 
                           n58309, ZN => n66240);
   U49559 : AOI22_X1 port map( A1 => n67392, A2 => n58789, B1 => n67386, B2 => 
                           n58441, ZN => n66241);
   U49560 : AOI22_X1 port map( A1 => n67368, A2 => n57977, B1 => n67362, B2 => 
                           n8956, ZN => n66242);
   U49561 : AOI22_X1 port map( A1 => n67416, A2 => n66316, B1 => n67410, B2 => 
                           n58310, ZN => n66222);
   U49562 : AOI22_X1 port map( A1 => n67392, A2 => n58790, B1 => n67386, B2 => 
                           n58442, ZN => n66223);
   U49563 : AOI22_X1 port map( A1 => n67368, A2 => n57953, B1 => n67362, B2 => 
                           n8955, ZN => n66224);
   U49564 : AOI22_X1 port map( A1 => n67416, A2 => n66317, B1 => n67410, B2 => 
                           n58311, ZN => n66204);
   U49565 : AOI22_X1 port map( A1 => n67392, A2 => n58791, B1 => n67386, B2 => 
                           n58443, ZN => n66205);
   U49566 : AOI22_X1 port map( A1 => n67368, A2 => n57929, B1 => n67362, B2 => 
                           n8954, ZN => n66206);
   U49567 : AOI22_X1 port map( A1 => n67416, A2 => n66318, B1 => n67410, B2 => 
                           n58312, ZN => n66186);
   U49568 : AOI22_X1 port map( A1 => n67392, A2 => n58792, B1 => n67386, B2 => 
                           n58444, ZN => n66187);
   U49569 : AOI22_X1 port map( A1 => n67368, A2 => n57905, B1 => n67362, B2 => 
                           n8953, ZN => n66188);
   U49570 : AOI22_X1 port map( A1 => n67416, A2 => n66319, B1 => n67410, B2 => 
                           n58313, ZN => n66168);
   U49571 : AOI22_X1 port map( A1 => n67392, A2 => n58793, B1 => n67386, B2 => 
                           n58445, ZN => n66169);
   U49572 : AOI22_X1 port map( A1 => n67368, A2 => n57881, B1 => n67362, B2 => 
                           n8952, ZN => n66170);
   U49573 : AOI22_X1 port map( A1 => n67416, A2 => n66320, B1 => n67410, B2 => 
                           n58314, ZN => n66150);
   U49574 : AOI22_X1 port map( A1 => n67392, A2 => n58794, B1 => n67386, B2 => 
                           n58446, ZN => n66151);
   U49575 : AOI22_X1 port map( A1 => n67368, A2 => n57857, B1 => n67362, B2 => 
                           n8951, ZN => n66152);
   U49576 : AOI22_X1 port map( A1 => n67416, A2 => n66321, B1 => n67410, B2 => 
                           n58315, ZN => n66132);
   U49577 : AOI22_X1 port map( A1 => n67392, A2 => n58795, B1 => n67386, B2 => 
                           n58447, ZN => n66133);
   U49578 : AOI22_X1 port map( A1 => n67368, A2 => n57833, B1 => n67362, B2 => 
                           n8950, ZN => n66134);
   U49579 : AOI22_X1 port map( A1 => n67416, A2 => n66322, B1 => n67410, B2 => 
                           n58316, ZN => n66114);
   U49580 : AOI22_X1 port map( A1 => n67392, A2 => n58796, B1 => n67386, B2 => 
                           n58448, ZN => n66115);
   U49581 : AOI22_X1 port map( A1 => n67368, A2 => n57809, B1 => n67362, B2 => 
                           n8949, ZN => n66116);
   U49582 : AOI22_X1 port map( A1 => n67416, A2 => n66323, B1 => n67410, B2 => 
                           n58317, ZN => n66096);
   U49583 : AOI22_X1 port map( A1 => n67392, A2 => n58797, B1 => n67386, B2 => 
                           n58449, ZN => n66097);
   U49584 : AOI22_X1 port map( A1 => n67368, A2 => n57785, B1 => n67362, B2 => 
                           n8948, ZN => n66098);
   U49585 : AOI22_X1 port map( A1 => n67416, A2 => n66324, B1 => n67410, B2 => 
                           n58318, ZN => n66078);
   U49586 : AOI22_X1 port map( A1 => n67392, A2 => n58798, B1 => n67386, B2 => 
                           n58450, ZN => n66079);
   U49587 : AOI22_X1 port map( A1 => n67368, A2 => n57761, B1 => n67362, B2 => 
                           n8947, ZN => n66080);
   U49588 : AOI22_X1 port map( A1 => n67441, A2 => n58391, B1 => n67435, B2 => 
                           OUT2_12_port, ZN => n66059);
   U49589 : AOI22_X1 port map( A1 => n67393, A2 => n56101, B1 => n67387, B2 => 
                           n58451, ZN => n66061);
   U49590 : AOI22_X1 port map( A1 => n67369, A2 => n57737, B1 => n67363, B2 => 
                           n8946, ZN => n66062);
   U49591 : AOI22_X1 port map( A1 => n67441, A2 => n58392, B1 => n67435, B2 => 
                           OUT2_13_port, ZN => n66041);
   U49592 : AOI22_X1 port map( A1 => n67393, A2 => n56074, B1 => n67387, B2 => 
                           n58452, ZN => n66043);
   U49593 : AOI22_X1 port map( A1 => n67369, A2 => n57713, B1 => n67363, B2 => 
                           n8945, ZN => n66044);
   U49594 : AOI22_X1 port map( A1 => n67441, A2 => n58393, B1 => n67435, B2 => 
                           OUT2_14_port, ZN => n66023);
   U49595 : AOI22_X1 port map( A1 => n67393, A2 => n56047, B1 => n67387, B2 => 
                           n58453, ZN => n66025);
   U49596 : AOI22_X1 port map( A1 => n67369, A2 => n57689, B1 => n67363, B2 => 
                           n8944, ZN => n66026);
   U49597 : AOI22_X1 port map( A1 => n67441, A2 => n58394, B1 => n67435, B2 => 
                           OUT2_15_port, ZN => n66005);
   U49598 : AOI22_X1 port map( A1 => n67393, A2 => n56020, B1 => n67387, B2 => 
                           n58454, ZN => n66007);
   U49599 : AOI22_X1 port map( A1 => n67369, A2 => n57665, B1 => n67363, B2 => 
                           n8943, ZN => n66008);
   U49600 : AOI22_X1 port map( A1 => n67441, A2 => n58395, B1 => n67435, B2 => 
                           OUT2_16_port, ZN => n65987);
   U49601 : AOI22_X1 port map( A1 => n67393, A2 => n58799, B1 => n67387, B2 => 
                           n58455, ZN => n65989);
   U49602 : AOI22_X1 port map( A1 => n67369, A2 => n57641, B1 => n67363, B2 => 
                           n8942, ZN => n65990);
   U49603 : AOI22_X1 port map( A1 => n67441, A2 => n58396, B1 => n67435, B2 => 
                           OUT2_17_port, ZN => n65969);
   U49604 : AOI22_X1 port map( A1 => n67393, A2 => n58800, B1 => n67387, B2 => 
                           n58456, ZN => n65971);
   U49605 : AOI22_X1 port map( A1 => n67369, A2 => n57617, B1 => n67363, B2 => 
                           n8941, ZN => n65972);
   U49606 : AOI22_X1 port map( A1 => n67441, A2 => n58397, B1 => n67435, B2 => 
                           OUT2_18_port, ZN => n65951);
   U49607 : AOI22_X1 port map( A1 => n67393, A2 => n58801, B1 => n67387, B2 => 
                           n58457, ZN => n65953);
   U49608 : AOI22_X1 port map( A1 => n67369, A2 => n57593, B1 => n67363, B2 => 
                           n8940, ZN => n65954);
   U49609 : AOI22_X1 port map( A1 => n67441, A2 => n58398, B1 => n67435, B2 => 
                           OUT2_19_port, ZN => n65933);
   U49610 : AOI22_X1 port map( A1 => n67393, A2 => n58802, B1 => n67387, B2 => 
                           n58458, ZN => n65935);
   U49611 : AOI22_X1 port map( A1 => n67369, A2 => n57569, B1 => n67363, B2 => 
                           n8939, ZN => n65936);
   U49612 : AOI22_X1 port map( A1 => n67441, A2 => n58399, B1 => n67435, B2 => 
                           OUT2_20_port, ZN => n65915);
   U49613 : AOI22_X1 port map( A1 => n67393, A2 => n58803, B1 => n67387, B2 => 
                           n58459, ZN => n65917);
   U49614 : AOI22_X1 port map( A1 => n67369, A2 => n57545, B1 => n67363, B2 => 
                           n8938, ZN => n65918);
   U49615 : AOI22_X1 port map( A1 => n67441, A2 => n58400, B1 => n67435, B2 => 
                           OUT2_21_port, ZN => n65897);
   U49616 : AOI22_X1 port map( A1 => n67393, A2 => n58804, B1 => n67387, B2 => 
                           n58460, ZN => n65899);
   U49617 : AOI22_X1 port map( A1 => n67369, A2 => n57521, B1 => n67363, B2 => 
                           n8937, ZN => n65900);
   U49618 : AOI22_X1 port map( A1 => n67441, A2 => n58401, B1 => n67436, B2 => 
                           OUT2_22_port, ZN => n65879);
   U49619 : AOI22_X1 port map( A1 => n67393, A2 => n58805, B1 => n67387, B2 => 
                           n58461, ZN => n65881);
   U49620 : AOI22_X1 port map( A1 => n67369, A2 => n57497, B1 => n67363, B2 => 
                           n8936, ZN => n65882);
   U49621 : AOI22_X1 port map( A1 => n67441, A2 => n58402, B1 => n67436, B2 => 
                           OUT2_23_port, ZN => n65861);
   U49622 : AOI22_X1 port map( A1 => n67393, A2 => n58806, B1 => n67387, B2 => 
                           n58462, ZN => n65863);
   U49623 : AOI22_X1 port map( A1 => n67369, A2 => n57473, B1 => n67363, B2 => 
                           n8935, ZN => n65864);
   U49624 : AOI22_X1 port map( A1 => n67442, A2 => n58403, B1 => n67436, B2 => 
                           OUT2_24_port, ZN => n65843);
   U49625 : AOI22_X1 port map( A1 => n67394, A2 => n58807, B1 => n67388, B2 => 
                           n58463, ZN => n65845);
   U49626 : AOI22_X1 port map( A1 => n67370, A2 => n57449, B1 => n67364, B2 => 
                           n8934, ZN => n65846);
   U49627 : AOI22_X1 port map( A1 => n67442, A2 => n58404, B1 => n67436, B2 => 
                           OUT2_25_port, ZN => n65825);
   U49628 : AOI22_X1 port map( A1 => n67394, A2 => n58808, B1 => n67388, B2 => 
                           n58464, ZN => n65827);
   U49629 : AOI22_X1 port map( A1 => n67370, A2 => n57425, B1 => n67364, B2 => 
                           n8933, ZN => n65828);
   U49630 : AOI22_X1 port map( A1 => n67442, A2 => n58405, B1 => n67436, B2 => 
                           OUT2_26_port, ZN => n65807);
   U49631 : AOI22_X1 port map( A1 => n67394, A2 => n58809, B1 => n67388, B2 => 
                           n58465, ZN => n65809);
   U49632 : AOI22_X1 port map( A1 => n67370, A2 => n57401, B1 => n67364, B2 => 
                           n8932, ZN => n65810);
   U49633 : AOI22_X1 port map( A1 => n67442, A2 => n58406, B1 => n67436, B2 => 
                           OUT2_27_port, ZN => n65789);
   U49634 : AOI22_X1 port map( A1 => n67394, A2 => n58810, B1 => n67388, B2 => 
                           n58466, ZN => n65791);
   U49635 : AOI22_X1 port map( A1 => n67370, A2 => n57377, B1 => n67364, B2 => 
                           n8931, ZN => n65792);
   U49636 : AOI22_X1 port map( A1 => n67442, A2 => n58407, B1 => n67436, B2 => 
                           OUT2_28_port, ZN => n65771);
   U49637 : AOI22_X1 port map( A1 => n67394, A2 => n58811, B1 => n67388, B2 => 
                           n58467, ZN => n65773);
   U49638 : AOI22_X1 port map( A1 => n67370, A2 => n57353, B1 => n67364, B2 => 
                           n8930, ZN => n65774);
   U49639 : AOI22_X1 port map( A1 => n67442, A2 => n58408, B1 => n67436, B2 => 
                           OUT2_29_port, ZN => n65753);
   U49640 : AOI22_X1 port map( A1 => n67394, A2 => n58812, B1 => n67388, B2 => 
                           n58468, ZN => n65755);
   U49641 : AOI22_X1 port map( A1 => n67370, A2 => n57329, B1 => n67364, B2 => 
                           n8929, ZN => n65756);
   U49642 : AOI22_X1 port map( A1 => n67442, A2 => n58409, B1 => n67436, B2 => 
                           OUT2_30_port, ZN => n65735);
   U49643 : AOI22_X1 port map( A1 => n67394, A2 => n58813, B1 => n67388, B2 => 
                           n58469, ZN => n65737);
   U49644 : AOI22_X1 port map( A1 => n67370, A2 => n57305, B1 => n67364, B2 => 
                           n8928, ZN => n65738);
   U49645 : AOI22_X1 port map( A1 => n67442, A2 => n58410, B1 => n67436, B2 => 
                           OUT2_31_port, ZN => n65717);
   U49646 : AOI22_X1 port map( A1 => n67394, A2 => n58814, B1 => n67388, B2 => 
                           n58470, ZN => n65719);
   U49647 : AOI22_X1 port map( A1 => n67370, A2 => n57281, B1 => n67364, B2 => 
                           n8927, ZN => n65720);
   U49648 : AOI22_X1 port map( A1 => n67442, A2 => n58411, B1 => n67436, B2 => 
                           OUT2_32_port, ZN => n65699);
   U49649 : AOI22_X1 port map( A1 => n67394, A2 => n58815, B1 => n67388, B2 => 
                           n58471, ZN => n65701);
   U49650 : AOI22_X1 port map( A1 => n67370, A2 => n57257, B1 => n67364, B2 => 
                           n8926, ZN => n65702);
   U49651 : AOI22_X1 port map( A1 => n67442, A2 => n58412, B1 => n67436, B2 => 
                           OUT2_33_port, ZN => n65681);
   U49652 : AOI22_X1 port map( A1 => n67394, A2 => n58816, B1 => n67388, B2 => 
                           n58472, ZN => n65683);
   U49653 : AOI22_X1 port map( A1 => n67370, A2 => n57233, B1 => n67364, B2 => 
                           n8925, ZN => n65684);
   U49654 : AOI22_X1 port map( A1 => n67442, A2 => n58413, B1 => n67436, B2 => 
                           OUT2_34_port, ZN => n65663);
   U49655 : AOI22_X1 port map( A1 => n67394, A2 => n58817, B1 => n67388, B2 => 
                           n58473, ZN => n65665);
   U49656 : AOI22_X1 port map( A1 => n67370, A2 => n57209, B1 => n67364, B2 => 
                           n8924, ZN => n65666);
   U49657 : AOI22_X1 port map( A1 => n67442, A2 => n58414, B1 => n67437, B2 => 
                           OUT2_35_port, ZN => n65645);
   U49658 : AOI22_X1 port map( A1 => n67394, A2 => n58818, B1 => n67388, B2 => 
                           n58474, ZN => n65647);
   U49659 : AOI22_X1 port map( A1 => n67370, A2 => n57185, B1 => n67364, B2 => 
                           n8923, ZN => n65648);
   U49660 : AOI22_X1 port map( A1 => n67443, A2 => n58415, B1 => n67437, B2 => 
                           OUT2_36_port, ZN => n65627);
   U49661 : AOI22_X1 port map( A1 => n67395, A2 => n58819, B1 => n67389, B2 => 
                           n58475, ZN => n65629);
   U49662 : AOI22_X1 port map( A1 => n67371, A2 => n57161, B1 => n67365, B2 => 
                           n8922, ZN => n65630);
   U49663 : AOI22_X1 port map( A1 => n67443, A2 => n58416, B1 => n67437, B2 => 
                           OUT2_37_port, ZN => n65609);
   U49664 : AOI22_X1 port map( A1 => n67395, A2 => n58820, B1 => n67389, B2 => 
                           n58476, ZN => n65611);
   U49665 : AOI22_X1 port map( A1 => n67371, A2 => n57137, B1 => n67365, B2 => 
                           n8921, ZN => n65612);
   U49666 : AOI22_X1 port map( A1 => n67443, A2 => n58417, B1 => n67437, B2 => 
                           OUT2_38_port, ZN => n65591);
   U49667 : AOI22_X1 port map( A1 => n67395, A2 => n58821, B1 => n67389, B2 => 
                           n58477, ZN => n65593);
   U49668 : AOI22_X1 port map( A1 => n67371, A2 => n57113, B1 => n67365, B2 => 
                           n8920, ZN => n65594);
   U49669 : AOI22_X1 port map( A1 => n67443, A2 => n58418, B1 => n67437, B2 => 
                           OUT2_39_port, ZN => n65573);
   U49670 : AOI22_X1 port map( A1 => n67395, A2 => n58822, B1 => n67389, B2 => 
                           n58478, ZN => n65575);
   U49671 : AOI22_X1 port map( A1 => n67371, A2 => n57089, B1 => n67365, B2 => 
                           n8919, ZN => n65576);
   U49672 : AOI22_X1 port map( A1 => n67443, A2 => n58419, B1 => n67437, B2 => 
                           OUT2_40_port, ZN => n65555);
   U49673 : AOI22_X1 port map( A1 => n67395, A2 => n58823, B1 => n67389, B2 => 
                           n58479, ZN => n65557);
   U49674 : AOI22_X1 port map( A1 => n67371, A2 => n57065, B1 => n67365, B2 => 
                           n8918, ZN => n65558);
   U49675 : AOI22_X1 port map( A1 => n67443, A2 => n58420, B1 => n67437, B2 => 
                           OUT2_41_port, ZN => n65537);
   U49676 : AOI22_X1 port map( A1 => n67395, A2 => n58824, B1 => n67389, B2 => 
                           n58480, ZN => n65539);
   U49677 : AOI22_X1 port map( A1 => n67371, A2 => n57041, B1 => n67365, B2 => 
                           n8917, ZN => n65540);
   U49678 : AOI22_X1 port map( A1 => n67443, A2 => n58421, B1 => n67437, B2 => 
                           OUT2_42_port, ZN => n65519);
   U49679 : AOI22_X1 port map( A1 => n67395, A2 => n58825, B1 => n67389, B2 => 
                           n58481, ZN => n65521);
   U49680 : AOI22_X1 port map( A1 => n67371, A2 => n57017, B1 => n67365, B2 => 
                           n8916, ZN => n65522);
   U49681 : AOI22_X1 port map( A1 => n67443, A2 => n58422, B1 => n67437, B2 => 
                           OUT2_43_port, ZN => n65501);
   U49682 : AOI22_X1 port map( A1 => n67395, A2 => n58826, B1 => n67389, B2 => 
                           n58482, ZN => n65503);
   U49683 : AOI22_X1 port map( A1 => n67371, A2 => n56993, B1 => n67365, B2 => 
                           n8915, ZN => n65504);
   U49684 : AOI22_X1 port map( A1 => n67443, A2 => n58423, B1 => n67437, B2 => 
                           OUT2_44_port, ZN => n65483);
   U49685 : AOI22_X1 port map( A1 => n67395, A2 => n58827, B1 => n67389, B2 => 
                           n58483, ZN => n65485);
   U49686 : AOI22_X1 port map( A1 => n67371, A2 => n56969, B1 => n67365, B2 => 
                           n8914, ZN => n65486);
   U49687 : AOI22_X1 port map( A1 => n67443, A2 => n58424, B1 => n67437, B2 => 
                           OUT2_45_port, ZN => n65465);
   U49688 : AOI22_X1 port map( A1 => n67395, A2 => n58828, B1 => n67389, B2 => 
                           n58484, ZN => n65467);
   U49689 : AOI22_X1 port map( A1 => n67371, A2 => n56945, B1 => n67365, B2 => 
                           n8913, ZN => n65468);
   U49690 : AOI22_X1 port map( A1 => n67443, A2 => n58425, B1 => n67437, B2 => 
                           OUT2_46_port, ZN => n65447);
   U49691 : AOI22_X1 port map( A1 => n67395, A2 => n58829, B1 => n67389, B2 => 
                           n58485, ZN => n65449);
   U49692 : AOI22_X1 port map( A1 => n67371, A2 => n56921, B1 => n67365, B2 => 
                           n8912, ZN => n65450);
   U49693 : AOI22_X1 port map( A1 => n67443, A2 => n58426, B1 => n67437, B2 => 
                           OUT2_47_port, ZN => n65429);
   U49694 : AOI22_X1 port map( A1 => n67395, A2 => n58830, B1 => n67389, B2 => 
                           n58486, ZN => n65431);
   U49695 : AOI22_X1 port map( A1 => n67371, A2 => n56897, B1 => n67365, B2 => 
                           n8911, ZN => n65432);
   U49696 : AOI22_X1 port map( A1 => n67444, A2 => n58427, B1 => n67438, B2 => 
                           OUT2_48_port, ZN => n65411);
   U49697 : AOI22_X1 port map( A1 => n67396, A2 => n58831, B1 => n67390, B2 => 
                           n58487, ZN => n65413);
   U49698 : AOI22_X1 port map( A1 => n67372, A2 => n56873, B1 => n67366, B2 => 
                           n8910, ZN => n65414);
   U49699 : AOI22_X1 port map( A1 => n67444, A2 => n58428, B1 => n67438, B2 => 
                           OUT2_49_port, ZN => n65393);
   U49700 : AOI22_X1 port map( A1 => n67396, A2 => n58832, B1 => n67390, B2 => 
                           n58488, ZN => n65395);
   U49701 : AOI22_X1 port map( A1 => n67372, A2 => n56849, B1 => n67366, B2 => 
                           n8909, ZN => n65396);
   U49702 : AOI22_X1 port map( A1 => n67444, A2 => n58429, B1 => n67438, B2 => 
                           OUT2_50_port, ZN => n65375);
   U49703 : AOI22_X1 port map( A1 => n67396, A2 => n58833, B1 => n67390, B2 => 
                           n58489, ZN => n65377);
   U49704 : AOI22_X1 port map( A1 => n67372, A2 => n56825, B1 => n67366, B2 => 
                           n8908, ZN => n65378);
   U49705 : AOI22_X1 port map( A1 => n67444, A2 => n58430, B1 => n67438, B2 => 
                           OUT2_51_port, ZN => n65357);
   U49706 : AOI22_X1 port map( A1 => n67396, A2 => n58834, B1 => n67390, B2 => 
                           n58490, ZN => n65359);
   U49707 : AOI22_X1 port map( A1 => n67372, A2 => n56801, B1 => n67366, B2 => 
                           n8907, ZN => n65360);
   U49708 : AOI22_X1 port map( A1 => n67444, A2 => n58431, B1 => n67438, B2 => 
                           OUT2_52_port, ZN => n65339);
   U49709 : AOI22_X1 port map( A1 => n67396, A2 => n58835, B1 => n67390, B2 => 
                           n58491, ZN => n65341);
   U49710 : AOI22_X1 port map( A1 => n67372, A2 => n56777, B1 => n67366, B2 => 
                           n8906, ZN => n65342);
   U49711 : AOI22_X1 port map( A1 => n67444, A2 => n58432, B1 => n67438, B2 => 
                           OUT2_53_port, ZN => n65321);
   U49712 : AOI22_X1 port map( A1 => n67396, A2 => n58836, B1 => n67390, B2 => 
                           n58492, ZN => n65323);
   U49713 : AOI22_X1 port map( A1 => n67372, A2 => n56753, B1 => n67366, B2 => 
                           n8905, ZN => n65324);
   U49714 : AOI22_X1 port map( A1 => n67444, A2 => n58433, B1 => n67438, B2 => 
                           OUT2_54_port, ZN => n65303);
   U49715 : AOI22_X1 port map( A1 => n67396, A2 => n58837, B1 => n67390, B2 => 
                           n58493, ZN => n65305);
   U49716 : AOI22_X1 port map( A1 => n67372, A2 => n56729, B1 => n67366, B2 => 
                           n8904, ZN => n65306);
   U49717 : AOI22_X1 port map( A1 => n67444, A2 => n58434, B1 => n67438, B2 => 
                           OUT2_55_port, ZN => n65285);
   U49718 : AOI22_X1 port map( A1 => n67396, A2 => n58838, B1 => n67390, B2 => 
                           n58494, ZN => n65287);
   U49719 : AOI22_X1 port map( A1 => n67372, A2 => n56705, B1 => n67366, B2 => 
                           n8903, ZN => n65288);
   U49720 : AOI22_X1 port map( A1 => n67444, A2 => n58435, B1 => n67438, B2 => 
                           OUT2_56_port, ZN => n65267);
   U49721 : AOI22_X1 port map( A1 => n67396, A2 => n58839, B1 => n67390, B2 => 
                           n58495, ZN => n65269);
   U49722 : AOI22_X1 port map( A1 => n67372, A2 => n56681, B1 => n67366, B2 => 
                           n8902, ZN => n65270);
   U49723 : AOI22_X1 port map( A1 => n67444, A2 => n58436, B1 => n67438, B2 => 
                           OUT2_57_port, ZN => n65249);
   U49724 : AOI22_X1 port map( A1 => n67396, A2 => n58840, B1 => n67390, B2 => 
                           n58496, ZN => n65251);
   U49725 : AOI22_X1 port map( A1 => n67372, A2 => n56657, B1 => n67366, B2 => 
                           n8901, ZN => n65252);
   U49726 : AOI22_X1 port map( A1 => n67444, A2 => n58437, B1 => n67438, B2 => 
                           OUT2_58_port, ZN => n65231);
   U49727 : AOI22_X1 port map( A1 => n67396, A2 => n58841, B1 => n67390, B2 => 
                           n58497, ZN => n65233);
   U49728 : AOI22_X1 port map( A1 => n67372, A2 => n56633, B1 => n67366, B2 => 
                           n8900, ZN => n65234);
   U49729 : AOI22_X1 port map( A1 => n67444, A2 => n58438, B1 => n67438, B2 => 
                           OUT2_59_port, ZN => n65213);
   U49730 : AOI22_X1 port map( A1 => n67396, A2 => n58842, B1 => n67390, B2 => 
                           n58498, ZN => n65215);
   U49731 : AOI22_X1 port map( A1 => n67372, A2 => n56609, B1 => n67366, B2 => 
                           n8899, ZN => n65216);
   U49732 : AOI22_X1 port map( A1 => n67590, A2 => n65084, B1 => n58379, B2 => 
                           n67584, ZN => n65083);
   U49733 : AOI22_X1 port map( A1 => n67636, A2 => n58013, B1 => n67632, B2 => 
                           OUT1_0_port, ZN => n65072);
   U49734 : AOI22_X1 port map( A1 => n67614, A2 => n58627, B1 => n67608, B2 => 
                           n58731, ZN => n65079);
   U49735 : AOI22_X1 port map( A1 => n67590, A2 => n65055, B1 => n58380, B2 => 
                           n67584, ZN => n65054);
   U49736 : AOI22_X1 port map( A1 => n67636, A2 => n57989, B1 => n67632, B2 => 
                           OUT1_1_port, ZN => n65052);
   U49737 : AOI22_X1 port map( A1 => n67614, A2 => n58628, B1 => n67608, B2 => 
                           n58732, ZN => n65053);
   U49738 : AOI22_X1 port map( A1 => n67590, A2 => n65035, B1 => n58381, B2 => 
                           n67584, ZN => n65034);
   U49739 : AOI22_X1 port map( A1 => n67636, A2 => n57965, B1 => n67632, B2 => 
                           OUT1_2_port, ZN => n65032);
   U49740 : AOI22_X1 port map( A1 => n67614, A2 => n58629, B1 => n67608, B2 => 
                           n58733, ZN => n65033);
   U49741 : AOI22_X1 port map( A1 => n67590, A2 => n65015, B1 => n58382, B2 => 
                           n67584, ZN => n65014);
   U49742 : AOI22_X1 port map( A1 => n67636, A2 => n57941, B1 => n67632, B2 => 
                           OUT1_3_port, ZN => n65012);
   U49743 : AOI22_X1 port map( A1 => n67614, A2 => n58630, B1 => n67608, B2 => 
                           n58734, ZN => n65013);
   U49744 : AOI22_X1 port map( A1 => n67590, A2 => n64995, B1 => n58383, B2 => 
                           n67584, ZN => n64994);
   U49745 : AOI22_X1 port map( A1 => n67636, A2 => n57917, B1 => n67632, B2 => 
                           OUT1_4_port, ZN => n64992);
   U49746 : AOI22_X1 port map( A1 => n67614, A2 => n58631, B1 => n67608, B2 => 
                           n58735, ZN => n64993);
   U49747 : AOI22_X1 port map( A1 => n67590, A2 => n64975, B1 => n58384, B2 => 
                           n67584, ZN => n64974);
   U49748 : AOI22_X1 port map( A1 => n67636, A2 => n57893, B1 => n67632, B2 => 
                           OUT1_5_port, ZN => n64972);
   U49749 : AOI22_X1 port map( A1 => n67614, A2 => n58632, B1 => n67608, B2 => 
                           n58736, ZN => n64973);
   U49750 : AOI22_X1 port map( A1 => n67590, A2 => n64955, B1 => n58385, B2 => 
                           n67584, ZN => n64954);
   U49751 : AOI22_X1 port map( A1 => n67636, A2 => n57869, B1 => n67632, B2 => 
                           OUT1_6_port, ZN => n64952);
   U49752 : AOI22_X1 port map( A1 => n67614, A2 => n58633, B1 => n67608, B2 => 
                           n58737, ZN => n64953);
   U49753 : AOI22_X1 port map( A1 => n67590, A2 => n64935, B1 => n58386, B2 => 
                           n67584, ZN => n64934);
   U49754 : AOI22_X1 port map( A1 => n67636, A2 => n57845, B1 => n67632, B2 => 
                           OUT1_7_port, ZN => n64932);
   U49755 : AOI22_X1 port map( A1 => n67614, A2 => n58634, B1 => n67608, B2 => 
                           n58738, ZN => n64933);
   U49756 : AOI22_X1 port map( A1 => n67590, A2 => n64915, B1 => n58387, B2 => 
                           n67584, ZN => n64914);
   U49757 : AOI22_X1 port map( A1 => n67636, A2 => n57821, B1 => n67632, B2 => 
                           OUT1_8_port, ZN => n64912);
   U49758 : AOI22_X1 port map( A1 => n67614, A2 => n58635, B1 => n67608, B2 => 
                           n58739, ZN => n64913);
   U49759 : AOI22_X1 port map( A1 => n67590, A2 => n64895, B1 => n58388, B2 => 
                           n67584, ZN => n64894);
   U49760 : AOI22_X1 port map( A1 => n67636, A2 => n57797, B1 => n67632, B2 => 
                           OUT1_9_port, ZN => n64892);
   U49761 : AOI22_X1 port map( A1 => n67614, A2 => n58636, B1 => n67608, B2 => 
                           n58740, ZN => n64893);
   U49762 : AOI22_X1 port map( A1 => n67590, A2 => n64875, B1 => n58389, B2 => 
                           n67584, ZN => n64874);
   U49763 : AOI22_X1 port map( A1 => n67636, A2 => n57773, B1 => n67632, B2 => 
                           OUT1_10_port, ZN => n64872);
   U49764 : AOI22_X1 port map( A1 => n67614, A2 => n58637, B1 => n67608, B2 => 
                           n58741, ZN => n64873);
   U49765 : AOI22_X1 port map( A1 => n67590, A2 => n64855, B1 => n58390, B2 => 
                           n67584, ZN => n64854);
   U49766 : AOI22_X1 port map( A1 => n67636, A2 => n57749, B1 => n67634, B2 => 
                           OUT1_11_port, ZN => n64852);
   U49767 : AOI22_X1 port map( A1 => n67614, A2 => n58638, B1 => n67608, B2 => 
                           n58742, ZN => n64853);
   U49768 : AOI22_X1 port map( A1 => n67567, A2 => n9061, B1 => n67561, B2 => 
                           n57737, ZN => n64836);
   U49769 : AOI22_X1 port map( A1 => n67591, A2 => n66514, B1 => n58391, B2 => 
                           n67585, ZN => n64834);
   U49770 : AOI22_X1 port map( A1 => n67615, A2 => n58639, B1 => n67609, B2 => 
                           n58667, ZN => n64833);
   U49771 : AOI22_X1 port map( A1 => n67567, A2 => n9059, B1 => n67561, B2 => 
                           n57713, ZN => n64816);
   U49772 : AOI22_X1 port map( A1 => n67591, A2 => n66515, B1 => n58392, B2 => 
                           n67585, ZN => n64814);
   U49773 : AOI22_X1 port map( A1 => n67615, A2 => n58640, B1 => n67609, B2 => 
                           n58668, ZN => n64813);
   U49774 : AOI22_X1 port map( A1 => n67567, A2 => n9057, B1 => n67561, B2 => 
                           n57689, ZN => n64796);
   U49775 : AOI22_X1 port map( A1 => n67591, A2 => n66516, B1 => n58393, B2 => 
                           n67585, ZN => n64794);
   U49776 : AOI22_X1 port map( A1 => n67615, A2 => n58641, B1 => n67609, B2 => 
                           n58669, ZN => n64793);
   U49777 : AOI22_X1 port map( A1 => n67567, A2 => n9055, B1 => n67561, B2 => 
                           n57665, ZN => n64776);
   U49778 : AOI22_X1 port map( A1 => n67591, A2 => n66517, B1 => n58394, B2 => 
                           n67585, ZN => n64774);
   U49779 : AOI22_X1 port map( A1 => n67615, A2 => n58642, B1 => n67609, B2 => 
                           n58670, ZN => n64773);
   U49780 : AOI22_X1 port map( A1 => n67567, A2 => n9053, B1 => n67561, B2 => 
                           n57641, ZN => n64756);
   U49781 : AOI22_X1 port map( A1 => n67591, A2 => n66518, B1 => n58395, B2 => 
                           n67585, ZN => n64754);
   U49782 : AOI22_X1 port map( A1 => n67615, A2 => n57631, B1 => n67609, B2 => 
                           n58671, ZN => n64753);
   U49783 : AOI22_X1 port map( A1 => n67567, A2 => n9051, B1 => n67561, B2 => 
                           n57617, ZN => n64736);
   U49784 : AOI22_X1 port map( A1 => n67591, A2 => n66519, B1 => n58396, B2 => 
                           n67585, ZN => n64734);
   U49785 : AOI22_X1 port map( A1 => n67615, A2 => n57607, B1 => n67609, B2 => 
                           n58672, ZN => n64733);
   U49786 : AOI22_X1 port map( A1 => n67567, A2 => n9049, B1 => n67561, B2 => 
                           n57593, ZN => n64716);
   U49787 : AOI22_X1 port map( A1 => n67591, A2 => n66520, B1 => n58397, B2 => 
                           n67585, ZN => n64714);
   U49788 : AOI22_X1 port map( A1 => n67615, A2 => n57583, B1 => n67609, B2 => 
                           n58673, ZN => n64713);
   U49789 : AOI22_X1 port map( A1 => n67567, A2 => n9047, B1 => n67561, B2 => 
                           n57569, ZN => n64696);
   U49790 : AOI22_X1 port map( A1 => n67591, A2 => n66521, B1 => n58398, B2 => 
                           n67585, ZN => n64694);
   U49791 : AOI22_X1 port map( A1 => n67615, A2 => n57559, B1 => n67609, B2 => 
                           n58674, ZN => n64693);
   U49792 : AOI22_X1 port map( A1 => n67567, A2 => n9045, B1 => n67561, B2 => 
                           n57545, ZN => n64676);
   U49793 : AOI22_X1 port map( A1 => n67591, A2 => n66522, B1 => n58399, B2 => 
                           n67585, ZN => n64674);
   U49794 : AOI22_X1 port map( A1 => n67615, A2 => n57535, B1 => n67609, B2 => 
                           n58675, ZN => n64673);
   U49795 : AOI22_X1 port map( A1 => n67567, A2 => n9043, B1 => n67561, B2 => 
                           n57521, ZN => n64656);
   U49796 : AOI22_X1 port map( A1 => n67591, A2 => n66523, B1 => n58400, B2 => 
                           n67585, ZN => n64654);
   U49797 : AOI22_X1 port map( A1 => n67615, A2 => n57511, B1 => n67609, B2 => 
                           n58676, ZN => n64653);
   U49798 : AOI22_X1 port map( A1 => n67567, A2 => n9041, B1 => n67561, B2 => 
                           n57497, ZN => n64636);
   U49799 : AOI22_X1 port map( A1 => n67591, A2 => n66524, B1 => n58401, B2 => 
                           n67585, ZN => n64634);
   U49800 : AOI22_X1 port map( A1 => n67615, A2 => n57487, B1 => n67609, B2 => 
                           n58677, ZN => n64633);
   U49801 : AOI22_X1 port map( A1 => n67567, A2 => n9039, B1 => n67561, B2 => 
                           n57473, ZN => n64616);
   U49802 : AOI22_X1 port map( A1 => n67591, A2 => n66525, B1 => n58402, B2 => 
                           n67585, ZN => n64614);
   U49803 : AOI22_X1 port map( A1 => n67615, A2 => n57463, B1 => n67609, B2 => 
                           n58678, ZN => n64613);
   U49804 : AOI22_X1 port map( A1 => n67568, A2 => n9037, B1 => n67562, B2 => 
                           n57449, ZN => n64596);
   U49805 : AOI22_X1 port map( A1 => n67592, A2 => n66526, B1 => n58403, B2 => 
                           n67586, ZN => n64594);
   U49806 : AOI22_X1 port map( A1 => n67616, A2 => n57439, B1 => n67610, B2 => 
                           n58679, ZN => n64593);
   U49807 : AOI22_X1 port map( A1 => n67568, A2 => n9035, B1 => n67562, B2 => 
                           n57425, ZN => n64576);
   U49808 : AOI22_X1 port map( A1 => n67592, A2 => n66527, B1 => n58404, B2 => 
                           n67586, ZN => n64574);
   U49809 : AOI22_X1 port map( A1 => n67616, A2 => n57415, B1 => n67610, B2 => 
                           n58680, ZN => n64573);
   U49810 : AOI22_X1 port map( A1 => n67568, A2 => n9033, B1 => n67562, B2 => 
                           n57401, ZN => n64556);
   U49811 : AOI22_X1 port map( A1 => n67592, A2 => n66528, B1 => n58405, B2 => 
                           n67586, ZN => n64554);
   U49812 : AOI22_X1 port map( A1 => n67616, A2 => n57391, B1 => n67610, B2 => 
                           n58681, ZN => n64553);
   U49813 : AOI22_X1 port map( A1 => n67568, A2 => n9031, B1 => n67562, B2 => 
                           n57377, ZN => n64536);
   U49814 : AOI22_X1 port map( A1 => n67592, A2 => n66529, B1 => n58406, B2 => 
                           n67586, ZN => n64534);
   U49815 : AOI22_X1 port map( A1 => n67616, A2 => n57367, B1 => n67610, B2 => 
                           n58682, ZN => n64533);
   U49816 : AOI22_X1 port map( A1 => n67568, A2 => n9029, B1 => n67562, B2 => 
                           n57353, ZN => n64516);
   U49817 : AOI22_X1 port map( A1 => n67592, A2 => n66530, B1 => n58407, B2 => 
                           n67586, ZN => n64514);
   U49818 : AOI22_X1 port map( A1 => n67616, A2 => n57343, B1 => n67610, B2 => 
                           n58683, ZN => n64513);
   U49819 : AOI22_X1 port map( A1 => n67568, A2 => n9027, B1 => n67562, B2 => 
                           n57329, ZN => n64496);
   U49820 : AOI22_X1 port map( A1 => n67592, A2 => n66531, B1 => n58408, B2 => 
                           n67586, ZN => n64494);
   U49821 : AOI22_X1 port map( A1 => n67616, A2 => n57319, B1 => n67610, B2 => 
                           n58684, ZN => n64493);
   U49822 : AOI22_X1 port map( A1 => n67568, A2 => n9025, B1 => n67562, B2 => 
                           n57305, ZN => n64476);
   U49823 : AOI22_X1 port map( A1 => n67592, A2 => n66532, B1 => n58409, B2 => 
                           n67586, ZN => n64474);
   U49824 : AOI22_X1 port map( A1 => n67616, A2 => n57295, B1 => n67610, B2 => 
                           n58685, ZN => n64473);
   U49825 : AOI22_X1 port map( A1 => n67568, A2 => n9023, B1 => n67562, B2 => 
                           n57281, ZN => n64456);
   U49826 : AOI22_X1 port map( A1 => n67592, A2 => n66533, B1 => n58410, B2 => 
                           n67586, ZN => n64454);
   U49827 : AOI22_X1 port map( A1 => n67616, A2 => n57271, B1 => n67610, B2 => 
                           n58686, ZN => n64453);
   U49828 : AOI22_X1 port map( A1 => n67568, A2 => n9021, B1 => n67562, B2 => 
                           n57257, ZN => n64436);
   U49829 : AOI22_X1 port map( A1 => n67592, A2 => n66534, B1 => n58411, B2 => 
                           n67586, ZN => n64434);
   U49830 : AOI22_X1 port map( A1 => n67616, A2 => n57247, B1 => n67610, B2 => 
                           n58687, ZN => n64433);
   U49831 : AOI22_X1 port map( A1 => n67568, A2 => n9019, B1 => n67562, B2 => 
                           n57233, ZN => n64416);
   U49832 : AOI22_X1 port map( A1 => n67592, A2 => n66535, B1 => n58412, B2 => 
                           n67586, ZN => n64414);
   U49833 : AOI22_X1 port map( A1 => n67616, A2 => n57223, B1 => n67610, B2 => 
                           n58688, ZN => n64413);
   U49834 : AOI22_X1 port map( A1 => n67568, A2 => n9017, B1 => n67562, B2 => 
                           n57209, ZN => n64396);
   U49835 : AOI22_X1 port map( A1 => n67592, A2 => n66536, B1 => n58413, B2 => 
                           n67586, ZN => n64394);
   U49836 : AOI22_X1 port map( A1 => n67616, A2 => n57199, B1 => n67610, B2 => 
                           n58689, ZN => n64393);
   U49837 : AOI22_X1 port map( A1 => n67568, A2 => n9015, B1 => n67562, B2 => 
                           n57185, ZN => n64376);
   U49838 : AOI22_X1 port map( A1 => n67592, A2 => n66537, B1 => n58414, B2 => 
                           n67586, ZN => n64374);
   U49839 : AOI22_X1 port map( A1 => n67616, A2 => n57175, B1 => n67610, B2 => 
                           n58690, ZN => n64373);
   U49840 : AOI22_X1 port map( A1 => n67569, A2 => n9013, B1 => n67563, B2 => 
                           n57161, ZN => n64356);
   U49841 : AOI22_X1 port map( A1 => n67593, A2 => n66538, B1 => n58415, B2 => 
                           n67587, ZN => n64354);
   U49842 : AOI22_X1 port map( A1 => n67617, A2 => n57151, B1 => n67611, B2 => 
                           n58691, ZN => n64353);
   U49843 : AOI22_X1 port map( A1 => n67569, A2 => n9011, B1 => n67563, B2 => 
                           n57137, ZN => n64336);
   U49844 : AOI22_X1 port map( A1 => n67593, A2 => n66539, B1 => n58416, B2 => 
                           n67587, ZN => n64334);
   U49845 : AOI22_X1 port map( A1 => n67617, A2 => n57127, B1 => n67611, B2 => 
                           n58692, ZN => n64333);
   U49846 : AOI22_X1 port map( A1 => n67569, A2 => n9009, B1 => n67563, B2 => 
                           n57113, ZN => n64316);
   U49847 : AOI22_X1 port map( A1 => n67593, A2 => n66540, B1 => n58417, B2 => 
                           n67587, ZN => n64314);
   U49848 : AOI22_X1 port map( A1 => n67617, A2 => n57103, B1 => n67611, B2 => 
                           n58693, ZN => n64313);
   U49849 : AOI22_X1 port map( A1 => n67569, A2 => n9007, B1 => n67563, B2 => 
                           n57089, ZN => n64296);
   U49850 : AOI22_X1 port map( A1 => n67593, A2 => n66541, B1 => n58418, B2 => 
                           n67587, ZN => n64294);
   U49851 : AOI22_X1 port map( A1 => n67617, A2 => n57079, B1 => n67611, B2 => 
                           n58694, ZN => n64293);
   U49852 : AOI22_X1 port map( A1 => n67569, A2 => n9005, B1 => n67563, B2 => 
                           n57065, ZN => n64276);
   U49853 : AOI22_X1 port map( A1 => n67593, A2 => n66542, B1 => n58419, B2 => 
                           n67587, ZN => n64274);
   U49854 : AOI22_X1 port map( A1 => n67617, A2 => n57055, B1 => n67611, B2 => 
                           n58695, ZN => n64273);
   U49855 : AOI22_X1 port map( A1 => n67569, A2 => n9003, B1 => n67563, B2 => 
                           n57041, ZN => n64256);
   U49856 : AOI22_X1 port map( A1 => n67593, A2 => n66543, B1 => n58420, B2 => 
                           n67587, ZN => n64254);
   U49857 : AOI22_X1 port map( A1 => n67617, A2 => n57031, B1 => n67611, B2 => 
                           n58696, ZN => n64253);
   U49858 : AOI22_X1 port map( A1 => n67569, A2 => n9001, B1 => n67563, B2 => 
                           n57017, ZN => n64236);
   U49859 : AOI22_X1 port map( A1 => n67593, A2 => n66544, B1 => n58421, B2 => 
                           n67587, ZN => n64234);
   U49860 : AOI22_X1 port map( A1 => n67617, A2 => n57007, B1 => n67611, B2 => 
                           n58697, ZN => n64233);
   U49861 : AOI22_X1 port map( A1 => n67569, A2 => n8999, B1 => n67563, B2 => 
                           n56993, ZN => n64216);
   U49862 : AOI22_X1 port map( A1 => n67593, A2 => n66545, B1 => n58422, B2 => 
                           n67587, ZN => n64214);
   U49863 : AOI22_X1 port map( A1 => n67617, A2 => n56983, B1 => n67611, B2 => 
                           n58698, ZN => n64213);
   U49864 : AOI22_X1 port map( A1 => n67569, A2 => n8997, B1 => n67563, B2 => 
                           n56969, ZN => n64196);
   U49865 : AOI22_X1 port map( A1 => n67593, A2 => n66546, B1 => n58423, B2 => 
                           n67587, ZN => n64194);
   U49866 : AOI22_X1 port map( A1 => n67617, A2 => n56959, B1 => n67611, B2 => 
                           n58699, ZN => n64193);
   U49867 : AOI22_X1 port map( A1 => n67569, A2 => n8995, B1 => n67563, B2 => 
                           n56945, ZN => n64176);
   U49868 : AOI22_X1 port map( A1 => n67593, A2 => n66547, B1 => n58424, B2 => 
                           n67587, ZN => n64174);
   U49869 : AOI22_X1 port map( A1 => n67617, A2 => n56935, B1 => n67611, B2 => 
                           n58700, ZN => n64173);
   U49870 : AOI22_X1 port map( A1 => n67569, A2 => n8993, B1 => n67563, B2 => 
                           n56921, ZN => n64156);
   U49871 : AOI22_X1 port map( A1 => n67593, A2 => n66548, B1 => n58425, B2 => 
                           n67587, ZN => n64154);
   U49872 : AOI22_X1 port map( A1 => n67617, A2 => n56911, B1 => n67611, B2 => 
                           n58701, ZN => n64153);
   U49873 : AOI22_X1 port map( A1 => n67569, A2 => n8991, B1 => n67563, B2 => 
                           n56897, ZN => n64136);
   U49874 : AOI22_X1 port map( A1 => n67593, A2 => n66549, B1 => n58426, B2 => 
                           n67587, ZN => n64134);
   U49875 : AOI22_X1 port map( A1 => n67617, A2 => n56887, B1 => n67611, B2 => 
                           n58702, ZN => n64133);
   U49876 : AOI22_X1 port map( A1 => n67570, A2 => n8989, B1 => n67564, B2 => 
                           n56873, ZN => n64116);
   U49877 : AOI22_X1 port map( A1 => n67618, A2 => n56863, B1 => n67612, B2 => 
                           n58703, ZN => n64113);
   U49878 : AOI22_X1 port map( A1 => n67570, A2 => n8987, B1 => n67564, B2 => 
                           n56849, ZN => n64096);
   U49879 : AOI22_X1 port map( A1 => n67618, A2 => n56839, B1 => n67612, B2 => 
                           n58704, ZN => n64093);
   U49880 : AOI22_X1 port map( A1 => n67570, A2 => n8985, B1 => n67564, B2 => 
                           n56825, ZN => n64076);
   U49881 : AOI22_X1 port map( A1 => n67618, A2 => n56815, B1 => n67612, B2 => 
                           n58705, ZN => n64073);
   U49882 : AOI22_X1 port map( A1 => n67570, A2 => n8983, B1 => n67564, B2 => 
                           n56801, ZN => n64056);
   U49883 : AOI22_X1 port map( A1 => n67618, A2 => n56791, B1 => n67612, B2 => 
                           n58706, ZN => n64053);
   U49884 : AOI22_X1 port map( A1 => n67570, A2 => n8981, B1 => n67564, B2 => 
                           n56777, ZN => n64036);
   U49885 : AOI22_X1 port map( A1 => n67618, A2 => n58643, B1 => n67612, B2 => 
                           n58707, ZN => n64033);
   U49886 : AOI22_X1 port map( A1 => n67570, A2 => n8979, B1 => n67564, B2 => 
                           n56753, ZN => n64016);
   U49887 : AOI22_X1 port map( A1 => n67618, A2 => n58644, B1 => n67612, B2 => 
                           n58708, ZN => n64013);
   U49888 : AOI22_X1 port map( A1 => n67570, A2 => n8977, B1 => n67564, B2 => 
                           n56729, ZN => n63996);
   U49889 : AOI22_X1 port map( A1 => n67618, A2 => n58645, B1 => n67612, B2 => 
                           n58709, ZN => n63993);
   U49890 : AOI22_X1 port map( A1 => n67570, A2 => n8975, B1 => n67564, B2 => 
                           n56705, ZN => n63976);
   U49891 : AOI22_X1 port map( A1 => n67618, A2 => n58646, B1 => n67612, B2 => 
                           n58710, ZN => n63973);
   U49892 : AOI22_X1 port map( A1 => n67570, A2 => n8973, B1 => n67564, B2 => 
                           n56681, ZN => n63956);
   U49893 : AOI22_X1 port map( A1 => n67618, A2 => n58647, B1 => n67612, B2 => 
                           n58711, ZN => n63953);
   U49894 : AOI22_X1 port map( A1 => n67570, A2 => n8971, B1 => n67564, B2 => 
                           n56657, ZN => n63936);
   U49895 : AOI22_X1 port map( A1 => n67618, A2 => n58648, B1 => n67612, B2 => 
                           n58712, ZN => n63933);
   U49896 : AOI22_X1 port map( A1 => n67570, A2 => n8969, B1 => n67564, B2 => 
                           n56633, ZN => n63916);
   U49897 : AOI22_X1 port map( A1 => n67618, A2 => n58649, B1 => n67612, B2 => 
                           n58713, ZN => n63913);
   U49898 : AOI22_X1 port map( A1 => n67570, A2 => n8967, B1 => n67564, B2 => 
                           n56609, ZN => n63896);
   U49899 : AOI22_X1 port map( A1 => n67618, A2 => n58650, B1 => n67612, B2 => 
                           n58714, ZN => n63893);
   U49900 : OAI221_X1 port map( B1 => n63427, B2 => n67452, C1 => n49232, C2 =>
                           n67446, A => n66275, ZN => n66274);
   U49901 : AOI22_X1 port map( A1 => n67440, A2 => n58379, B1 => n67434, B2 => 
                           OUT2_0_port, ZN => n66275);
   U49902 : OAI221_X1 port map( B1 => n63426, B2 => n67452, C1 => n49233, C2 =>
                           n67446, A => n66257, ZN => n66256);
   U49903 : AOI22_X1 port map( A1 => n67440, A2 => n58380, B1 => n67434, B2 => 
                           OUT2_1_port, ZN => n66257);
   U49904 : OAI221_X1 port map( B1 => n63425, B2 => n67452, C1 => n49234, C2 =>
                           n67446, A => n66239, ZN => n66238);
   U49905 : AOI22_X1 port map( A1 => n67440, A2 => n58381, B1 => n67434, B2 => 
                           OUT2_2_port, ZN => n66239);
   U49906 : OAI221_X1 port map( B1 => n63424, B2 => n67452, C1 => n49235, C2 =>
                           n67446, A => n66221, ZN => n66220);
   U49907 : AOI22_X1 port map( A1 => n67440, A2 => n58382, B1 => n67434, B2 => 
                           OUT2_3_port, ZN => n66221);
   U49908 : OAI221_X1 port map( B1 => n63423, B2 => n67452, C1 => n49236, C2 =>
                           n67446, A => n66203, ZN => n66202);
   U49909 : AOI22_X1 port map( A1 => n67440, A2 => n58383, B1 => n67434, B2 => 
                           OUT2_4_port, ZN => n66203);
   U49910 : OAI221_X1 port map( B1 => n63422, B2 => n67452, C1 => n49237, C2 =>
                           n67446, A => n66185, ZN => n66184);
   U49911 : AOI22_X1 port map( A1 => n67440, A2 => n58384, B1 => n67434, B2 => 
                           OUT2_5_port, ZN => n66185);
   U49912 : OAI221_X1 port map( B1 => n63421, B2 => n67452, C1 => n49238, C2 =>
                           n67446, A => n66167, ZN => n66166);
   U49913 : AOI22_X1 port map( A1 => n67440, A2 => n58385, B1 => n67434, B2 => 
                           OUT2_6_port, ZN => n66167);
   U49914 : OAI221_X1 port map( B1 => n63420, B2 => n67452, C1 => n49239, C2 =>
                           n67446, A => n66149, ZN => n66148);
   U49915 : AOI22_X1 port map( A1 => n67440, A2 => n58386, B1 => n67434, B2 => 
                           OUT2_7_port, ZN => n66149);
   U49916 : OAI221_X1 port map( B1 => n63419, B2 => n67452, C1 => n49240, C2 =>
                           n67446, A => n66131, ZN => n66130);
   U49917 : AOI22_X1 port map( A1 => n67440, A2 => n58387, B1 => n67434, B2 => 
                           OUT2_8_port, ZN => n66131);
   U49918 : OAI221_X1 port map( B1 => n63418, B2 => n67452, C1 => n49241, C2 =>
                           n67446, A => n66113, ZN => n66112);
   U49919 : AOI22_X1 port map( A1 => n67440, A2 => n58388, B1 => n67435, B2 => 
                           OUT2_9_port, ZN => n66113);
   U49920 : OAI221_X1 port map( B1 => n63417, B2 => n67452, C1 => n49242, C2 =>
                           n67446, A => n66095, ZN => n66094);
   U49921 : AOI22_X1 port map( A1 => n67440, A2 => n58389, B1 => n67435, B2 => 
                           OUT2_10_port, ZN => n66095);
   U49922 : OAI221_X1 port map( B1 => n63416, B2 => n67452, C1 => n49243, C2 =>
                           n67446, A => n66077, ZN => n66076);
   U49923 : AOI22_X1 port map( A1 => n67440, A2 => n58390, B1 => n67435, B2 => 
                           OUT2_11_port, ZN => n66077);
   U49924 : OAI221_X1 port map( B1 => n63100, B2 => n67631, C1 => n62229, C2 =>
                           n67625, A => n63872, ZN => n63869);
   U49925 : AOI22_X1 port map( A1 => n67619, A2 => n58651, B1 => n67613, B2 => 
                           n58715, ZN => n63872);
   U49926 : OAI221_X1 port map( B1 => n63099, B2 => n67631, C1 => n62228, C2 =>
                           n67625, A => n63851, ZN => n63848);
   U49927 : AOI22_X1 port map( A1 => n67619, A2 => n58652, B1 => n67613, B2 => 
                           n58716, ZN => n63851);
   U49928 : OAI221_X1 port map( B1 => n63098, B2 => n67631, C1 => n62227, C2 =>
                           n67625, A => n63830, ZN => n63827);
   U49929 : AOI22_X1 port map( A1 => n67619, A2 => n58653, B1 => n67613, B2 => 
                           n58717, ZN => n63830);
   U49930 : OAI221_X1 port map( B1 => n62424, B2 => n67607, C1 => n63501, C2 =>
                           n67601, A => n63787, ZN => n63772);
   U49931 : AOI22_X1 port map( A1 => n67595, A2 => n66550, B1 => n67589, B2 => 
                           n58378, ZN => n63787);
   U49932 : OAI221_X1 port map( B1 => n63096, B2 => n67631, C1 => n62225, C2 =>
                           n67625, A => n63782, ZN => n63773);
   U49933 : AOI22_X1 port map( A1 => n67619, A2 => n58654, B1 => n67613, B2 => 
                           n58718, ZN => n63782);
   U49934 : OAI22_X1 port map( A1 => n54670, A2 => n67725, B1 => n68060, B2 => 
                           n67719, ZN => n5759);
   U49935 : OAI22_X1 port map( A1 => n54669, A2 => n67725, B1 => n68063, B2 => 
                           n67719, ZN => n5760);
   U49936 : OAI22_X1 port map( A1 => n54668, A2 => n67725, B1 => n68066, B2 => 
                           n67719, ZN => n5761);
   U49937 : OAI22_X1 port map( A1 => n54667, A2 => n67725, B1 => n68069, B2 => 
                           n67719, ZN => n5762);
   U49938 : OAI22_X1 port map( A1 => n54666, A2 => n67725, B1 => n68072, B2 => 
                           n67719, ZN => n5763);
   U49939 : OAI22_X1 port map( A1 => n54665, A2 => n67725, B1 => n68075, B2 => 
                           n67719, ZN => n5764);
   U49940 : OAI22_X1 port map( A1 => n54664, A2 => n67725, B1 => n68078, B2 => 
                           n67719, ZN => n5765);
   U49941 : OAI22_X1 port map( A1 => n54663, A2 => n67725, B1 => n68081, B2 => 
                           n67719, ZN => n5766);
   U49942 : OAI22_X1 port map( A1 => n54662, A2 => n67725, B1 => n68084, B2 => 
                           n67719, ZN => n5767);
   U49943 : OAI22_X1 port map( A1 => n54661, A2 => n67725, B1 => n68087, B2 => 
                           n67719, ZN => n5768);
   U49944 : OAI22_X1 port map( A1 => n54660, A2 => n67725, B1 => n68090, B2 => 
                           n67719, ZN => n5769);
   U49945 : OAI22_X1 port map( A1 => n54659, A2 => n67726, B1 => n68093, B2 => 
                           n67719, ZN => n5770);
   U49946 : OAI22_X1 port map( A1 => n54658, A2 => n67726, B1 => n68096, B2 => 
                           n67720, ZN => n5771);
   U49947 : OAI22_X1 port map( A1 => n54657, A2 => n67726, B1 => n68099, B2 => 
                           n67720, ZN => n5772);
   U49948 : OAI22_X1 port map( A1 => n54656, A2 => n67726, B1 => n68102, B2 => 
                           n67720, ZN => n5773);
   U49949 : OAI22_X1 port map( A1 => n54655, A2 => n67726, B1 => n68105, B2 => 
                           n67720, ZN => n5774);
   U49950 : OAI22_X1 port map( A1 => n54654, A2 => n67726, B1 => n68108, B2 => 
                           n67720, ZN => n5775);
   U49951 : OAI22_X1 port map( A1 => n54653, A2 => n67726, B1 => n68111, B2 => 
                           n67720, ZN => n5776);
   U49952 : OAI22_X1 port map( A1 => n54652, A2 => n67726, B1 => n68114, B2 => 
                           n67720, ZN => n5777);
   U49953 : OAI22_X1 port map( A1 => n54651, A2 => n67726, B1 => n68117, B2 => 
                           n67720, ZN => n5778);
   U49954 : OAI22_X1 port map( A1 => n54650, A2 => n67726, B1 => n68120, B2 => 
                           n67720, ZN => n5779);
   U49955 : OAI22_X1 port map( A1 => n54649, A2 => n67726, B1 => n68123, B2 => 
                           n67720, ZN => n5780);
   U49956 : OAI22_X1 port map( A1 => n54648, A2 => n67726, B1 => n68126, B2 => 
                           n67720, ZN => n5781);
   U49957 : OAI22_X1 port map( A1 => n54647, A2 => n67727, B1 => n68129, B2 => 
                           n67720, ZN => n5782);
   U49958 : OAI22_X1 port map( A1 => n54646, A2 => n67727, B1 => n68132, B2 => 
                           n67721, ZN => n5783);
   U49959 : OAI22_X1 port map( A1 => n54645, A2 => n67727, B1 => n68135, B2 => 
                           n67721, ZN => n5784);
   U49960 : OAI22_X1 port map( A1 => n54644, A2 => n67727, B1 => n68138, B2 => 
                           n67721, ZN => n5785);
   U49961 : OAI22_X1 port map( A1 => n54643, A2 => n67727, B1 => n68141, B2 => 
                           n67721, ZN => n5786);
   U49962 : OAI22_X1 port map( A1 => n54642, A2 => n67727, B1 => n68144, B2 => 
                           n67721, ZN => n5787);
   U49963 : OAI22_X1 port map( A1 => n54641, A2 => n67727, B1 => n68147, B2 => 
                           n67721, ZN => n5788);
   U49964 : OAI22_X1 port map( A1 => n54640, A2 => n67727, B1 => n68150, B2 => 
                           n67721, ZN => n5789);
   U49965 : OAI22_X1 port map( A1 => n54639, A2 => n67727, B1 => n68153, B2 => 
                           n67721, ZN => n5790);
   U49966 : OAI22_X1 port map( A1 => n54638, A2 => n67727, B1 => n68156, B2 => 
                           n67721, ZN => n5791);
   U49967 : OAI22_X1 port map( A1 => n54637, A2 => n67727, B1 => n68159, B2 => 
                           n67721, ZN => n5792);
   U49968 : OAI22_X1 port map( A1 => n54636, A2 => n67727, B1 => n68162, B2 => 
                           n67721, ZN => n5793);
   U49969 : OAI22_X1 port map( A1 => n54635, A2 => n67728, B1 => n68165, B2 => 
                           n67721, ZN => n5794);
   U49970 : OAI22_X1 port map( A1 => n54634, A2 => n67728, B1 => n68168, B2 => 
                           n67722, ZN => n5795);
   U49971 : OAI22_X1 port map( A1 => n54633, A2 => n67728, B1 => n68171, B2 => 
                           n67722, ZN => n5796);
   U49972 : OAI22_X1 port map( A1 => n54632, A2 => n67728, B1 => n68174, B2 => 
                           n67722, ZN => n5797);
   U49973 : OAI22_X1 port map( A1 => n54631, A2 => n67728, B1 => n68177, B2 => 
                           n67722, ZN => n5798);
   U49974 : OAI22_X1 port map( A1 => n54630, A2 => n67728, B1 => n68180, B2 => 
                           n67722, ZN => n5799);
   U49975 : OAI22_X1 port map( A1 => n54629, A2 => n67728, B1 => n68183, B2 => 
                           n67722, ZN => n5800);
   U49976 : OAI22_X1 port map( A1 => n54628, A2 => n67728, B1 => n68186, B2 => 
                           n67722, ZN => n5801);
   U49977 : OAI22_X1 port map( A1 => n54627, A2 => n67728, B1 => n68189, B2 => 
                           n67722, ZN => n5802);
   U49978 : OAI22_X1 port map( A1 => n54626, A2 => n67728, B1 => n68192, B2 => 
                           n67722, ZN => n5803);
   U49979 : OAI22_X1 port map( A1 => n54625, A2 => n67728, B1 => n68195, B2 => 
                           n67722, ZN => n5804);
   U49980 : OAI22_X1 port map( A1 => n54624, A2 => n67728, B1 => n68198, B2 => 
                           n67722, ZN => n5805);
   U49981 : OAI22_X1 port map( A1 => n54623, A2 => n67729, B1 => n68201, B2 => 
                           n67722, ZN => n5806);
   U49982 : OAI22_X1 port map( A1 => n54622, A2 => n67729, B1 => n68204, B2 => 
                           n67723, ZN => n5807);
   U49983 : OAI22_X1 port map( A1 => n54621, A2 => n67729, B1 => n68207, B2 => 
                           n67723, ZN => n5808);
   U49984 : OAI22_X1 port map( A1 => n54620, A2 => n67729, B1 => n68210, B2 => 
                           n67723, ZN => n5809);
   U49985 : OAI22_X1 port map( A1 => n54619, A2 => n67729, B1 => n68213, B2 => 
                           n67723, ZN => n5810);
   U49986 : OAI22_X1 port map( A1 => n54618, A2 => n67729, B1 => n68216, B2 => 
                           n67723, ZN => n5811);
   U49987 : OAI22_X1 port map( A1 => n54617, A2 => n67729, B1 => n68219, B2 => 
                           n67723, ZN => n5812);
   U49988 : OAI22_X1 port map( A1 => n54616, A2 => n67729, B1 => n68222, B2 => 
                           n67723, ZN => n5813);
   U49989 : OAI22_X1 port map( A1 => n54615, A2 => n67729, B1 => n68225, B2 => 
                           n67723, ZN => n5814);
   U49990 : OAI22_X1 port map( A1 => n54614, A2 => n67729, B1 => n68228, B2 => 
                           n67723, ZN => n5815);
   U49991 : OAI22_X1 port map( A1 => n54613, A2 => n67729, B1 => n68231, B2 => 
                           n67723, ZN => n5816);
   U49992 : OAI22_X1 port map( A1 => n54612, A2 => n67729, B1 => n68234, B2 => 
                           n67723, ZN => n5817);
   U49993 : OAI22_X1 port map( A1 => n54611, A2 => n67730, B1 => n68237, B2 => 
                           n67723, ZN => n5818);
   U49994 : OAI22_X1 port map( A1 => n67662, A2 => n65063, B1 => n68060, B2 => 
                           n67654, ZN => n5376);
   U49995 : OAI22_X1 port map( A1 => n67662, A2 => n65043, B1 => n68063, B2 => 
                           n67654, ZN => n5378);
   U49996 : OAI22_X1 port map( A1 => n67662, A2 => n65023, B1 => n68066, B2 => 
                           n67654, ZN => n5380);
   U49997 : OAI22_X1 port map( A1 => n67662, A2 => n65003, B1 => n68069, B2 => 
                           n67654, ZN => n5382);
   U49998 : OAI22_X1 port map( A1 => n67662, A2 => n64983, B1 => n68072, B2 => 
                           n67654, ZN => n5384);
   U49999 : OAI22_X1 port map( A1 => n67662, A2 => n64963, B1 => n68075, B2 => 
                           n67654, ZN => n5386);
   U50000 : OAI22_X1 port map( A1 => n67662, A2 => n64943, B1 => n68078, B2 => 
                           n67654, ZN => n5388);
   U50001 : OAI22_X1 port map( A1 => n67662, A2 => n64923, B1 => n68081, B2 => 
                           n67654, ZN => n5390);
   U50002 : OAI22_X1 port map( A1 => n67662, A2 => n64903, B1 => n68084, B2 => 
                           n67654, ZN => n5392);
   U50003 : OAI22_X1 port map( A1 => n67662, A2 => n64883, B1 => n68087, B2 => 
                           n67654, ZN => n5394);
   U50004 : OAI22_X1 port map( A1 => n67662, A2 => n64863, B1 => n68090, B2 => 
                           n67654, ZN => n5396);
   U50005 : OAI22_X1 port map( A1 => n67662, A2 => n64843, B1 => n68093, B2 => 
                           n67654, ZN => n5398);
   U50006 : OAI22_X1 port map( A1 => n67663, A2 => n64823, B1 => n68096, B2 => 
                           n67655, ZN => n5400);
   U50007 : OAI22_X1 port map( A1 => n67663, A2 => n64803, B1 => n68099, B2 => 
                           n67655, ZN => n5402);
   U50008 : OAI22_X1 port map( A1 => n67663, A2 => n64783, B1 => n68102, B2 => 
                           n67655, ZN => n5404);
   U50009 : OAI22_X1 port map( A1 => n67663, A2 => n64763, B1 => n68105, B2 => 
                           n67655, ZN => n5406);
   U50010 : OAI22_X1 port map( A1 => n67663, A2 => n64743, B1 => n68108, B2 => 
                           n67655, ZN => n5408);
   U50011 : OAI22_X1 port map( A1 => n67663, A2 => n64723, B1 => n68111, B2 => 
                           n67655, ZN => n5410);
   U50012 : OAI22_X1 port map( A1 => n67663, A2 => n64703, B1 => n68114, B2 => 
                           n67655, ZN => n5412);
   U50013 : OAI22_X1 port map( A1 => n67663, A2 => n64683, B1 => n68117, B2 => 
                           n67655, ZN => n5414);
   U50014 : OAI22_X1 port map( A1 => n67663, A2 => n64663, B1 => n68120, B2 => 
                           n67655, ZN => n5416);
   U50015 : OAI22_X1 port map( A1 => n67663, A2 => n64643, B1 => n68123, B2 => 
                           n67655, ZN => n5418);
   U50016 : OAI22_X1 port map( A1 => n67663, A2 => n64623, B1 => n68126, B2 => 
                           n67655, ZN => n5420);
   U50017 : OAI22_X1 port map( A1 => n67663, A2 => n64603, B1 => n68129, B2 => 
                           n67655, ZN => n5422);
   U50018 : OAI22_X1 port map( A1 => n67663, A2 => n64583, B1 => n68132, B2 => 
                           n67656, ZN => n5424);
   U50019 : OAI22_X1 port map( A1 => n67664, A2 => n64563, B1 => n68135, B2 => 
                           n67656, ZN => n5426);
   U50020 : OAI22_X1 port map( A1 => n67664, A2 => n64543, B1 => n68138, B2 => 
                           n67656, ZN => n5428);
   U50021 : OAI22_X1 port map( A1 => n67664, A2 => n64523, B1 => n68141, B2 => 
                           n67656, ZN => n5430);
   U50022 : OAI22_X1 port map( A1 => n67664, A2 => n64503, B1 => n68144, B2 => 
                           n67656, ZN => n5432);
   U50023 : OAI22_X1 port map( A1 => n67664, A2 => n64483, B1 => n68147, B2 => 
                           n67656, ZN => n5434);
   U50024 : OAI22_X1 port map( A1 => n67664, A2 => n64463, B1 => n68150, B2 => 
                           n67656, ZN => n5436);
   U50025 : OAI22_X1 port map( A1 => n67664, A2 => n64443, B1 => n68153, B2 => 
                           n67656, ZN => n5438);
   U50026 : OAI22_X1 port map( A1 => n67664, A2 => n64423, B1 => n68156, B2 => 
                           n67656, ZN => n5440);
   U50027 : OAI22_X1 port map( A1 => n67664, A2 => n64403, B1 => n68159, B2 => 
                           n67656, ZN => n5442);
   U50028 : OAI22_X1 port map( A1 => n67664, A2 => n64383, B1 => n68162, B2 => 
                           n67656, ZN => n5444);
   U50029 : OAI22_X1 port map( A1 => n67664, A2 => n64363, B1 => n68165, B2 => 
                           n67656, ZN => n5446);
   U50030 : OAI22_X1 port map( A1 => n67664, A2 => n64343, B1 => n68168, B2 => 
                           n67657, ZN => n5448);
   U50031 : OAI22_X1 port map( A1 => n67664, A2 => n64323, B1 => n68171, B2 => 
                           n67657, ZN => n5450);
   U50032 : OAI22_X1 port map( A1 => n67665, A2 => n64303, B1 => n68174, B2 => 
                           n67657, ZN => n5452);
   U50033 : OAI22_X1 port map( A1 => n67665, A2 => n64283, B1 => n68177, B2 => 
                           n67657, ZN => n5454);
   U50034 : OAI22_X1 port map( A1 => n67665, A2 => n64263, B1 => n68180, B2 => 
                           n67657, ZN => n5456);
   U50035 : OAI22_X1 port map( A1 => n67665, A2 => n64243, B1 => n68183, B2 => 
                           n67657, ZN => n5458);
   U50036 : OAI22_X1 port map( A1 => n67665, A2 => n64223, B1 => n68186, B2 => 
                           n67657, ZN => n5460);
   U50037 : OAI22_X1 port map( A1 => n67665, A2 => n64203, B1 => n68189, B2 => 
                           n67657, ZN => n5462);
   U50038 : OAI22_X1 port map( A1 => n67665, A2 => n64183, B1 => n68192, B2 => 
                           n67657, ZN => n5464);
   U50039 : OAI22_X1 port map( A1 => n67665, A2 => n64163, B1 => n68195, B2 => 
                           n67657, ZN => n5466);
   U50040 : OAI22_X1 port map( A1 => n67665, A2 => n64143, B1 => n68198, B2 => 
                           n67657, ZN => n5468);
   U50041 : OAI22_X1 port map( A1 => n67665, A2 => n64123, B1 => n68201, B2 => 
                           n67657, ZN => n5470);
   U50042 : OAI22_X1 port map( A1 => n67665, A2 => n64103, B1 => n68204, B2 => 
                           n67658, ZN => n5472);
   U50043 : OAI22_X1 port map( A1 => n67665, A2 => n64083, B1 => n68207, B2 => 
                           n67658, ZN => n5474);
   U50044 : OAI22_X1 port map( A1 => n67665, A2 => n64063, B1 => n68210, B2 => 
                           n67658, ZN => n5476);
   U50045 : OAI22_X1 port map( A1 => n67666, A2 => n64043, B1 => n68213, B2 => 
                           n67658, ZN => n5478);
   U50046 : OAI22_X1 port map( A1 => n67666, A2 => n64023, B1 => n68216, B2 => 
                           n67658, ZN => n5480);
   U50047 : OAI22_X1 port map( A1 => n67666, A2 => n64003, B1 => n68219, B2 => 
                           n67658, ZN => n5482);
   U50048 : OAI22_X1 port map( A1 => n67666, A2 => n63983, B1 => n68222, B2 => 
                           n67658, ZN => n5484);
   U50049 : OAI22_X1 port map( A1 => n67666, A2 => n63963, B1 => n68225, B2 => 
                           n67658, ZN => n5486);
   U50050 : OAI22_X1 port map( A1 => n67666, A2 => n63943, B1 => n68228, B2 => 
                           n67658, ZN => n5488);
   U50051 : OAI22_X1 port map( A1 => n67666, A2 => n63923, B1 => n68231, B2 => 
                           n67658, ZN => n5490);
   U50052 : OAI22_X1 port map( A1 => n67666, A2 => n63903, B1 => n68234, B2 => 
                           n67658, ZN => n5492);
   U50053 : OAI22_X1 port map( A1 => n67666, A2 => n63883, B1 => n68237, B2 => 
                           n67658, ZN => n5494);
   U50054 : OAI22_X1 port map( A1 => n67675, A2 => n63763, B1 => n68060, B2 => 
                           n67667, ZN => n5503);
   U50055 : OAI22_X1 port map( A1 => n67675, A2 => n63762, B1 => n68063, B2 => 
                           n67667, ZN => n5504);
   U50056 : OAI22_X1 port map( A1 => n67675, A2 => n63761, B1 => n68066, B2 => 
                           n67667, ZN => n5505);
   U50057 : OAI22_X1 port map( A1 => n67675, A2 => n63760, B1 => n68069, B2 => 
                           n67667, ZN => n5506);
   U50058 : OAI22_X1 port map( A1 => n67675, A2 => n63759, B1 => n68072, B2 => 
                           n67667, ZN => n5507);
   U50059 : OAI22_X1 port map( A1 => n67675, A2 => n63758, B1 => n68075, B2 => 
                           n67667, ZN => n5508);
   U50060 : OAI22_X1 port map( A1 => n67675, A2 => n63757, B1 => n68078, B2 => 
                           n67667, ZN => n5509);
   U50061 : OAI22_X1 port map( A1 => n67675, A2 => n63756, B1 => n68081, B2 => 
                           n67667, ZN => n5510);
   U50062 : OAI22_X1 port map( A1 => n67675, A2 => n63755, B1 => n68084, B2 => 
                           n67667, ZN => n5511);
   U50063 : OAI22_X1 port map( A1 => n67675, A2 => n63754, B1 => n68087, B2 => 
                           n67667, ZN => n5512);
   U50064 : OAI22_X1 port map( A1 => n67675, A2 => n63753, B1 => n68090, B2 => 
                           n67667, ZN => n5513);
   U50065 : OAI22_X1 port map( A1 => n67675, A2 => n63752, B1 => n68093, B2 => 
                           n67667, ZN => n5514);
   U50066 : OAI22_X1 port map( A1 => n67676, A2 => n63751, B1 => n68096, B2 => 
                           n67668, ZN => n5515);
   U50067 : OAI22_X1 port map( A1 => n67676, A2 => n63750, B1 => n68099, B2 => 
                           n67668, ZN => n5516);
   U50068 : OAI22_X1 port map( A1 => n67676, A2 => n63749, B1 => n68102, B2 => 
                           n67668, ZN => n5517);
   U50069 : OAI22_X1 port map( A1 => n67676, A2 => n63748, B1 => n68105, B2 => 
                           n67668, ZN => n5518);
   U50070 : OAI22_X1 port map( A1 => n67676, A2 => n63747, B1 => n68108, B2 => 
                           n67668, ZN => n5519);
   U50071 : OAI22_X1 port map( A1 => n67676, A2 => n63746, B1 => n68111, B2 => 
                           n67668, ZN => n5520);
   U50072 : OAI22_X1 port map( A1 => n67676, A2 => n63745, B1 => n68114, B2 => 
                           n67668, ZN => n5521);
   U50073 : OAI22_X1 port map( A1 => n67676, A2 => n63744, B1 => n68117, B2 => 
                           n67668, ZN => n5522);
   U50074 : OAI22_X1 port map( A1 => n67676, A2 => n63743, B1 => n68120, B2 => 
                           n67668, ZN => n5523);
   U50075 : OAI22_X1 port map( A1 => n67676, A2 => n63742, B1 => n68123, B2 => 
                           n67668, ZN => n5524);
   U50076 : OAI22_X1 port map( A1 => n67676, A2 => n63741, B1 => n68126, B2 => 
                           n67668, ZN => n5525);
   U50077 : OAI22_X1 port map( A1 => n67676, A2 => n63740, B1 => n68129, B2 => 
                           n67668, ZN => n5526);
   U50078 : OAI22_X1 port map( A1 => n67676, A2 => n63739, B1 => n68132, B2 => 
                           n67669, ZN => n5527);
   U50079 : OAI22_X1 port map( A1 => n67677, A2 => n63738, B1 => n68135, B2 => 
                           n67669, ZN => n5528);
   U50080 : OAI22_X1 port map( A1 => n67677, A2 => n63737, B1 => n68138, B2 => 
                           n67669, ZN => n5529);
   U50081 : OAI22_X1 port map( A1 => n67677, A2 => n63736, B1 => n68141, B2 => 
                           n67669, ZN => n5530);
   U50082 : OAI22_X1 port map( A1 => n67677, A2 => n63735, B1 => n68144, B2 => 
                           n67669, ZN => n5531);
   U50083 : OAI22_X1 port map( A1 => n67677, A2 => n63734, B1 => n68147, B2 => 
                           n67669, ZN => n5532);
   U50084 : OAI22_X1 port map( A1 => n67677, A2 => n63733, B1 => n68150, B2 => 
                           n67669, ZN => n5533);
   U50085 : OAI22_X1 port map( A1 => n67677, A2 => n63732, B1 => n68153, B2 => 
                           n67669, ZN => n5534);
   U50086 : OAI22_X1 port map( A1 => n67677, A2 => n63731, B1 => n68156, B2 => 
                           n67669, ZN => n5535);
   U50087 : OAI22_X1 port map( A1 => n67677, A2 => n63730, B1 => n68159, B2 => 
                           n67669, ZN => n5536);
   U50088 : OAI22_X1 port map( A1 => n67677, A2 => n63729, B1 => n68162, B2 => 
                           n67669, ZN => n5537);
   U50089 : OAI22_X1 port map( A1 => n67677, A2 => n63728, B1 => n68165, B2 => 
                           n67669, ZN => n5538);
   U50090 : OAI22_X1 port map( A1 => n67677, A2 => n63727, B1 => n68168, B2 => 
                           n67670, ZN => n5539);
   U50091 : OAI22_X1 port map( A1 => n67677, A2 => n63726, B1 => n68171, B2 => 
                           n67670, ZN => n5540);
   U50092 : OAI22_X1 port map( A1 => n67678, A2 => n63725, B1 => n68174, B2 => 
                           n67670, ZN => n5541);
   U50093 : OAI22_X1 port map( A1 => n67678, A2 => n63724, B1 => n68177, B2 => 
                           n67670, ZN => n5542);
   U50094 : OAI22_X1 port map( A1 => n67678, A2 => n63723, B1 => n68180, B2 => 
                           n67670, ZN => n5543);
   U50095 : OAI22_X1 port map( A1 => n67678, A2 => n63722, B1 => n68183, B2 => 
                           n67670, ZN => n5544);
   U50096 : OAI22_X1 port map( A1 => n67678, A2 => n63721, B1 => n68186, B2 => 
                           n67670, ZN => n5545);
   U50097 : OAI22_X1 port map( A1 => n67678, A2 => n63720, B1 => n68189, B2 => 
                           n67670, ZN => n5546);
   U50098 : OAI22_X1 port map( A1 => n67678, A2 => n63719, B1 => n68192, B2 => 
                           n67670, ZN => n5547);
   U50099 : OAI22_X1 port map( A1 => n67678, A2 => n63718, B1 => n68195, B2 => 
                           n67670, ZN => n5548);
   U50100 : OAI22_X1 port map( A1 => n67678, A2 => n63717, B1 => n68198, B2 => 
                           n67670, ZN => n5549);
   U50101 : OAI22_X1 port map( A1 => n67678, A2 => n63716, B1 => n68201, B2 => 
                           n67670, ZN => n5550);
   U50102 : OAI22_X1 port map( A1 => n67678, A2 => n63715, B1 => n68204, B2 => 
                           n67671, ZN => n5551);
   U50103 : OAI22_X1 port map( A1 => n67678, A2 => n63714, B1 => n68207, B2 => 
                           n67671, ZN => n5552);
   U50104 : OAI22_X1 port map( A1 => n67678, A2 => n63713, B1 => n68210, B2 => 
                           n67671, ZN => n5553);
   U50105 : OAI22_X1 port map( A1 => n67679, A2 => n63712, B1 => n68213, B2 => 
                           n67671, ZN => n5554);
   U50106 : OAI22_X1 port map( A1 => n67679, A2 => n63711, B1 => n68216, B2 => 
                           n67671, ZN => n5555);
   U50107 : OAI22_X1 port map( A1 => n67679, A2 => n63710, B1 => n68219, B2 => 
                           n67671, ZN => n5556);
   U50108 : OAI22_X1 port map( A1 => n67679, A2 => n63709, B1 => n68222, B2 => 
                           n67671, ZN => n5557);
   U50109 : OAI22_X1 port map( A1 => n67679, A2 => n63708, B1 => n68225, B2 => 
                           n67671, ZN => n5558);
   U50110 : OAI22_X1 port map( A1 => n67679, A2 => n63707, B1 => n68228, B2 => 
                           n67671, ZN => n5559);
   U50111 : OAI22_X1 port map( A1 => n67679, A2 => n63706, B1 => n68231, B2 => 
                           n67671, ZN => n5560);
   U50112 : OAI22_X1 port map( A1 => n67679, A2 => n63705, B1 => n68234, B2 => 
                           n67671, ZN => n5561);
   U50113 : OAI22_X1 port map( A1 => n67679, A2 => n63704, B1 => n68237, B2 => 
                           n67671, ZN => n5562);
   U50114 : OAI22_X1 port map( A1 => n54246, A2 => n67929, B1 => n68058, B2 => 
                           n67923, ZN => n6783);
   U50115 : OAI22_X1 port map( A1 => n54245, A2 => n67929, B1 => n68061, B2 => 
                           n67923, ZN => n6784);
   U50116 : OAI22_X1 port map( A1 => n54244, A2 => n67929, B1 => n68064, B2 => 
                           n67923, ZN => n6785);
   U50117 : OAI22_X1 port map( A1 => n54243, A2 => n67929, B1 => n68067, B2 => 
                           n67923, ZN => n6786);
   U50118 : OAI22_X1 port map( A1 => n54242, A2 => n67929, B1 => n68070, B2 => 
                           n67923, ZN => n6787);
   U50119 : OAI22_X1 port map( A1 => n54241, A2 => n67929, B1 => n68073, B2 => 
                           n67923, ZN => n6788);
   U50120 : OAI22_X1 port map( A1 => n54240, A2 => n67929, B1 => n68076, B2 => 
                           n67923, ZN => n6789);
   U50121 : OAI22_X1 port map( A1 => n54239, A2 => n67929, B1 => n68079, B2 => 
                           n67923, ZN => n6790);
   U50122 : OAI22_X1 port map( A1 => n54238, A2 => n67929, B1 => n68082, B2 => 
                           n67923, ZN => n6791);
   U50123 : OAI22_X1 port map( A1 => n54237, A2 => n67929, B1 => n68085, B2 => 
                           n67923, ZN => n6792);
   U50124 : OAI22_X1 port map( A1 => n54236, A2 => n67929, B1 => n68088, B2 => 
                           n67923, ZN => n6793);
   U50125 : OAI22_X1 port map( A1 => n54235, A2 => n67930, B1 => n68091, B2 => 
                           n67923, ZN => n6794);
   U50126 : OAI22_X1 port map( A1 => n54234, A2 => n67930, B1 => n68094, B2 => 
                           n67924, ZN => n6795);
   U50127 : OAI22_X1 port map( A1 => n54233, A2 => n67930, B1 => n68097, B2 => 
                           n67924, ZN => n6796);
   U50128 : OAI22_X1 port map( A1 => n54232, A2 => n67930, B1 => n68100, B2 => 
                           n67924, ZN => n6797);
   U50129 : OAI22_X1 port map( A1 => n54231, A2 => n67930, B1 => n68103, B2 => 
                           n67924, ZN => n6798);
   U50130 : OAI22_X1 port map( A1 => n54230, A2 => n67930, B1 => n68106, B2 => 
                           n67924, ZN => n6799);
   U50131 : OAI22_X1 port map( A1 => n54229, A2 => n67930, B1 => n68109, B2 => 
                           n67924, ZN => n6800);
   U50132 : OAI22_X1 port map( A1 => n54228, A2 => n67930, B1 => n68112, B2 => 
                           n67924, ZN => n6801);
   U50133 : OAI22_X1 port map( A1 => n54227, A2 => n67930, B1 => n68115, B2 => 
                           n67924, ZN => n6802);
   U50134 : OAI22_X1 port map( A1 => n54226, A2 => n67930, B1 => n68118, B2 => 
                           n67924, ZN => n6803);
   U50135 : OAI22_X1 port map( A1 => n54225, A2 => n67930, B1 => n68121, B2 => 
                           n67924, ZN => n6804);
   U50136 : OAI22_X1 port map( A1 => n54224, A2 => n67930, B1 => n68124, B2 => 
                           n67924, ZN => n6805);
   U50137 : OAI22_X1 port map( A1 => n54223, A2 => n67931, B1 => n68127, B2 => 
                           n67924, ZN => n6806);
   U50138 : OAI22_X1 port map( A1 => n54222, A2 => n67931, B1 => n68130, B2 => 
                           n67925, ZN => n6807);
   U50139 : OAI22_X1 port map( A1 => n54221, A2 => n67931, B1 => n68133, B2 => 
                           n67925, ZN => n6808);
   U50140 : OAI22_X1 port map( A1 => n54220, A2 => n67931, B1 => n68136, B2 => 
                           n67925, ZN => n6809);
   U50141 : OAI22_X1 port map( A1 => n54219, A2 => n67931, B1 => n68139, B2 => 
                           n67925, ZN => n6810);
   U50142 : OAI22_X1 port map( A1 => n54218, A2 => n67931, B1 => n68142, B2 => 
                           n67925, ZN => n6811);
   U50143 : OAI22_X1 port map( A1 => n54217, A2 => n67931, B1 => n68145, B2 => 
                           n67925, ZN => n6812);
   U50144 : OAI22_X1 port map( A1 => n54216, A2 => n67931, B1 => n68148, B2 => 
                           n67925, ZN => n6813);
   U50145 : OAI22_X1 port map( A1 => n54215, A2 => n67931, B1 => n68151, B2 => 
                           n67925, ZN => n6814);
   U50146 : OAI22_X1 port map( A1 => n54214, A2 => n67931, B1 => n68154, B2 => 
                           n67925, ZN => n6815);
   U50147 : OAI22_X1 port map( A1 => n54213, A2 => n67931, B1 => n68157, B2 => 
                           n67925, ZN => n6816);
   U50148 : OAI22_X1 port map( A1 => n54212, A2 => n67931, B1 => n68160, B2 => 
                           n67925, ZN => n6817);
   U50149 : OAI22_X1 port map( A1 => n54211, A2 => n67932, B1 => n68163, B2 => 
                           n67925, ZN => n6818);
   U50150 : OAI22_X1 port map( A1 => n54210, A2 => n67932, B1 => n68166, B2 => 
                           n67926, ZN => n6819);
   U50151 : OAI22_X1 port map( A1 => n54209, A2 => n67932, B1 => n68169, B2 => 
                           n67926, ZN => n6820);
   U50152 : OAI22_X1 port map( A1 => n54208, A2 => n67932, B1 => n68172, B2 => 
                           n67926, ZN => n6821);
   U50153 : OAI22_X1 port map( A1 => n54207, A2 => n67932, B1 => n68175, B2 => 
                           n67926, ZN => n6822);
   U50154 : OAI22_X1 port map( A1 => n54206, A2 => n67932, B1 => n68178, B2 => 
                           n67926, ZN => n6823);
   U50155 : OAI22_X1 port map( A1 => n54205, A2 => n67932, B1 => n68181, B2 => 
                           n67926, ZN => n6824);
   U50156 : OAI22_X1 port map( A1 => n54204, A2 => n67932, B1 => n68184, B2 => 
                           n67926, ZN => n6825);
   U50157 : OAI22_X1 port map( A1 => n54203, A2 => n67932, B1 => n68187, B2 => 
                           n67926, ZN => n6826);
   U50158 : OAI22_X1 port map( A1 => n54202, A2 => n67932, B1 => n68190, B2 => 
                           n67926, ZN => n6827);
   U50159 : OAI22_X1 port map( A1 => n54201, A2 => n67932, B1 => n68193, B2 => 
                           n67926, ZN => n6828);
   U50160 : OAI22_X1 port map( A1 => n54200, A2 => n67932, B1 => n68196, B2 => 
                           n67926, ZN => n6829);
   U50161 : OAI22_X1 port map( A1 => n54199, A2 => n67933, B1 => n68199, B2 => 
                           n67926, ZN => n6830);
   U50162 : OAI22_X1 port map( A1 => n54198, A2 => n67933, B1 => n68202, B2 => 
                           n67927, ZN => n6831);
   U50163 : OAI22_X1 port map( A1 => n54197, A2 => n67933, B1 => n68205, B2 => 
                           n67927, ZN => n6832);
   U50164 : OAI22_X1 port map( A1 => n54196, A2 => n67933, B1 => n68208, B2 => 
                           n67927, ZN => n6833);
   U50165 : OAI22_X1 port map( A1 => n54195, A2 => n67933, B1 => n68211, B2 => 
                           n67927, ZN => n6834);
   U50166 : OAI22_X1 port map( A1 => n54194, A2 => n67933, B1 => n68214, B2 => 
                           n67927, ZN => n6835);
   U50167 : OAI22_X1 port map( A1 => n54193, A2 => n67933, B1 => n68217, B2 => 
                           n67927, ZN => n6836);
   U50168 : OAI22_X1 port map( A1 => n54192, A2 => n67933, B1 => n68220, B2 => 
                           n67927, ZN => n6837);
   U50169 : OAI22_X1 port map( A1 => n54191, A2 => n67933, B1 => n68223, B2 => 
                           n67927, ZN => n6838);
   U50170 : OAI22_X1 port map( A1 => n54190, A2 => n67933, B1 => n68226, B2 => 
                           n67927, ZN => n6839);
   U50171 : OAI22_X1 port map( A1 => n54189, A2 => n67933, B1 => n68229, B2 => 
                           n67927, ZN => n6840);
   U50172 : OAI22_X1 port map( A1 => n54188, A2 => n67933, B1 => n68232, B2 => 
                           n67927, ZN => n6841);
   U50173 : OAI22_X1 port map( A1 => n54187, A2 => n67934, B1 => n68235, B2 => 
                           n67927, ZN => n6842);
   U50174 : OAI22_X1 port map( A1 => n49232, A2 => n67904, B1 => n68059, B2 => 
                           n67898, ZN => n6655);
   U50175 : OAI22_X1 port map( A1 => n49233, A2 => n67904, B1 => n68062, B2 => 
                           n67898, ZN => n6656);
   U50176 : OAI22_X1 port map( A1 => n49234, A2 => n67904, B1 => n68065, B2 => 
                           n67898, ZN => n6657);
   U50177 : OAI22_X1 port map( A1 => n49235, A2 => n67904, B1 => n68068, B2 => 
                           n67898, ZN => n6658);
   U50178 : OAI22_X1 port map( A1 => n49236, A2 => n67904, B1 => n68071, B2 => 
                           n67898, ZN => n6659);
   U50179 : OAI22_X1 port map( A1 => n49237, A2 => n67904, B1 => n68074, B2 => 
                           n67898, ZN => n6660);
   U50180 : OAI22_X1 port map( A1 => n49238, A2 => n67904, B1 => n68077, B2 => 
                           n67898, ZN => n6661);
   U50181 : OAI22_X1 port map( A1 => n49239, A2 => n67904, B1 => n68080, B2 => 
                           n67898, ZN => n6662);
   U50182 : OAI22_X1 port map( A1 => n49240, A2 => n67904, B1 => n68083, B2 => 
                           n67898, ZN => n6663);
   U50183 : OAI22_X1 port map( A1 => n49241, A2 => n67904, B1 => n68086, B2 => 
                           n67898, ZN => n6664);
   U50184 : OAI22_X1 port map( A1 => n49242, A2 => n67904, B1 => n68089, B2 => 
                           n67898, ZN => n6665);
   U50185 : OAI22_X1 port map( A1 => n49243, A2 => n67905, B1 => n68092, B2 => 
                           n67898, ZN => n6666);
   U50186 : OAI22_X1 port map( A1 => n49244, A2 => n67905, B1 => n68095, B2 => 
                           n67899, ZN => n6667);
   U50187 : OAI22_X1 port map( A1 => n49245, A2 => n67905, B1 => n68098, B2 => 
                           n67899, ZN => n6668);
   U50188 : OAI22_X1 port map( A1 => n49246, A2 => n67905, B1 => n68101, B2 => 
                           n67899, ZN => n6669);
   U50189 : OAI22_X1 port map( A1 => n49247, A2 => n67905, B1 => n68104, B2 => 
                           n67899, ZN => n6670);
   U50190 : OAI22_X1 port map( A1 => n49248, A2 => n67905, B1 => n68107, B2 => 
                           n67899, ZN => n6671);
   U50191 : OAI22_X1 port map( A1 => n49249, A2 => n67905, B1 => n68110, B2 => 
                           n67899, ZN => n6672);
   U50192 : OAI22_X1 port map( A1 => n49250, A2 => n67905, B1 => n68113, B2 => 
                           n67899, ZN => n6673);
   U50193 : OAI22_X1 port map( A1 => n49251, A2 => n67905, B1 => n68116, B2 => 
                           n67899, ZN => n6674);
   U50194 : OAI22_X1 port map( A1 => n49252, A2 => n67905, B1 => n68119, B2 => 
                           n67899, ZN => n6675);
   U50195 : OAI22_X1 port map( A1 => n49253, A2 => n67905, B1 => n68122, B2 => 
                           n67899, ZN => n6676);
   U50196 : OAI22_X1 port map( A1 => n49254, A2 => n67905, B1 => n68125, B2 => 
                           n67899, ZN => n6677);
   U50197 : OAI22_X1 port map( A1 => n49255, A2 => n67906, B1 => n68128, B2 => 
                           n67899, ZN => n6678);
   U50198 : OAI22_X1 port map( A1 => n49256, A2 => n67906, B1 => n68131, B2 => 
                           n67900, ZN => n6679);
   U50199 : OAI22_X1 port map( A1 => n49257, A2 => n67906, B1 => n68134, B2 => 
                           n67900, ZN => n6680);
   U50200 : OAI22_X1 port map( A1 => n49258, A2 => n67906, B1 => n68137, B2 => 
                           n67900, ZN => n6681);
   U50201 : OAI22_X1 port map( A1 => n49259, A2 => n67906, B1 => n68140, B2 => 
                           n67900, ZN => n6682);
   U50202 : OAI22_X1 port map( A1 => n49260, A2 => n67906, B1 => n68143, B2 => 
                           n67900, ZN => n6683);
   U50203 : OAI22_X1 port map( A1 => n49261, A2 => n67906, B1 => n68146, B2 => 
                           n67900, ZN => n6684);
   U50204 : OAI22_X1 port map( A1 => n49262, A2 => n67906, B1 => n68149, B2 => 
                           n67900, ZN => n6685);
   U50205 : OAI22_X1 port map( A1 => n49263, A2 => n67906, B1 => n68152, B2 => 
                           n67900, ZN => n6686);
   U50206 : OAI22_X1 port map( A1 => n49264, A2 => n67906, B1 => n68155, B2 => 
                           n67900, ZN => n6687);
   U50207 : OAI22_X1 port map( A1 => n49265, A2 => n67906, B1 => n68158, B2 => 
                           n67900, ZN => n6688);
   U50208 : OAI22_X1 port map( A1 => n49266, A2 => n67906, B1 => n68161, B2 => 
                           n67900, ZN => n6689);
   U50209 : OAI22_X1 port map( A1 => n49267, A2 => n67907, B1 => n68164, B2 => 
                           n67900, ZN => n6690);
   U50210 : OAI22_X1 port map( A1 => n49268, A2 => n67907, B1 => n68167, B2 => 
                           n67901, ZN => n6691);
   U50211 : OAI22_X1 port map( A1 => n49269, A2 => n67907, B1 => n68170, B2 => 
                           n67901, ZN => n6692);
   U50212 : OAI22_X1 port map( A1 => n49270, A2 => n67907, B1 => n68173, B2 => 
                           n67901, ZN => n6693);
   U50213 : OAI22_X1 port map( A1 => n49271, A2 => n67907, B1 => n68176, B2 => 
                           n67901, ZN => n6694);
   U50214 : OAI22_X1 port map( A1 => n49272, A2 => n67907, B1 => n68179, B2 => 
                           n67901, ZN => n6695);
   U50215 : OAI22_X1 port map( A1 => n49273, A2 => n67907, B1 => n68182, B2 => 
                           n67901, ZN => n6696);
   U50216 : OAI22_X1 port map( A1 => n49274, A2 => n67907, B1 => n68185, B2 => 
                           n67901, ZN => n6697);
   U50217 : OAI22_X1 port map( A1 => n49275, A2 => n67907, B1 => n68188, B2 => 
                           n67901, ZN => n6698);
   U50218 : OAI22_X1 port map( A1 => n49276, A2 => n67907, B1 => n68191, B2 => 
                           n67901, ZN => n6699);
   U50219 : OAI22_X1 port map( A1 => n49277, A2 => n67907, B1 => n68194, B2 => 
                           n67901, ZN => n6700);
   U50220 : OAI22_X1 port map( A1 => n49278, A2 => n67907, B1 => n68197, B2 => 
                           n67901, ZN => n6701);
   U50221 : OAI22_X1 port map( A1 => n49279, A2 => n67908, B1 => n68200, B2 => 
                           n67901, ZN => n6702);
   U50222 : OAI22_X1 port map( A1 => n49280, A2 => n67908, B1 => n68203, B2 => 
                           n67902, ZN => n6703);
   U50223 : OAI22_X1 port map( A1 => n49281, A2 => n67908, B1 => n68206, B2 => 
                           n67902, ZN => n6704);
   U50224 : OAI22_X1 port map( A1 => n49282, A2 => n67908, B1 => n68209, B2 => 
                           n67902, ZN => n6705);
   U50225 : OAI22_X1 port map( A1 => n49283, A2 => n67908, B1 => n68212, B2 => 
                           n67902, ZN => n6706);
   U50226 : OAI22_X1 port map( A1 => n49284, A2 => n67908, B1 => n68215, B2 => 
                           n67902, ZN => n6707);
   U50227 : OAI22_X1 port map( A1 => n49285, A2 => n67908, B1 => n68218, B2 => 
                           n67902, ZN => n6708);
   U50228 : OAI22_X1 port map( A1 => n49286, A2 => n67908, B1 => n68221, B2 => 
                           n67902, ZN => n6709);
   U50229 : OAI22_X1 port map( A1 => n49287, A2 => n67908, B1 => n68224, B2 => 
                           n67902, ZN => n6710);
   U50230 : OAI22_X1 port map( A1 => n49288, A2 => n67908, B1 => n68227, B2 => 
                           n67902, ZN => n6711);
   U50231 : OAI22_X1 port map( A1 => n49289, A2 => n67908, B1 => n68230, B2 => 
                           n67902, ZN => n6712);
   U50232 : OAI22_X1 port map( A1 => n49290, A2 => n67908, B1 => n68233, B2 => 
                           n67902, ZN => n6713);
   U50233 : OAI22_X1 port map( A1 => n49291, A2 => n67909, B1 => n68236, B2 => 
                           n67902, ZN => n6714);
   U50234 : OAI22_X1 port map( A1 => n68258, A2 => n62085, B1 => n68250, B2 => 
                           n68058, ZN => n7423);
   U50235 : OAI22_X1 port map( A1 => n68258, A2 => n62083, B1 => n68250, B2 => 
                           n68061, ZN => n7424);
   U50236 : OAI22_X1 port map( A1 => n68258, A2 => n62081, B1 => n68250, B2 => 
                           n68064, ZN => n7425);
   U50237 : OAI22_X1 port map( A1 => n68258, A2 => n62079, B1 => n68250, B2 => 
                           n68067, ZN => n7426);
   U50238 : OAI22_X1 port map( A1 => n68258, A2 => n62077, B1 => n68250, B2 => 
                           n68070, ZN => n7427);
   U50239 : OAI22_X1 port map( A1 => n68258, A2 => n62075, B1 => n68250, B2 => 
                           n68073, ZN => n7428);
   U50240 : OAI22_X1 port map( A1 => n68258, A2 => n62073, B1 => n68250, B2 => 
                           n68076, ZN => n7429);
   U50241 : OAI22_X1 port map( A1 => n68258, A2 => n62071, B1 => n68250, B2 => 
                           n68079, ZN => n7430);
   U50242 : OAI22_X1 port map( A1 => n68258, A2 => n62069, B1 => n68250, B2 => 
                           n68082, ZN => n7431);
   U50243 : OAI22_X1 port map( A1 => n68258, A2 => n62067, B1 => n68250, B2 => 
                           n68085, ZN => n7432);
   U50244 : OAI22_X1 port map( A1 => n68258, A2 => n62065, B1 => n68250, B2 => 
                           n68088, ZN => n7433);
   U50245 : OAI22_X1 port map( A1 => n68258, A2 => n62063, B1 => n68250, B2 => 
                           n68091, ZN => n7434);
   U50246 : OAI22_X1 port map( A1 => n49420, A2 => n67827, B1 => n68059, B2 => 
                           n67821, ZN => n6271);
   U50247 : OAI22_X1 port map( A1 => n49421, A2 => n67827, B1 => n68062, B2 => 
                           n67821, ZN => n6272);
   U50248 : OAI22_X1 port map( A1 => n49422, A2 => n67827, B1 => n68065, B2 => 
                           n67821, ZN => n6273);
   U50249 : OAI22_X1 port map( A1 => n49423, A2 => n67827, B1 => n68068, B2 => 
                           n67821, ZN => n6274);
   U50250 : OAI22_X1 port map( A1 => n49424, A2 => n67827, B1 => n68071, B2 => 
                           n67821, ZN => n6275);
   U50251 : OAI22_X1 port map( A1 => n49425, A2 => n67827, B1 => n68074, B2 => 
                           n67821, ZN => n6276);
   U50252 : OAI22_X1 port map( A1 => n49426, A2 => n67827, B1 => n68077, B2 => 
                           n67821, ZN => n6277);
   U50253 : OAI22_X1 port map( A1 => n49427, A2 => n67827, B1 => n68080, B2 => 
                           n67821, ZN => n6278);
   U50254 : OAI22_X1 port map( A1 => n49428, A2 => n67827, B1 => n68083, B2 => 
                           n67821, ZN => n6279);
   U50255 : OAI22_X1 port map( A1 => n49429, A2 => n67827, B1 => n68086, B2 => 
                           n67821, ZN => n6280);
   U50256 : OAI22_X1 port map( A1 => n49430, A2 => n67827, B1 => n68089, B2 => 
                           n67821, ZN => n6281);
   U50257 : OAI22_X1 port map( A1 => n49431, A2 => n67828, B1 => n68092, B2 => 
                           n67821, ZN => n6282);
   U50258 : OAI22_X1 port map( A1 => n49432, A2 => n67828, B1 => n68095, B2 => 
                           n67822, ZN => n6283);
   U50259 : OAI22_X1 port map( A1 => n49433, A2 => n67828, B1 => n68098, B2 => 
                           n67822, ZN => n6284);
   U50260 : OAI22_X1 port map( A1 => n49434, A2 => n67828, B1 => n68101, B2 => 
                           n67822, ZN => n6285);
   U50261 : OAI22_X1 port map( A1 => n49435, A2 => n67828, B1 => n68104, B2 => 
                           n67822, ZN => n6286);
   U50262 : OAI22_X1 port map( A1 => n49436, A2 => n67828, B1 => n68107, B2 => 
                           n67822, ZN => n6287);
   U50263 : OAI22_X1 port map( A1 => n49437, A2 => n67828, B1 => n68110, B2 => 
                           n67822, ZN => n6288);
   U50264 : OAI22_X1 port map( A1 => n49438, A2 => n67828, B1 => n68113, B2 => 
                           n67822, ZN => n6289);
   U50265 : OAI22_X1 port map( A1 => n49439, A2 => n67828, B1 => n68116, B2 => 
                           n67822, ZN => n6290);
   U50266 : OAI22_X1 port map( A1 => n49440, A2 => n67828, B1 => n68119, B2 => 
                           n67822, ZN => n6291);
   U50267 : OAI22_X1 port map( A1 => n49441, A2 => n67828, B1 => n68122, B2 => 
                           n67822, ZN => n6292);
   U50268 : OAI22_X1 port map( A1 => n49442, A2 => n67828, B1 => n68125, B2 => 
                           n67822, ZN => n6293);
   U50269 : OAI22_X1 port map( A1 => n49443, A2 => n67829, B1 => n68128, B2 => 
                           n67822, ZN => n6294);
   U50270 : OAI22_X1 port map( A1 => n49444, A2 => n67829, B1 => n68131, B2 => 
                           n67823, ZN => n6295);
   U50271 : OAI22_X1 port map( A1 => n49445, A2 => n67829, B1 => n68134, B2 => 
                           n67823, ZN => n6296);
   U50272 : OAI22_X1 port map( A1 => n49446, A2 => n67829, B1 => n68137, B2 => 
                           n67823, ZN => n6297);
   U50273 : OAI22_X1 port map( A1 => n49447, A2 => n67829, B1 => n68140, B2 => 
                           n67823, ZN => n6298);
   U50274 : OAI22_X1 port map( A1 => n49448, A2 => n67829, B1 => n68143, B2 => 
                           n67823, ZN => n6299);
   U50275 : OAI22_X1 port map( A1 => n49449, A2 => n67829, B1 => n68146, B2 => 
                           n67823, ZN => n6300);
   U50276 : OAI22_X1 port map( A1 => n49450, A2 => n67829, B1 => n68149, B2 => 
                           n67823, ZN => n6301);
   U50277 : OAI22_X1 port map( A1 => n49451, A2 => n67829, B1 => n68152, B2 => 
                           n67823, ZN => n6302);
   U50278 : OAI22_X1 port map( A1 => n49452, A2 => n67829, B1 => n68155, B2 => 
                           n67823, ZN => n6303);
   U50279 : OAI22_X1 port map( A1 => n49453, A2 => n67829, B1 => n68158, B2 => 
                           n67823, ZN => n6304);
   U50280 : OAI22_X1 port map( A1 => n49454, A2 => n67829, B1 => n68161, B2 => 
                           n67823, ZN => n6305);
   U50281 : OAI22_X1 port map( A1 => n49455, A2 => n67830, B1 => n68164, B2 => 
                           n67823, ZN => n6306);
   U50282 : OAI22_X1 port map( A1 => n49456, A2 => n67830, B1 => n68167, B2 => 
                           n67824, ZN => n6307);
   U50283 : OAI22_X1 port map( A1 => n49457, A2 => n67830, B1 => n68170, B2 => 
                           n67824, ZN => n6308);
   U50284 : OAI22_X1 port map( A1 => n49458, A2 => n67830, B1 => n68173, B2 => 
                           n67824, ZN => n6309);
   U50285 : OAI22_X1 port map( A1 => n49459, A2 => n67830, B1 => n68176, B2 => 
                           n67824, ZN => n6310);
   U50286 : OAI22_X1 port map( A1 => n49460, A2 => n67830, B1 => n68179, B2 => 
                           n67824, ZN => n6311);
   U50287 : OAI22_X1 port map( A1 => n49461, A2 => n67830, B1 => n68182, B2 => 
                           n67824, ZN => n6312);
   U50288 : OAI22_X1 port map( A1 => n49462, A2 => n67830, B1 => n68185, B2 => 
                           n67824, ZN => n6313);
   U50289 : OAI22_X1 port map( A1 => n49463, A2 => n67830, B1 => n68188, B2 => 
                           n67824, ZN => n6314);
   U50290 : OAI22_X1 port map( A1 => n49464, A2 => n67830, B1 => n68191, B2 => 
                           n67824, ZN => n6315);
   U50291 : OAI22_X1 port map( A1 => n49465, A2 => n67830, B1 => n68194, B2 => 
                           n67824, ZN => n6316);
   U50292 : OAI22_X1 port map( A1 => n49466, A2 => n67830, B1 => n68197, B2 => 
                           n67824, ZN => n6317);
   U50293 : OAI22_X1 port map( A1 => n49467, A2 => n67831, B1 => n68200, B2 => 
                           n67824, ZN => n6318);
   U50294 : OAI22_X1 port map( A1 => n49468, A2 => n67831, B1 => n68203, B2 => 
                           n67825, ZN => n6319);
   U50295 : OAI22_X1 port map( A1 => n49469, A2 => n67831, B1 => n68206, B2 => 
                           n67825, ZN => n6320);
   U50296 : OAI22_X1 port map( A1 => n49470, A2 => n67831, B1 => n68209, B2 => 
                           n67825, ZN => n6321);
   U50297 : OAI22_X1 port map( A1 => n49471, A2 => n67831, B1 => n68212, B2 => 
                           n67825, ZN => n6322);
   U50298 : OAI22_X1 port map( A1 => n49472, A2 => n67831, B1 => n68215, B2 => 
                           n67825, ZN => n6323);
   U50299 : OAI22_X1 port map( A1 => n49473, A2 => n67831, B1 => n68218, B2 => 
                           n67825, ZN => n6324);
   U50300 : OAI22_X1 port map( A1 => n49474, A2 => n67831, B1 => n68221, B2 => 
                           n67825, ZN => n6325);
   U50301 : OAI22_X1 port map( A1 => n49475, A2 => n67831, B1 => n68224, B2 => 
                           n67825, ZN => n6326);
   U50302 : OAI22_X1 port map( A1 => n49476, A2 => n67831, B1 => n68227, B2 => 
                           n67825, ZN => n6327);
   U50303 : OAI22_X1 port map( A1 => n49477, A2 => n67831, B1 => n68230, B2 => 
                           n67825, ZN => n6328);
   U50304 : OAI22_X1 port map( A1 => n49478, A2 => n67831, B1 => n68233, B2 => 
                           n67825, ZN => n6329);
   U50305 : OAI22_X1 port map( A1 => n49479, A2 => n67832, B1 => n68236, B2 => 
                           n67825, ZN => n6330);
   U50306 : OAI22_X1 port map( A1 => n67778, A2 => n63294, B1 => n68059, B2 => 
                           n67770, ZN => n6015);
   U50307 : OAI22_X1 port map( A1 => n67778, A2 => n63293, B1 => n68062, B2 => 
                           n67770, ZN => n6016);
   U50308 : OAI22_X1 port map( A1 => n67778, A2 => n63292, B1 => n68065, B2 => 
                           n67770, ZN => n6017);
   U50309 : OAI22_X1 port map( A1 => n67778, A2 => n63291, B1 => n68068, B2 => 
                           n67770, ZN => n6018);
   U50310 : OAI22_X1 port map( A1 => n67778, A2 => n63290, B1 => n68071, B2 => 
                           n67770, ZN => n6019);
   U50311 : OAI22_X1 port map( A1 => n67778, A2 => n63289, B1 => n68074, B2 => 
                           n67770, ZN => n6020);
   U50312 : OAI22_X1 port map( A1 => n67778, A2 => n63288, B1 => n68077, B2 => 
                           n67770, ZN => n6021);
   U50313 : OAI22_X1 port map( A1 => n67778, A2 => n63287, B1 => n68080, B2 => 
                           n67770, ZN => n6022);
   U50314 : OAI22_X1 port map( A1 => n67778, A2 => n63286, B1 => n68083, B2 => 
                           n67770, ZN => n6023);
   U50315 : OAI22_X1 port map( A1 => n67778, A2 => n63285, B1 => n68086, B2 => 
                           n67770, ZN => n6024);
   U50316 : OAI22_X1 port map( A1 => n67778, A2 => n63284, B1 => n68089, B2 => 
                           n67770, ZN => n6025);
   U50317 : OAI22_X1 port map( A1 => n67778, A2 => n63283, B1 => n68092, B2 => 
                           n67770, ZN => n6026);
   U50318 : OAI22_X1 port map( A1 => n67779, A2 => n63282, B1 => n68095, B2 => 
                           n67771, ZN => n6027);
   U50319 : OAI22_X1 port map( A1 => n67779, A2 => n63281, B1 => n68098, B2 => 
                           n67771, ZN => n6028);
   U50320 : OAI22_X1 port map( A1 => n67779, A2 => n63280, B1 => n68101, B2 => 
                           n67771, ZN => n6029);
   U50321 : OAI22_X1 port map( A1 => n67779, A2 => n63279, B1 => n68104, B2 => 
                           n67771, ZN => n6030);
   U50322 : OAI22_X1 port map( A1 => n67779, A2 => n63278, B1 => n68107, B2 => 
                           n67771, ZN => n6031);
   U50323 : OAI22_X1 port map( A1 => n67779, A2 => n63277, B1 => n68110, B2 => 
                           n67771, ZN => n6032);
   U50324 : OAI22_X1 port map( A1 => n67779, A2 => n63276, B1 => n68113, B2 => 
                           n67771, ZN => n6033);
   U50325 : OAI22_X1 port map( A1 => n67779, A2 => n63275, B1 => n68116, B2 => 
                           n67771, ZN => n6034);
   U50326 : OAI22_X1 port map( A1 => n67779, A2 => n63274, B1 => n68119, B2 => 
                           n67771, ZN => n6035);
   U50327 : OAI22_X1 port map( A1 => n67779, A2 => n63273, B1 => n68122, B2 => 
                           n67771, ZN => n6036);
   U50328 : OAI22_X1 port map( A1 => n67779, A2 => n63272, B1 => n68125, B2 => 
                           n67771, ZN => n6037);
   U50329 : OAI22_X1 port map( A1 => n67779, A2 => n63271, B1 => n68128, B2 => 
                           n67771, ZN => n6038);
   U50330 : OAI22_X1 port map( A1 => n67779, A2 => n63270, B1 => n68131, B2 => 
                           n67772, ZN => n6039);
   U50331 : OAI22_X1 port map( A1 => n67780, A2 => n63269, B1 => n68134, B2 => 
                           n67772, ZN => n6040);
   U50332 : OAI22_X1 port map( A1 => n67780, A2 => n63268, B1 => n68137, B2 => 
                           n67772, ZN => n6041);
   U50333 : OAI22_X1 port map( A1 => n67780, A2 => n63267, B1 => n68140, B2 => 
                           n67772, ZN => n6042);
   U50334 : OAI22_X1 port map( A1 => n67780, A2 => n63266, B1 => n68143, B2 => 
                           n67772, ZN => n6043);
   U50335 : OAI22_X1 port map( A1 => n67780, A2 => n63265, B1 => n68146, B2 => 
                           n67772, ZN => n6044);
   U50336 : OAI22_X1 port map( A1 => n67780, A2 => n63264, B1 => n68149, B2 => 
                           n67772, ZN => n6045);
   U50337 : OAI22_X1 port map( A1 => n67780, A2 => n63263, B1 => n68152, B2 => 
                           n67772, ZN => n6046);
   U50338 : OAI22_X1 port map( A1 => n67780, A2 => n63262, B1 => n68155, B2 => 
                           n67772, ZN => n6047);
   U50339 : OAI22_X1 port map( A1 => n67780, A2 => n63261, B1 => n68158, B2 => 
                           n67772, ZN => n6048);
   U50340 : OAI22_X1 port map( A1 => n67780, A2 => n63260, B1 => n68161, B2 => 
                           n67772, ZN => n6049);
   U50341 : OAI22_X1 port map( A1 => n67780, A2 => n63259, B1 => n68164, B2 => 
                           n67772, ZN => n6050);
   U50342 : OAI22_X1 port map( A1 => n67780, A2 => n63258, B1 => n68167, B2 => 
                           n67773, ZN => n6051);
   U50343 : OAI22_X1 port map( A1 => n67780, A2 => n63257, B1 => n68170, B2 => 
                           n67773, ZN => n6052);
   U50344 : OAI22_X1 port map( A1 => n67781, A2 => n63256, B1 => n68173, B2 => 
                           n67773, ZN => n6053);
   U50345 : OAI22_X1 port map( A1 => n67781, A2 => n63255, B1 => n68176, B2 => 
                           n67773, ZN => n6054);
   U50346 : OAI22_X1 port map( A1 => n67781, A2 => n63254, B1 => n68179, B2 => 
                           n67773, ZN => n6055);
   U50347 : OAI22_X1 port map( A1 => n67781, A2 => n63253, B1 => n68182, B2 => 
                           n67773, ZN => n6056);
   U50348 : OAI22_X1 port map( A1 => n67781, A2 => n63252, B1 => n68185, B2 => 
                           n67773, ZN => n6057);
   U50349 : OAI22_X1 port map( A1 => n67781, A2 => n63251, B1 => n68188, B2 => 
                           n67773, ZN => n6058);
   U50350 : OAI22_X1 port map( A1 => n67781, A2 => n63250, B1 => n68191, B2 => 
                           n67773, ZN => n6059);
   U50351 : OAI22_X1 port map( A1 => n67781, A2 => n63249, B1 => n68194, B2 => 
                           n67773, ZN => n6060);
   U50352 : OAI22_X1 port map( A1 => n67781, A2 => n63248, B1 => n68197, B2 => 
                           n67773, ZN => n6061);
   U50353 : OAI22_X1 port map( A1 => n67781, A2 => n63247, B1 => n68200, B2 => 
                           n67773, ZN => n6062);
   U50354 : OAI22_X1 port map( A1 => n67781, A2 => n63246, B1 => n68203, B2 => 
                           n67774, ZN => n6063);
   U50355 : OAI22_X1 port map( A1 => n67781, A2 => n63245, B1 => n68206, B2 => 
                           n67774, ZN => n6064);
   U50356 : OAI22_X1 port map( A1 => n67781, A2 => n63244, B1 => n68209, B2 => 
                           n67774, ZN => n6065);
   U50357 : OAI22_X1 port map( A1 => n67782, A2 => n63243, B1 => n68212, B2 => 
                           n67774, ZN => n6066);
   U50358 : OAI22_X1 port map( A1 => n67782, A2 => n63242, B1 => n68215, B2 => 
                           n67774, ZN => n6067);
   U50359 : OAI22_X1 port map( A1 => n67782, A2 => n63241, B1 => n68218, B2 => 
                           n67774, ZN => n6068);
   U50360 : OAI22_X1 port map( A1 => n67782, A2 => n63240, B1 => n68221, B2 => 
                           n67774, ZN => n6069);
   U50361 : OAI22_X1 port map( A1 => n67782, A2 => n63239, B1 => n68224, B2 => 
                           n67774, ZN => n6070);
   U50362 : OAI22_X1 port map( A1 => n67782, A2 => n63238, B1 => n68227, B2 => 
                           n67774, ZN => n6071);
   U50363 : OAI22_X1 port map( A1 => n67782, A2 => n63237, B1 => n68230, B2 => 
                           n67774, ZN => n6072);
   U50364 : OAI22_X1 port map( A1 => n67782, A2 => n63236, B1 => n68233, B2 => 
                           n67774, ZN => n6073);
   U50365 : OAI22_X1 port map( A1 => n67782, A2 => n63235, B1 => n68236, B2 => 
                           n67774, ZN => n6074);
   U50366 : OAI22_X1 port map( A1 => n7489, A2 => n67789, B1 => n68059, B2 => 
                           n67783, ZN => n6079);
   U50367 : OAI22_X1 port map( A1 => n7505, A2 => n67789, B1 => n68062, B2 => 
                           n67783, ZN => n6080);
   U50368 : OAI22_X1 port map( A1 => n7521, A2 => n67789, B1 => n68065, B2 => 
                           n67783, ZN => n6081);
   U50369 : OAI22_X1 port map( A1 => n7537, A2 => n67789, B1 => n68068, B2 => 
                           n67783, ZN => n6082);
   U50370 : OAI22_X1 port map( A1 => n7553, A2 => n67789, B1 => n68071, B2 => 
                           n67783, ZN => n6083);
   U50371 : OAI22_X1 port map( A1 => n7569, A2 => n67789, B1 => n68074, B2 => 
                           n67783, ZN => n6084);
   U50372 : OAI22_X1 port map( A1 => n7585, A2 => n67789, B1 => n68077, B2 => 
                           n67783, ZN => n6085);
   U50373 : OAI22_X1 port map( A1 => n7601, A2 => n67789, B1 => n68080, B2 => 
                           n67783, ZN => n6086);
   U50374 : OAI22_X1 port map( A1 => n7617, A2 => n67789, B1 => n68083, B2 => 
                           n67783, ZN => n6087);
   U50375 : OAI22_X1 port map( A1 => n7633, A2 => n67789, B1 => n68086, B2 => 
                           n67783, ZN => n6088);
   U50376 : OAI22_X1 port map( A1 => n7649, A2 => n67789, B1 => n68089, B2 => 
                           n67783, ZN => n6089);
   U50377 : OAI22_X1 port map( A1 => n7665, A2 => n67790, B1 => n68092, B2 => 
                           n67783, ZN => n6090);
   U50378 : OAI22_X1 port map( A1 => n7681, A2 => n67790, B1 => n68095, B2 => 
                           n67784, ZN => n6091);
   U50379 : OAI22_X1 port map( A1 => n7697, A2 => n67790, B1 => n68098, B2 => 
                           n67784, ZN => n6092);
   U50380 : OAI22_X1 port map( A1 => n7713, A2 => n67790, B1 => n68101, B2 => 
                           n67784, ZN => n6093);
   U50381 : OAI22_X1 port map( A1 => n7729, A2 => n67790, B1 => n68104, B2 => 
                           n67784, ZN => n6094);
   U50382 : OAI22_X1 port map( A1 => n7745, A2 => n67790, B1 => n68107, B2 => 
                           n67784, ZN => n6095);
   U50383 : OAI22_X1 port map( A1 => n7761, A2 => n67790, B1 => n68110, B2 => 
                           n67784, ZN => n6096);
   U50384 : OAI22_X1 port map( A1 => n7777, A2 => n67790, B1 => n68113, B2 => 
                           n67784, ZN => n6097);
   U50385 : OAI22_X1 port map( A1 => n7793, A2 => n67790, B1 => n68116, B2 => 
                           n67784, ZN => n6098);
   U50386 : OAI22_X1 port map( A1 => n7809, A2 => n67790, B1 => n68119, B2 => 
                           n67784, ZN => n6099);
   U50387 : OAI22_X1 port map( A1 => n7825, A2 => n67790, B1 => n68122, B2 => 
                           n67784, ZN => n6100);
   U50388 : OAI22_X1 port map( A1 => n7841, A2 => n67790, B1 => n68125, B2 => 
                           n67784, ZN => n6101);
   U50389 : OAI22_X1 port map( A1 => n7857, A2 => n67791, B1 => n68128, B2 => 
                           n67784, ZN => n6102);
   U50390 : OAI22_X1 port map( A1 => n7873, A2 => n67791, B1 => n68131, B2 => 
                           n67785, ZN => n6103);
   U50391 : OAI22_X1 port map( A1 => n7889, A2 => n67791, B1 => n68134, B2 => 
                           n67785, ZN => n6104);
   U50392 : OAI22_X1 port map( A1 => n7905, A2 => n67791, B1 => n68137, B2 => 
                           n67785, ZN => n6105);
   U50393 : OAI22_X1 port map( A1 => n7921, A2 => n67791, B1 => n68140, B2 => 
                           n67785, ZN => n6106);
   U50394 : OAI22_X1 port map( A1 => n7937, A2 => n67791, B1 => n68143, B2 => 
                           n67785, ZN => n6107);
   U50395 : OAI22_X1 port map( A1 => n7953, A2 => n67791, B1 => n68146, B2 => 
                           n67785, ZN => n6108);
   U50396 : OAI22_X1 port map( A1 => n7969, A2 => n67791, B1 => n68149, B2 => 
                           n67785, ZN => n6109);
   U50397 : OAI22_X1 port map( A1 => n7985, A2 => n67791, B1 => n68152, B2 => 
                           n67785, ZN => n6110);
   U50398 : OAI22_X1 port map( A1 => n8001, A2 => n67791, B1 => n68155, B2 => 
                           n67785, ZN => n6111);
   U50399 : OAI22_X1 port map( A1 => n8017, A2 => n67791, B1 => n68158, B2 => 
                           n67785, ZN => n6112);
   U50400 : OAI22_X1 port map( A1 => n8033, A2 => n67791, B1 => n68161, B2 => 
                           n67785, ZN => n6113);
   U50401 : OAI22_X1 port map( A1 => n8049, A2 => n67792, B1 => n68164, B2 => 
                           n67785, ZN => n6114);
   U50402 : OAI22_X1 port map( A1 => n8065, A2 => n67792, B1 => n68167, B2 => 
                           n67786, ZN => n6115);
   U50403 : OAI22_X1 port map( A1 => n8081, A2 => n67792, B1 => n68170, B2 => 
                           n67786, ZN => n6116);
   U50404 : OAI22_X1 port map( A1 => n8097, A2 => n67792, B1 => n68173, B2 => 
                           n67786, ZN => n6117);
   U50405 : OAI22_X1 port map( A1 => n8113, A2 => n67792, B1 => n68176, B2 => 
                           n67786, ZN => n6118);
   U50406 : OAI22_X1 port map( A1 => n8129, A2 => n67792, B1 => n68179, B2 => 
                           n67786, ZN => n6119);
   U50407 : OAI22_X1 port map( A1 => n8145, A2 => n67792, B1 => n68182, B2 => 
                           n67786, ZN => n6120);
   U50408 : OAI22_X1 port map( A1 => n8161, A2 => n67792, B1 => n68185, B2 => 
                           n67786, ZN => n6121);
   U50409 : OAI22_X1 port map( A1 => n8177, A2 => n67792, B1 => n68188, B2 => 
                           n67786, ZN => n6122);
   U50410 : OAI22_X1 port map( A1 => n8193, A2 => n67792, B1 => n68191, B2 => 
                           n67786, ZN => n6123);
   U50411 : OAI22_X1 port map( A1 => n8209, A2 => n67792, B1 => n68194, B2 => 
                           n67786, ZN => n6124);
   U50412 : OAI22_X1 port map( A1 => n8225, A2 => n67792, B1 => n68197, B2 => 
                           n67786, ZN => n6125);
   U50413 : OAI22_X1 port map( A1 => n8241, A2 => n67793, B1 => n68200, B2 => 
                           n67786, ZN => n6126);
   U50414 : OAI22_X1 port map( A1 => n8257, A2 => n67793, B1 => n68203, B2 => 
                           n67787, ZN => n6127);
   U50415 : OAI22_X1 port map( A1 => n8273, A2 => n67793, B1 => n68206, B2 => 
                           n67787, ZN => n6128);
   U50416 : OAI22_X1 port map( A1 => n8289, A2 => n67793, B1 => n68209, B2 => 
                           n67787, ZN => n6129);
   U50417 : OAI22_X1 port map( A1 => n8305, A2 => n67793, B1 => n68212, B2 => 
                           n67787, ZN => n6130);
   U50418 : OAI22_X1 port map( A1 => n8321, A2 => n67793, B1 => n68215, B2 => 
                           n67787, ZN => n6131);
   U50419 : OAI22_X1 port map( A1 => n8337, A2 => n67793, B1 => n68218, B2 => 
                           n67787, ZN => n6132);
   U50420 : OAI22_X1 port map( A1 => n8353, A2 => n67793, B1 => n68221, B2 => 
                           n67787, ZN => n6133);
   U50421 : OAI22_X1 port map( A1 => n8369, A2 => n67793, B1 => n68224, B2 => 
                           n67787, ZN => n6134);
   U50422 : OAI22_X1 port map( A1 => n8385, A2 => n67793, B1 => n68227, B2 => 
                           n67787, ZN => n6135);
   U50423 : OAI22_X1 port map( A1 => n8401, A2 => n67793, B1 => n68230, B2 => 
                           n67787, ZN => n6136);
   U50424 : OAI22_X1 port map( A1 => n8417, A2 => n67793, B1 => n68233, B2 => 
                           n67787, ZN => n6137);
   U50425 : OAI22_X1 port map( A1 => n8433, A2 => n67794, B1 => n68236, B2 => 
                           n67787, ZN => n6138);
   U50426 : OAI22_X1 port map( A1 => n67893, A2 => n62825, B1 => n68059, B2 => 
                           n67885, ZN => n6591);
   U50427 : OAI22_X1 port map( A1 => n67897, A2 => n62824, B1 => n68062, B2 => 
                           n67885, ZN => n6592);
   U50428 : OAI22_X1 port map( A1 => n67897, A2 => n62823, B1 => n68065, B2 => 
                           n67885, ZN => n6593);
   U50429 : OAI22_X1 port map( A1 => n67897, A2 => n62822, B1 => n68068, B2 => 
                           n67885, ZN => n6594);
   U50430 : OAI22_X1 port map( A1 => n67897, A2 => n62821, B1 => n68071, B2 => 
                           n67885, ZN => n6595);
   U50431 : OAI22_X1 port map( A1 => n67897, A2 => n62820, B1 => n68074, B2 => 
                           n67885, ZN => n6596);
   U50432 : OAI22_X1 port map( A1 => n67897, A2 => n62819, B1 => n68077, B2 => 
                           n67885, ZN => n6597);
   U50433 : OAI22_X1 port map( A1 => n67897, A2 => n62818, B1 => n68080, B2 => 
                           n67885, ZN => n6598);
   U50434 : OAI22_X1 port map( A1 => n67897, A2 => n62817, B1 => n68083, B2 => 
                           n67885, ZN => n6599);
   U50435 : OAI22_X1 port map( A1 => n67897, A2 => n62816, B1 => n68086, B2 => 
                           n67885, ZN => n6600);
   U50436 : OAI22_X1 port map( A1 => n67897, A2 => n62815, B1 => n68089, B2 => 
                           n67885, ZN => n6601);
   U50437 : OAI22_X1 port map( A1 => n67897, A2 => n62814, B1 => n68092, B2 => 
                           n67885, ZN => n6602);
   U50438 : OAI22_X1 port map( A1 => n67897, A2 => n62813, B1 => n68095, B2 => 
                           n67886, ZN => n6603);
   U50439 : OAI22_X1 port map( A1 => n67897, A2 => n62812, B1 => n68098, B2 => 
                           n67886, ZN => n6604);
   U50440 : OAI22_X1 port map( A1 => n67896, A2 => n62811, B1 => n68101, B2 => 
                           n67886, ZN => n6605);
   U50441 : OAI22_X1 port map( A1 => n67896, A2 => n62810, B1 => n68104, B2 => 
                           n67886, ZN => n6606);
   U50442 : OAI22_X1 port map( A1 => n67896, A2 => n62809, B1 => n68107, B2 => 
                           n67886, ZN => n6607);
   U50443 : OAI22_X1 port map( A1 => n67896, A2 => n62808, B1 => n68110, B2 => 
                           n67886, ZN => n6608);
   U50444 : OAI22_X1 port map( A1 => n67896, A2 => n62807, B1 => n68113, B2 => 
                           n67886, ZN => n6609);
   U50445 : OAI22_X1 port map( A1 => n67896, A2 => n62806, B1 => n68116, B2 => 
                           n67886, ZN => n6610);
   U50446 : OAI22_X1 port map( A1 => n67896, A2 => n62805, B1 => n68119, B2 => 
                           n67886, ZN => n6611);
   U50447 : OAI22_X1 port map( A1 => n67896, A2 => n62804, B1 => n68122, B2 => 
                           n67886, ZN => n6612);
   U50448 : OAI22_X1 port map( A1 => n67896, A2 => n62803, B1 => n68125, B2 => 
                           n67886, ZN => n6613);
   U50449 : OAI22_X1 port map( A1 => n67896, A2 => n62802, B1 => n68128, B2 => 
                           n67886, ZN => n6614);
   U50450 : OAI22_X1 port map( A1 => n67896, A2 => n62801, B1 => n68131, B2 => 
                           n67887, ZN => n6615);
   U50451 : OAI22_X1 port map( A1 => n67896, A2 => n62800, B1 => n68134, B2 => 
                           n67887, ZN => n6616);
   U50452 : OAI22_X1 port map( A1 => n67896, A2 => n62799, B1 => n68137, B2 => 
                           n67887, ZN => n6617);
   U50453 : OAI22_X1 port map( A1 => n67895, A2 => n62798, B1 => n68140, B2 => 
                           n67887, ZN => n6618);
   U50454 : OAI22_X1 port map( A1 => n67895, A2 => n62797, B1 => n68143, B2 => 
                           n67887, ZN => n6619);
   U50455 : OAI22_X1 port map( A1 => n67895, A2 => n62796, B1 => n68146, B2 => 
                           n67887, ZN => n6620);
   U50456 : OAI22_X1 port map( A1 => n67895, A2 => n62795, B1 => n68149, B2 => 
                           n67887, ZN => n6621);
   U50457 : OAI22_X1 port map( A1 => n67895, A2 => n62794, B1 => n68152, B2 => 
                           n67887, ZN => n6622);
   U50458 : OAI22_X1 port map( A1 => n67895, A2 => n62793, B1 => n68155, B2 => 
                           n67887, ZN => n6623);
   U50459 : OAI22_X1 port map( A1 => n67895, A2 => n62792, B1 => n68158, B2 => 
                           n67887, ZN => n6624);
   U50460 : OAI22_X1 port map( A1 => n67895, A2 => n62791, B1 => n68161, B2 => 
                           n67887, ZN => n6625);
   U50461 : OAI22_X1 port map( A1 => n67895, A2 => n62790, B1 => n68164, B2 => 
                           n67887, ZN => n6626);
   U50462 : OAI22_X1 port map( A1 => n67895, A2 => n62789, B1 => n68167, B2 => 
                           n67888, ZN => n6627);
   U50463 : OAI22_X1 port map( A1 => n67895, A2 => n62788, B1 => n68170, B2 => 
                           n67888, ZN => n6628);
   U50464 : OAI22_X1 port map( A1 => n67895, A2 => n62787, B1 => n68173, B2 => 
                           n67888, ZN => n6629);
   U50465 : OAI22_X1 port map( A1 => n67894, A2 => n62786, B1 => n68176, B2 => 
                           n67888, ZN => n6630);
   U50466 : OAI22_X1 port map( A1 => n67894, A2 => n62785, B1 => n68179, B2 => 
                           n67888, ZN => n6631);
   U50467 : OAI22_X1 port map( A1 => n67894, A2 => n62784, B1 => n68182, B2 => 
                           n67888, ZN => n6632);
   U50468 : OAI22_X1 port map( A1 => n67894, A2 => n62783, B1 => n68185, B2 => 
                           n67888, ZN => n6633);
   U50469 : OAI22_X1 port map( A1 => n67894, A2 => n62782, B1 => n68188, B2 => 
                           n67888, ZN => n6634);
   U50470 : OAI22_X1 port map( A1 => n67894, A2 => n62781, B1 => n68191, B2 => 
                           n67888, ZN => n6635);
   U50471 : OAI22_X1 port map( A1 => n67894, A2 => n62780, B1 => n68194, B2 => 
                           n67888, ZN => n6636);
   U50472 : OAI22_X1 port map( A1 => n67894, A2 => n62779, B1 => n68197, B2 => 
                           n67888, ZN => n6637);
   U50473 : OAI22_X1 port map( A1 => n67895, A2 => n62778, B1 => n68200, B2 => 
                           n67888, ZN => n6638);
   U50474 : OAI22_X1 port map( A1 => n67894, A2 => n62777, B1 => n68203, B2 => 
                           n67889, ZN => n6639);
   U50475 : OAI22_X1 port map( A1 => n67894, A2 => n62776, B1 => n68206, B2 => 
                           n67889, ZN => n6640);
   U50476 : OAI22_X1 port map( A1 => n67894, A2 => n62775, B1 => n68209, B2 => 
                           n67889, ZN => n6641);
   U50477 : OAI22_X1 port map( A1 => n67894, A2 => n62774, B1 => n68212, B2 => 
                           n67889, ZN => n6642);
   U50478 : OAI22_X1 port map( A1 => n67894, A2 => n62773, B1 => n68215, B2 => 
                           n67889, ZN => n6643);
   U50479 : OAI22_X1 port map( A1 => n67893, A2 => n62772, B1 => n68218, B2 => 
                           n67889, ZN => n6644);
   U50480 : OAI22_X1 port map( A1 => n67893, A2 => n62771, B1 => n68221, B2 => 
                           n67889, ZN => n6645);
   U50481 : OAI22_X1 port map( A1 => n67893, A2 => n62770, B1 => n68224, B2 => 
                           n67889, ZN => n6646);
   U50482 : OAI22_X1 port map( A1 => n67893, A2 => n62769, B1 => n68227, B2 => 
                           n67889, ZN => n6647);
   U50483 : OAI22_X1 port map( A1 => n67893, A2 => n62768, B1 => n68230, B2 => 
                           n67889, ZN => n6648);
   U50484 : OAI22_X1 port map( A1 => n67893, A2 => n62767, B1 => n68233, B2 => 
                           n67889, ZN => n6649);
   U50485 : OAI22_X1 port map( A1 => n67893, A2 => n62766, B1 => n68236, B2 => 
                           n67889, ZN => n6650);
   U50486 : INV_X1 port map( A => ADD_RD2(3), ZN => n66292);
   U50487 : INV_X1 port map( A => ADD_RD1(3), ZN => n65093);
   U50488 : INV_X1 port map( A => ADD_RD2(4), ZN => n66291);
   U50489 : INV_X1 port map( A => ADD_RD1(4), ZN => n65095);
   U50490 : INV_X1 port map( A => ADD_RD2(0), ZN => n66297);
   U50491 : INV_X1 port map( A => ADD_RD1(0), ZN => n65094);
   U50492 : NAND4_X1 port map( A1 => n65151, A2 => n65152, A3 => n65153, A4 => 
                           n65154, ZN => n5373);
   U50493 : NOR4_X1 port map( A1 => n65155, A2 => n65156, A3 => n65157, A4 => 
                           n65158, ZN => n65154);
   U50494 : AOI221_X1 port map( B1 => n67283, B2 => n56531, C1 => n67277, C2 =>
                           n58049, A => n65168, ZN => n65151);
   U50495 : NOR4_X1 port map( A1 => n65163, A2 => n65164, A3 => n65165, A4 => 
                           n65166, ZN => n65153);
   U50496 : NAND4_X1 port map( A1 => n65100, A2 => n65101, A3 => n65102, A4 => 
                           n65103, ZN => n5374);
   U50497 : NOR4_X1 port map( A1 => n65104, A2 => n65105, A3 => n65106, A4 => 
                           n65107, ZN => n65103);
   U50498 : AOI221_X1 port map( B1 => n67283, B2 => n56490, C1 => n67277, C2 =>
                           n58050, A => n65148, ZN => n65100);
   U50499 : NOR4_X1 port map( A1 => n65128, A2 => n65129, A3 => n65130, A4 => 
                           n65131, ZN => n65102);
   U50500 : NAND4_X1 port map( A1 => n66267, A2 => n66268, A3 => n66269, A4 => 
                           n66270, ZN => n5311);
   U50501 : AOI221_X1 port map( B1 => n67278, B2 => n58028, C1 => n67272, C2 =>
                           n58051, A => n66300, ZN => n66267);
   U50502 : NOR4_X1 port map( A1 => n66293, A2 => n66294, A3 => n66295, A4 => 
                           n66296, ZN => n66269);
   U50503 : AOI221_X1 port map( B1 => n67302, B2 => n58731, C1 => n67296, C2 =>
                           n58283, A => n66298, ZN => n66268);
   U50504 : NAND4_X1 port map( A1 => n66249, A2 => n66250, A3 => n66251, A4 => 
                           n66252, ZN => n5312);
   U50505 : AOI221_X1 port map( B1 => n67278, B2 => n57995, C1 => n67272, C2 =>
                           n58052, A => n66266, ZN => n66249);
   U50506 : NOR4_X1 port map( A1 => n66261, A2 => n66262, A3 => n66263, A4 => 
                           n66264, ZN => n66251);
   U50507 : AOI221_X1 port map( B1 => n67302, B2 => n58732, C1 => n67296, C2 =>
                           n58284, A => n66265, ZN => n66250);
   U50508 : NAND4_X1 port map( A1 => n66231, A2 => n66232, A3 => n66233, A4 => 
                           n66234, ZN => n5313);
   U50509 : AOI221_X1 port map( B1 => n67278, B2 => n57971, C1 => n67272, C2 =>
                           n58053, A => n66248, ZN => n66231);
   U50510 : NOR4_X1 port map( A1 => n66243, A2 => n66244, A3 => n66245, A4 => 
                           n66246, ZN => n66233);
   U50511 : AOI221_X1 port map( B1 => n67302, B2 => n58733, C1 => n67296, C2 =>
                           n58285, A => n66247, ZN => n66232);
   U50512 : NAND4_X1 port map( A1 => n66213, A2 => n66214, A3 => n66215, A4 => 
                           n66216, ZN => n5314);
   U50513 : AOI221_X1 port map( B1 => n67278, B2 => n57947, C1 => n67272, C2 =>
                           n58054, A => n66230, ZN => n66213);
   U50514 : NOR4_X1 port map( A1 => n66225, A2 => n66226, A3 => n66227, A4 => 
                           n66228, ZN => n66215);
   U50515 : AOI221_X1 port map( B1 => n67302, B2 => n58734, C1 => n67296, C2 =>
                           n58286, A => n66229, ZN => n66214);
   U50516 : NAND4_X1 port map( A1 => n66195, A2 => n66196, A3 => n66197, A4 => 
                           n66198, ZN => n5315);
   U50517 : AOI221_X1 port map( B1 => n67278, B2 => n57923, C1 => n67272, C2 =>
                           n58055, A => n66212, ZN => n66195);
   U50518 : NOR4_X1 port map( A1 => n66207, A2 => n66208, A3 => n66209, A4 => 
                           n66210, ZN => n66197);
   U50519 : AOI221_X1 port map( B1 => n67302, B2 => n58735, C1 => n67296, C2 =>
                           n58287, A => n66211, ZN => n66196);
   U50520 : NAND4_X1 port map( A1 => n66177, A2 => n66178, A3 => n66179, A4 => 
                           n66180, ZN => n5316);
   U50521 : AOI221_X1 port map( B1 => n67278, B2 => n57899, C1 => n67272, C2 =>
                           n58056, A => n66194, ZN => n66177);
   U50522 : NOR4_X1 port map( A1 => n66189, A2 => n66190, A3 => n66191, A4 => 
                           n66192, ZN => n66179);
   U50523 : AOI221_X1 port map( B1 => n67302, B2 => n58736, C1 => n67296, C2 =>
                           n58288, A => n66193, ZN => n66178);
   U50524 : NAND4_X1 port map( A1 => n66159, A2 => n66160, A3 => n66161, A4 => 
                           n66162, ZN => n5317);
   U50525 : AOI221_X1 port map( B1 => n67278, B2 => n57875, C1 => n67272, C2 =>
                           n58057, A => n66176, ZN => n66159);
   U50526 : NOR4_X1 port map( A1 => n66171, A2 => n66172, A3 => n66173, A4 => 
                           n66174, ZN => n66161);
   U50527 : AOI221_X1 port map( B1 => n67302, B2 => n58737, C1 => n67296, C2 =>
                           n58289, A => n66175, ZN => n66160);
   U50528 : NAND4_X1 port map( A1 => n66141, A2 => n66142, A3 => n66143, A4 => 
                           n66144, ZN => n5318);
   U50529 : AOI221_X1 port map( B1 => n67278, B2 => n57851, C1 => n67272, C2 =>
                           n58058, A => n66158, ZN => n66141);
   U50530 : NOR4_X1 port map( A1 => n66153, A2 => n66154, A3 => n66155, A4 => 
                           n66156, ZN => n66143);
   U50531 : AOI221_X1 port map( B1 => n67302, B2 => n58738, C1 => n67296, C2 =>
                           n58290, A => n66157, ZN => n66142);
   U50532 : NAND4_X1 port map( A1 => n66123, A2 => n66124, A3 => n66125, A4 => 
                           n66126, ZN => n5319);
   U50533 : AOI221_X1 port map( B1 => n67278, B2 => n57827, C1 => n67272, C2 =>
                           n58059, A => n66140, ZN => n66123);
   U50534 : NOR4_X1 port map( A1 => n66135, A2 => n66136, A3 => n66137, A4 => 
                           n66138, ZN => n66125);
   U50535 : AOI221_X1 port map( B1 => n67302, B2 => n58739, C1 => n67296, C2 =>
                           n58291, A => n66139, ZN => n66124);
   U50536 : NAND4_X1 port map( A1 => n66105, A2 => n66106, A3 => n66107, A4 => 
                           n66108, ZN => n5320);
   U50537 : AOI221_X1 port map( B1 => n67278, B2 => n57803, C1 => n67272, C2 =>
                           n58060, A => n66122, ZN => n66105);
   U50538 : NOR4_X1 port map( A1 => n66117, A2 => n66118, A3 => n66119, A4 => 
                           n66120, ZN => n66107);
   U50539 : AOI221_X1 port map( B1 => n67302, B2 => n58740, C1 => n67296, C2 =>
                           n58292, A => n66121, ZN => n66106);
   U50540 : NAND4_X1 port map( A1 => n66087, A2 => n66088, A3 => n66089, A4 => 
                           n66090, ZN => n5321);
   U50541 : AOI221_X1 port map( B1 => n67278, B2 => n57779, C1 => n67272, C2 =>
                           n58061, A => n66104, ZN => n66087);
   U50542 : NOR4_X1 port map( A1 => n66099, A2 => n66100, A3 => n66101, A4 => 
                           n66102, ZN => n66089);
   U50543 : AOI221_X1 port map( B1 => n67302, B2 => n58741, C1 => n67296, C2 =>
                           n58293, A => n66103, ZN => n66088);
   U50544 : NAND4_X1 port map( A1 => n66069, A2 => n66070, A3 => n66071, A4 => 
                           n66072, ZN => n5322);
   U50545 : AOI221_X1 port map( B1 => n67278, B2 => n57755, C1 => n67272, C2 =>
                           n58062, A => n66086, ZN => n66069);
   U50546 : NOR4_X1 port map( A1 => n66081, A2 => n66082, A3 => n66083, A4 => 
                           n66084, ZN => n66071);
   U50547 : AOI221_X1 port map( B1 => n67302, B2 => n58742, C1 => n67296, C2 =>
                           n58294, A => n66085, ZN => n66070);
   U50548 : NAND4_X1 port map( A1 => n66051, A2 => n66052, A3 => n66053, A4 => 
                           n66054, ZN => n5323);
   U50549 : AOI221_X1 port map( B1 => n67279, B2 => n57731, C1 => n67273, C2 =>
                           n58063, A => n66068, ZN => n66051);
   U50550 : NOR4_X1 port map( A1 => n66063, A2 => n66064, A3 => n66065, A4 => 
                           n66066, ZN => n66053);
   U50551 : AOI221_X1 port map( B1 => n67303, B2 => n58667, C1 => n67297, C2 =>
                           n58235, A => n66067, ZN => n66052);
   U50552 : NAND4_X1 port map( A1 => n66033, A2 => n66034, A3 => n66035, A4 => 
                           n66036, ZN => n5324);
   U50553 : AOI221_X1 port map( B1 => n67279, B2 => n57707, C1 => n67273, C2 =>
                           n58064, A => n66050, ZN => n66033);
   U50554 : NOR4_X1 port map( A1 => n66045, A2 => n66046, A3 => n66047, A4 => 
                           n66048, ZN => n66035);
   U50555 : AOI221_X1 port map( B1 => n67303, B2 => n58668, C1 => n67297, C2 =>
                           n58236, A => n66049, ZN => n66034);
   U50556 : NAND4_X1 port map( A1 => n66015, A2 => n66016, A3 => n66017, A4 => 
                           n66018, ZN => n5325);
   U50557 : AOI221_X1 port map( B1 => n67279, B2 => n57683, C1 => n67273, C2 =>
                           n58065, A => n66032, ZN => n66015);
   U50558 : NOR4_X1 port map( A1 => n66027, A2 => n66028, A3 => n66029, A4 => 
                           n66030, ZN => n66017);
   U50559 : AOI221_X1 port map( B1 => n67303, B2 => n58669, C1 => n67297, C2 =>
                           n58237, A => n66031, ZN => n66016);
   U50560 : NAND4_X1 port map( A1 => n65997, A2 => n65998, A3 => n65999, A4 => 
                           n66000, ZN => n5326);
   U50561 : AOI221_X1 port map( B1 => n67279, B2 => n57659, C1 => n67273, C2 =>
                           n58066, A => n66014, ZN => n65997);
   U50562 : NOR4_X1 port map( A1 => n66009, A2 => n66010, A3 => n66011, A4 => 
                           n66012, ZN => n65999);
   U50563 : AOI221_X1 port map( B1 => n67303, B2 => n58670, C1 => n67297, C2 =>
                           n58238, A => n66013, ZN => n65998);
   U50564 : NAND4_X1 port map( A1 => n65979, A2 => n65980, A3 => n65981, A4 => 
                           n65982, ZN => n5327);
   U50565 : AOI221_X1 port map( B1 => n67279, B2 => n57635, C1 => n67273, C2 =>
                           n58067, A => n65996, ZN => n65979);
   U50566 : NOR4_X1 port map( A1 => n65991, A2 => n65992, A3 => n65993, A4 => 
                           n65994, ZN => n65981);
   U50567 : AOI221_X1 port map( B1 => n67303, B2 => n58671, C1 => n67297, C2 =>
                           n58239, A => n65995, ZN => n65980);
   U50568 : NAND4_X1 port map( A1 => n65961, A2 => n65962, A3 => n65963, A4 => 
                           n65964, ZN => n5328);
   U50569 : AOI221_X1 port map( B1 => n67279, B2 => n57611, C1 => n67273, C2 =>
                           n58068, A => n65978, ZN => n65961);
   U50570 : NOR4_X1 port map( A1 => n65973, A2 => n65974, A3 => n65975, A4 => 
                           n65976, ZN => n65963);
   U50571 : AOI221_X1 port map( B1 => n67303, B2 => n58672, C1 => n67297, C2 =>
                           n58240, A => n65977, ZN => n65962);
   U50572 : NAND4_X1 port map( A1 => n65943, A2 => n65944, A3 => n65945, A4 => 
                           n65946, ZN => n5329);
   U50573 : AOI221_X1 port map( B1 => n67279, B2 => n57587, C1 => n67273, C2 =>
                           n58069, A => n65960, ZN => n65943);
   U50574 : NOR4_X1 port map( A1 => n65955, A2 => n65956, A3 => n65957, A4 => 
                           n65958, ZN => n65945);
   U50575 : AOI221_X1 port map( B1 => n67303, B2 => n58673, C1 => n67297, C2 =>
                           n58241, A => n65959, ZN => n65944);
   U50576 : NAND4_X1 port map( A1 => n65925, A2 => n65926, A3 => n65927, A4 => 
                           n65928, ZN => n5330);
   U50577 : AOI221_X1 port map( B1 => n67279, B2 => n57563, C1 => n67273, C2 =>
                           n58070, A => n65942, ZN => n65925);
   U50578 : NOR4_X1 port map( A1 => n65937, A2 => n65938, A3 => n65939, A4 => 
                           n65940, ZN => n65927);
   U50579 : AOI221_X1 port map( B1 => n67303, B2 => n58674, C1 => n67297, C2 =>
                           n58242, A => n65941, ZN => n65926);
   U50580 : NAND4_X1 port map( A1 => n65907, A2 => n65908, A3 => n65909, A4 => 
                           n65910, ZN => n5331);
   U50581 : AOI221_X1 port map( B1 => n67279, B2 => n57539, C1 => n67273, C2 =>
                           n58071, A => n65924, ZN => n65907);
   U50582 : NOR4_X1 port map( A1 => n65919, A2 => n65920, A3 => n65921, A4 => 
                           n65922, ZN => n65909);
   U50583 : AOI221_X1 port map( B1 => n67303, B2 => n58675, C1 => n67297, C2 =>
                           n58243, A => n65923, ZN => n65908);
   U50584 : NAND4_X1 port map( A1 => n65889, A2 => n65890, A3 => n65891, A4 => 
                           n65892, ZN => n5332);
   U50585 : AOI221_X1 port map( B1 => n67279, B2 => n57515, C1 => n67273, C2 =>
                           n58072, A => n65906, ZN => n65889);
   U50586 : NOR4_X1 port map( A1 => n65901, A2 => n65902, A3 => n65903, A4 => 
                           n65904, ZN => n65891);
   U50587 : AOI221_X1 port map( B1 => n67303, B2 => n58676, C1 => n67297, C2 =>
                           n58244, A => n65905, ZN => n65890);
   U50588 : NAND4_X1 port map( A1 => n65871, A2 => n65872, A3 => n65873, A4 => 
                           n65874, ZN => n5333);
   U50589 : AOI221_X1 port map( B1 => n67279, B2 => n57491, C1 => n67273, C2 =>
                           n58073, A => n65888, ZN => n65871);
   U50590 : NOR4_X1 port map( A1 => n65883, A2 => n65884, A3 => n65885, A4 => 
                           n65886, ZN => n65873);
   U50591 : AOI221_X1 port map( B1 => n67303, B2 => n58677, C1 => n67297, C2 =>
                           n58245, A => n65887, ZN => n65872);
   U50592 : NAND4_X1 port map( A1 => n65853, A2 => n65854, A3 => n65855, A4 => 
                           n65856, ZN => n5334);
   U50593 : AOI221_X1 port map( B1 => n67279, B2 => n57467, C1 => n67273, C2 =>
                           n58074, A => n65870, ZN => n65853);
   U50594 : NOR4_X1 port map( A1 => n65865, A2 => n65866, A3 => n65867, A4 => 
                           n65868, ZN => n65855);
   U50595 : AOI221_X1 port map( B1 => n67303, B2 => n58678, C1 => n67297, C2 =>
                           n58246, A => n65869, ZN => n65854);
   U50596 : NAND4_X1 port map( A1 => n65835, A2 => n65836, A3 => n65837, A4 => 
                           n65838, ZN => n5335);
   U50597 : AOI221_X1 port map( B1 => n67280, B2 => n57443, C1 => n67274, C2 =>
                           n58075, A => n65852, ZN => n65835);
   U50598 : NOR4_X1 port map( A1 => n65847, A2 => n65848, A3 => n65849, A4 => 
                           n65850, ZN => n65837);
   U50599 : AOI221_X1 port map( B1 => n67304, B2 => n58679, C1 => n67298, C2 =>
                           n58247, A => n65851, ZN => n65836);
   U50600 : NAND4_X1 port map( A1 => n65817, A2 => n65818, A3 => n65819, A4 => 
                           n65820, ZN => n5336);
   U50601 : AOI221_X1 port map( B1 => n67280, B2 => n57419, C1 => n67274, C2 =>
                           n58076, A => n65834, ZN => n65817);
   U50602 : NOR4_X1 port map( A1 => n65829, A2 => n65830, A3 => n65831, A4 => 
                           n65832, ZN => n65819);
   U50603 : AOI221_X1 port map( B1 => n67304, B2 => n58680, C1 => n67298, C2 =>
                           n58248, A => n65833, ZN => n65818);
   U50604 : NAND4_X1 port map( A1 => n65799, A2 => n65800, A3 => n65801, A4 => 
                           n65802, ZN => n5337);
   U50605 : AOI221_X1 port map( B1 => n67280, B2 => n57395, C1 => n67274, C2 =>
                           n58077, A => n65816, ZN => n65799);
   U50606 : NOR4_X1 port map( A1 => n65811, A2 => n65812, A3 => n65813, A4 => 
                           n65814, ZN => n65801);
   U50607 : AOI221_X1 port map( B1 => n67304, B2 => n58681, C1 => n67298, C2 =>
                           n58249, A => n65815, ZN => n65800);
   U50608 : NAND4_X1 port map( A1 => n65781, A2 => n65782, A3 => n65783, A4 => 
                           n65784, ZN => n5338);
   U50609 : AOI221_X1 port map( B1 => n67280, B2 => n57371, C1 => n67274, C2 =>
                           n58078, A => n65798, ZN => n65781);
   U50610 : NOR4_X1 port map( A1 => n65793, A2 => n65794, A3 => n65795, A4 => 
                           n65796, ZN => n65783);
   U50611 : AOI221_X1 port map( B1 => n67304, B2 => n58682, C1 => n67298, C2 =>
                           n58250, A => n65797, ZN => n65782);
   U50612 : NAND4_X1 port map( A1 => n65763, A2 => n65764, A3 => n65765, A4 => 
                           n65766, ZN => n5339);
   U50613 : AOI221_X1 port map( B1 => n67280, B2 => n57347, C1 => n67274, C2 =>
                           n58079, A => n65780, ZN => n65763);
   U50614 : NOR4_X1 port map( A1 => n65775, A2 => n65776, A3 => n65777, A4 => 
                           n65778, ZN => n65765);
   U50615 : AOI221_X1 port map( B1 => n67304, B2 => n58683, C1 => n67298, C2 =>
                           n58251, A => n65779, ZN => n65764);
   U50616 : NAND4_X1 port map( A1 => n65745, A2 => n65746, A3 => n65747, A4 => 
                           n65748, ZN => n5340);
   U50617 : AOI221_X1 port map( B1 => n67280, B2 => n57323, C1 => n67274, C2 =>
                           n58080, A => n65762, ZN => n65745);
   U50618 : NOR4_X1 port map( A1 => n65757, A2 => n65758, A3 => n65759, A4 => 
                           n65760, ZN => n65747);
   U50619 : AOI221_X1 port map( B1 => n67304, B2 => n58684, C1 => n67298, C2 =>
                           n58252, A => n65761, ZN => n65746);
   U50620 : NAND4_X1 port map( A1 => n65727, A2 => n65728, A3 => n65729, A4 => 
                           n65730, ZN => n5341);
   U50621 : AOI221_X1 port map( B1 => n67280, B2 => n57299, C1 => n67274, C2 =>
                           n58081, A => n65744, ZN => n65727);
   U50622 : NOR4_X1 port map( A1 => n65739, A2 => n65740, A3 => n65741, A4 => 
                           n65742, ZN => n65729);
   U50623 : AOI221_X1 port map( B1 => n67304, B2 => n58685, C1 => n67298, C2 =>
                           n58253, A => n65743, ZN => n65728);
   U50624 : NAND4_X1 port map( A1 => n65709, A2 => n65710, A3 => n65711, A4 => 
                           n65712, ZN => n5342);
   U50625 : AOI221_X1 port map( B1 => n67280, B2 => n57275, C1 => n67274, C2 =>
                           n58082, A => n65726, ZN => n65709);
   U50626 : NOR4_X1 port map( A1 => n65721, A2 => n65722, A3 => n65723, A4 => 
                           n65724, ZN => n65711);
   U50627 : AOI221_X1 port map( B1 => n67304, B2 => n58686, C1 => n67298, C2 =>
                           n58254, A => n65725, ZN => n65710);
   U50628 : NAND4_X1 port map( A1 => n65691, A2 => n65692, A3 => n65693, A4 => 
                           n65694, ZN => n5343);
   U50629 : AOI221_X1 port map( B1 => n67280, B2 => n57251, C1 => n67274, C2 =>
                           n58083, A => n65708, ZN => n65691);
   U50630 : NOR4_X1 port map( A1 => n65703, A2 => n65704, A3 => n65705, A4 => 
                           n65706, ZN => n65693);
   U50631 : AOI221_X1 port map( B1 => n67304, B2 => n58687, C1 => n67298, C2 =>
                           n58255, A => n65707, ZN => n65692);
   U50632 : NAND4_X1 port map( A1 => n65673, A2 => n65674, A3 => n65675, A4 => 
                           n65676, ZN => n5344);
   U50633 : AOI221_X1 port map( B1 => n67280, B2 => n57227, C1 => n67274, C2 =>
                           n58084, A => n65690, ZN => n65673);
   U50634 : NOR4_X1 port map( A1 => n65685, A2 => n65686, A3 => n65687, A4 => 
                           n65688, ZN => n65675);
   U50635 : AOI221_X1 port map( B1 => n67304, B2 => n58688, C1 => n67298, C2 =>
                           n58256, A => n65689, ZN => n65674);
   U50636 : NAND4_X1 port map( A1 => n65655, A2 => n65656, A3 => n65657, A4 => 
                           n65658, ZN => n5345);
   U50637 : AOI221_X1 port map( B1 => n67280, B2 => n57203, C1 => n67274, C2 =>
                           n58085, A => n65672, ZN => n65655);
   U50638 : NOR4_X1 port map( A1 => n65667, A2 => n65668, A3 => n65669, A4 => 
                           n65670, ZN => n65657);
   U50639 : AOI221_X1 port map( B1 => n67304, B2 => n58689, C1 => n67298, C2 =>
                           n58257, A => n65671, ZN => n65656);
   U50640 : NAND4_X1 port map( A1 => n65637, A2 => n65638, A3 => n65639, A4 => 
                           n65640, ZN => n5346);
   U50641 : AOI221_X1 port map( B1 => n67280, B2 => n57179, C1 => n67274, C2 =>
                           n58086, A => n65654, ZN => n65637);
   U50642 : NOR4_X1 port map( A1 => n65649, A2 => n65650, A3 => n65651, A4 => 
                           n65652, ZN => n65639);
   U50643 : AOI221_X1 port map( B1 => n67304, B2 => n58690, C1 => n67298, C2 =>
                           n58258, A => n65653, ZN => n65638);
   U50644 : NAND4_X1 port map( A1 => n65619, A2 => n65620, A3 => n65621, A4 => 
                           n65622, ZN => n5347);
   U50645 : AOI221_X1 port map( B1 => n67281, B2 => n57155, C1 => n67275, C2 =>
                           n58087, A => n65636, ZN => n65619);
   U50646 : NOR4_X1 port map( A1 => n65631, A2 => n65632, A3 => n65633, A4 => 
                           n65634, ZN => n65621);
   U50647 : AOI221_X1 port map( B1 => n67305, B2 => n58691, C1 => n67299, C2 =>
                           n58259, A => n65635, ZN => n65620);
   U50648 : NAND4_X1 port map( A1 => n65601, A2 => n65602, A3 => n65603, A4 => 
                           n65604, ZN => n5348);
   U50649 : AOI221_X1 port map( B1 => n67281, B2 => n57131, C1 => n67275, C2 =>
                           n58088, A => n65618, ZN => n65601);
   U50650 : NOR4_X1 port map( A1 => n65613, A2 => n65614, A3 => n65615, A4 => 
                           n65616, ZN => n65603);
   U50651 : AOI221_X1 port map( B1 => n67305, B2 => n58692, C1 => n67299, C2 =>
                           n58260, A => n65617, ZN => n65602);
   U50652 : NAND4_X1 port map( A1 => n65583, A2 => n65584, A3 => n65585, A4 => 
                           n65586, ZN => n5349);
   U50653 : AOI221_X1 port map( B1 => n67281, B2 => n57107, C1 => n67275, C2 =>
                           n58089, A => n65600, ZN => n65583);
   U50654 : NOR4_X1 port map( A1 => n65595, A2 => n65596, A3 => n65597, A4 => 
                           n65598, ZN => n65585);
   U50655 : AOI221_X1 port map( B1 => n67305, B2 => n58693, C1 => n67299, C2 =>
                           n58261, A => n65599, ZN => n65584);
   U50656 : NAND4_X1 port map( A1 => n65565, A2 => n65566, A3 => n65567, A4 => 
                           n65568, ZN => n5350);
   U50657 : AOI221_X1 port map( B1 => n67281, B2 => n57083, C1 => n67275, C2 =>
                           n58090, A => n65582, ZN => n65565);
   U50658 : NOR4_X1 port map( A1 => n65577, A2 => n65578, A3 => n65579, A4 => 
                           n65580, ZN => n65567);
   U50659 : AOI221_X1 port map( B1 => n67305, B2 => n58694, C1 => n67299, C2 =>
                           n58262, A => n65581, ZN => n65566);
   U50660 : NAND4_X1 port map( A1 => n65547, A2 => n65548, A3 => n65549, A4 => 
                           n65550, ZN => n5351);
   U50661 : AOI221_X1 port map( B1 => n67281, B2 => n57059, C1 => n67275, C2 =>
                           n58091, A => n65564, ZN => n65547);
   U50662 : NOR4_X1 port map( A1 => n65559, A2 => n65560, A3 => n65561, A4 => 
                           n65562, ZN => n65549);
   U50663 : AOI221_X1 port map( B1 => n67305, B2 => n58695, C1 => n67299, C2 =>
                           n58263, A => n65563, ZN => n65548);
   U50664 : NAND4_X1 port map( A1 => n65529, A2 => n65530, A3 => n65531, A4 => 
                           n65532, ZN => n5352);
   U50665 : AOI221_X1 port map( B1 => n67281, B2 => n57035, C1 => n67275, C2 =>
                           n58092, A => n65546, ZN => n65529);
   U50666 : NOR4_X1 port map( A1 => n65541, A2 => n65542, A3 => n65543, A4 => 
                           n65544, ZN => n65531);
   U50667 : AOI221_X1 port map( B1 => n67305, B2 => n58696, C1 => n67299, C2 =>
                           n58264, A => n65545, ZN => n65530);
   U50668 : NAND4_X1 port map( A1 => n65511, A2 => n65512, A3 => n65513, A4 => 
                           n65514, ZN => n5353);
   U50669 : AOI221_X1 port map( B1 => n67281, B2 => n57011, C1 => n67275, C2 =>
                           n58093, A => n65528, ZN => n65511);
   U50670 : NOR4_X1 port map( A1 => n65523, A2 => n65524, A3 => n65525, A4 => 
                           n65526, ZN => n65513);
   U50671 : AOI221_X1 port map( B1 => n67305, B2 => n58697, C1 => n67299, C2 =>
                           n58265, A => n65527, ZN => n65512);
   U50672 : NAND4_X1 port map( A1 => n65493, A2 => n65494, A3 => n65495, A4 => 
                           n65496, ZN => n5354);
   U50673 : AOI221_X1 port map( B1 => n67281, B2 => n56987, C1 => n67275, C2 =>
                           n58094, A => n65510, ZN => n65493);
   U50674 : NOR4_X1 port map( A1 => n65505, A2 => n65506, A3 => n65507, A4 => 
                           n65508, ZN => n65495);
   U50675 : AOI221_X1 port map( B1 => n67305, B2 => n58698, C1 => n67299, C2 =>
                           n58266, A => n65509, ZN => n65494);
   U50676 : NAND4_X1 port map( A1 => n65475, A2 => n65476, A3 => n65477, A4 => 
                           n65478, ZN => n5355);
   U50677 : AOI221_X1 port map( B1 => n67281, B2 => n56963, C1 => n67275, C2 =>
                           n58095, A => n65492, ZN => n65475);
   U50678 : NOR4_X1 port map( A1 => n65487, A2 => n65488, A3 => n65489, A4 => 
                           n65490, ZN => n65477);
   U50679 : AOI221_X1 port map( B1 => n67305, B2 => n58699, C1 => n67299, C2 =>
                           n58267, A => n65491, ZN => n65476);
   U50680 : NAND4_X1 port map( A1 => n65457, A2 => n65458, A3 => n65459, A4 => 
                           n65460, ZN => n5356);
   U50681 : AOI221_X1 port map( B1 => n67281, B2 => n56939, C1 => n67275, C2 =>
                           n58096, A => n65474, ZN => n65457);
   U50682 : NOR4_X1 port map( A1 => n65469, A2 => n65470, A3 => n65471, A4 => 
                           n65472, ZN => n65459);
   U50683 : AOI221_X1 port map( B1 => n67305, B2 => n58700, C1 => n67299, C2 =>
                           n58268, A => n65473, ZN => n65458);
   U50684 : NAND4_X1 port map( A1 => n65439, A2 => n65440, A3 => n65441, A4 => 
                           n65442, ZN => n5357);
   U50685 : AOI221_X1 port map( B1 => n67281, B2 => n56915, C1 => n67275, C2 =>
                           n58097, A => n65456, ZN => n65439);
   U50686 : NOR4_X1 port map( A1 => n65451, A2 => n65452, A3 => n65453, A4 => 
                           n65454, ZN => n65441);
   U50687 : AOI221_X1 port map( B1 => n67305, B2 => n58701, C1 => n67299, C2 =>
                           n58269, A => n65455, ZN => n65440);
   U50688 : NAND4_X1 port map( A1 => n65421, A2 => n65422, A3 => n65423, A4 => 
                           n65424, ZN => n5358);
   U50689 : AOI221_X1 port map( B1 => n67281, B2 => n56891, C1 => n67275, C2 =>
                           n58098, A => n65438, ZN => n65421);
   U50690 : NOR4_X1 port map( A1 => n65433, A2 => n65434, A3 => n65435, A4 => 
                           n65436, ZN => n65423);
   U50691 : AOI221_X1 port map( B1 => n67305, B2 => n58702, C1 => n67299, C2 =>
                           n58270, A => n65437, ZN => n65422);
   U50692 : NAND4_X1 port map( A1 => n65403, A2 => n65404, A3 => n65405, A4 => 
                           n65406, ZN => n5359);
   U50693 : AOI221_X1 port map( B1 => n67282, B2 => n56867, C1 => n67276, C2 =>
                           n58099, A => n65420, ZN => n65403);
   U50694 : NOR4_X1 port map( A1 => n65415, A2 => n65416, A3 => n65417, A4 => 
                           n65418, ZN => n65405);
   U50695 : AOI221_X1 port map( B1 => n67306, B2 => n58703, C1 => n67300, C2 =>
                           n58271, A => n65419, ZN => n65404);
   U50696 : NAND4_X1 port map( A1 => n65385, A2 => n65386, A3 => n65387, A4 => 
                           n65388, ZN => n5360);
   U50697 : AOI221_X1 port map( B1 => n67282, B2 => n56843, C1 => n67276, C2 =>
                           n58100, A => n65402, ZN => n65385);
   U50698 : NOR4_X1 port map( A1 => n65397, A2 => n65398, A3 => n65399, A4 => 
                           n65400, ZN => n65387);
   U50699 : AOI221_X1 port map( B1 => n67306, B2 => n58704, C1 => n67300, C2 =>
                           n58272, A => n65401, ZN => n65386);
   U50700 : NAND4_X1 port map( A1 => n65367, A2 => n65368, A3 => n65369, A4 => 
                           n65370, ZN => n5361);
   U50701 : AOI221_X1 port map( B1 => n67282, B2 => n56819, C1 => n67276, C2 =>
                           n58101, A => n65384, ZN => n65367);
   U50702 : NOR4_X1 port map( A1 => n65379, A2 => n65380, A3 => n65381, A4 => 
                           n65382, ZN => n65369);
   U50703 : AOI221_X1 port map( B1 => n67306, B2 => n58705, C1 => n67300, C2 =>
                           n58273, A => n65383, ZN => n65368);
   U50704 : NAND4_X1 port map( A1 => n65349, A2 => n65350, A3 => n65351, A4 => 
                           n65352, ZN => n5362);
   U50705 : AOI221_X1 port map( B1 => n67282, B2 => n56795, C1 => n67276, C2 =>
                           n58102, A => n65366, ZN => n65349);
   U50706 : NOR4_X1 port map( A1 => n65361, A2 => n65362, A3 => n65363, A4 => 
                           n65364, ZN => n65351);
   U50707 : AOI221_X1 port map( B1 => n67306, B2 => n58706, C1 => n67300, C2 =>
                           n58274, A => n65365, ZN => n65350);
   U50708 : NAND4_X1 port map( A1 => n65331, A2 => n65332, A3 => n65333, A4 => 
                           n65334, ZN => n5363);
   U50709 : AOI221_X1 port map( B1 => n67282, B2 => n56771, C1 => n67276, C2 =>
                           n58103, A => n65348, ZN => n65331);
   U50710 : NOR4_X1 port map( A1 => n65343, A2 => n65344, A3 => n65345, A4 => 
                           n65346, ZN => n65333);
   U50711 : AOI221_X1 port map( B1 => n67306, B2 => n58707, C1 => n67300, C2 =>
                           n58275, A => n65347, ZN => n65332);
   U50712 : NAND4_X1 port map( A1 => n65313, A2 => n65314, A3 => n65315, A4 => 
                           n65316, ZN => n5364);
   U50713 : AOI221_X1 port map( B1 => n67282, B2 => n56747, C1 => n67276, C2 =>
                           n58104, A => n65330, ZN => n65313);
   U50714 : NOR4_X1 port map( A1 => n65325, A2 => n65326, A3 => n65327, A4 => 
                           n65328, ZN => n65315);
   U50715 : AOI221_X1 port map( B1 => n67306, B2 => n58708, C1 => n67300, C2 =>
                           n58276, A => n65329, ZN => n65314);
   U50716 : NAND4_X1 port map( A1 => n65295, A2 => n65296, A3 => n65297, A4 => 
                           n65298, ZN => n5365);
   U50717 : AOI221_X1 port map( B1 => n67282, B2 => n56723, C1 => n67276, C2 =>
                           n58105, A => n65312, ZN => n65295);
   U50718 : NOR4_X1 port map( A1 => n65307, A2 => n65308, A3 => n65309, A4 => 
                           n65310, ZN => n65297);
   U50719 : AOI221_X1 port map( B1 => n67306, B2 => n58709, C1 => n67300, C2 =>
                           n58277, A => n65311, ZN => n65296);
   U50720 : NAND4_X1 port map( A1 => n65277, A2 => n65278, A3 => n65279, A4 => 
                           n65280, ZN => n5366);
   U50721 : AOI221_X1 port map( B1 => n67282, B2 => n56699, C1 => n67276, C2 =>
                           n58106, A => n65294, ZN => n65277);
   U50722 : NOR4_X1 port map( A1 => n65289, A2 => n65290, A3 => n65291, A4 => 
                           n65292, ZN => n65279);
   U50723 : AOI221_X1 port map( B1 => n67306, B2 => n58710, C1 => n67300, C2 =>
                           n58278, A => n65293, ZN => n65278);
   U50724 : NAND4_X1 port map( A1 => n65259, A2 => n65260, A3 => n65261, A4 => 
                           n65262, ZN => n5367);
   U50725 : AOI221_X1 port map( B1 => n67282, B2 => n56675, C1 => n67276, C2 =>
                           n58107, A => n65276, ZN => n65259);
   U50726 : NOR4_X1 port map( A1 => n65271, A2 => n65272, A3 => n65273, A4 => 
                           n65274, ZN => n65261);
   U50727 : AOI221_X1 port map( B1 => n67306, B2 => n58711, C1 => n67300, C2 =>
                           n58279, A => n65275, ZN => n65260);
   U50728 : NAND4_X1 port map( A1 => n65241, A2 => n65242, A3 => n65243, A4 => 
                           n65244, ZN => n5368);
   U50729 : AOI221_X1 port map( B1 => n67282, B2 => n56651, C1 => n67276, C2 =>
                           n58108, A => n65258, ZN => n65241);
   U50730 : NOR4_X1 port map( A1 => n65253, A2 => n65254, A3 => n65255, A4 => 
                           n65256, ZN => n65243);
   U50731 : AOI221_X1 port map( B1 => n67306, B2 => n58712, C1 => n67300, C2 =>
                           n58280, A => n65257, ZN => n65242);
   U50732 : NAND4_X1 port map( A1 => n65223, A2 => n65224, A3 => n65225, A4 => 
                           n65226, ZN => n5369);
   U50733 : AOI221_X1 port map( B1 => n67282, B2 => n56627, C1 => n67276, C2 =>
                           n58109, A => n65240, ZN => n65223);
   U50734 : NOR4_X1 port map( A1 => n65235, A2 => n65236, A3 => n65237, A4 => 
                           n65238, ZN => n65225);
   U50735 : AOI221_X1 port map( B1 => n67306, B2 => n58713, C1 => n67300, C2 =>
                           n58281, A => n65239, ZN => n65224);
   U50736 : NAND4_X1 port map( A1 => n65205, A2 => n65206, A3 => n65207, A4 => 
                           n65208, ZN => n5370);
   U50737 : AOI221_X1 port map( B1 => n67282, B2 => n56603, C1 => n67276, C2 =>
                           n58110, A => n65222, ZN => n65205);
   U50738 : NOR4_X1 port map( A1 => n65217, A2 => n65218, A3 => n65219, A4 => 
                           n65220, ZN => n65207);
   U50739 : AOI221_X1 port map( B1 => n67306, B2 => n58714, C1 => n67300, C2 =>
                           n58282, A => n65221, ZN => n65206);
   U50740 : NAND4_X1 port map( A1 => n65187, A2 => n65188, A3 => n65189, A4 => 
                           n65190, ZN => n5371);
   U50741 : NOR4_X1 port map( A1 => n65191, A2 => n65192, A3 => n65193, A4 => 
                           n65194, ZN => n65190);
   U50742 : AOI221_X1 port map( B1 => n67283, B2 => n56579, C1 => n67277, C2 =>
                           n58047, A => n65204, ZN => n65187);
   U50743 : NOR4_X1 port map( A1 => n65199, A2 => n65200, A3 => n65201, A4 => 
                           n65202, ZN => n65189);
   U50744 : NAND4_X1 port map( A1 => n65169, A2 => n65170, A3 => n65171, A4 => 
                           n65172, ZN => n5372);
   U50745 : NOR4_X1 port map( A1 => n65173, A2 => n65174, A3 => n65175, A4 => 
                           n65176, ZN => n65172);
   U50746 : AOI221_X1 port map( B1 => n67283, B2 => n56555, C1 => n67277, C2 =>
                           n58048, A => n65186, ZN => n65169);
   U50747 : NOR4_X1 port map( A1 => n65181, A2 => n65182, A3 => n65183, A4 => 
                           n65184, ZN => n65171);
   U50748 : NAND4_X1 port map( A1 => n65064, A2 => n65065, A3 => n65066, A4 => 
                           n65067, ZN => n5375);
   U50749 : AOI221_X1 port map( B1 => n67476, B2 => n58028, C1 => n67470, C2 =>
                           n59029, A => n65098, ZN => n65064);
   U50750 : AOI221_X1 port map( B1 => n67500, B2 => n66313, C1 => n67494, C2 =>
                           n58112, A => n65096, ZN => n65065);
   U50751 : NOR4_X1 port map( A1 => n65089, A2 => n65090, A3 => n65091, A4 => 
                           n65092, ZN => n65066);
   U50752 : NAND4_X1 port map( A1 => n65044, A2 => n65045, A3 => n65046, A4 => 
                           n65047, ZN => n5377);
   U50753 : AOI221_X1 port map( B1 => n67476, B2 => n57995, C1 => n67470, C2 =>
                           n59030, A => n65062, ZN => n65044);
   U50754 : AOI221_X1 port map( B1 => n67500, B2 => n66314, C1 => n67494, C2 =>
                           n58114, A => n65061, ZN => n65045);
   U50755 : NOR4_X1 port map( A1 => n65057, A2 => n65058, A3 => n65059, A4 => 
                           n65060, ZN => n65046);
   U50756 : NAND4_X1 port map( A1 => n65024, A2 => n65025, A3 => n65026, A4 => 
                           n65027, ZN => n5379);
   U50757 : AOI221_X1 port map( B1 => n67476, B2 => n57971, C1 => n67470, C2 =>
                           n59031, A => n65042, ZN => n65024);
   U50758 : AOI221_X1 port map( B1 => n67500, B2 => n66315, C1 => n67494, C2 =>
                           n58116, A => n65041, ZN => n65025);
   U50759 : NOR4_X1 port map( A1 => n65037, A2 => n65038, A3 => n65039, A4 => 
                           n65040, ZN => n65026);
   U50760 : NAND4_X1 port map( A1 => n65004, A2 => n65005, A3 => n65006, A4 => 
                           n65007, ZN => n5381);
   U50761 : AOI221_X1 port map( B1 => n67476, B2 => n57947, C1 => n67470, C2 =>
                           n59032, A => n65022, ZN => n65004);
   U50762 : AOI221_X1 port map( B1 => n67500, B2 => n66316, C1 => n67494, C2 =>
                           n58118, A => n65021, ZN => n65005);
   U50763 : NOR4_X1 port map( A1 => n65017, A2 => n65018, A3 => n65019, A4 => 
                           n65020, ZN => n65006);
   U50764 : NAND4_X1 port map( A1 => n64984, A2 => n64985, A3 => n64986, A4 => 
                           n64987, ZN => n5383);
   U50765 : AOI221_X1 port map( B1 => n67476, B2 => n57923, C1 => n67470, C2 =>
                           n59033, A => n65002, ZN => n64984);
   U50766 : AOI221_X1 port map( B1 => n67500, B2 => n66317, C1 => n67494, C2 =>
                           n58120, A => n65001, ZN => n64985);
   U50767 : NOR4_X1 port map( A1 => n64997, A2 => n64998, A3 => n64999, A4 => 
                           n65000, ZN => n64986);
   U50768 : NAND4_X1 port map( A1 => n64964, A2 => n64965, A3 => n64966, A4 => 
                           n64967, ZN => n5385);
   U50769 : AOI221_X1 port map( B1 => n67476, B2 => n57899, C1 => n67470, C2 =>
                           n59034, A => n64982, ZN => n64964);
   U50770 : AOI221_X1 port map( B1 => n67500, B2 => n66318, C1 => n67494, C2 =>
                           n58122, A => n64981, ZN => n64965);
   U50771 : NOR4_X1 port map( A1 => n64977, A2 => n64978, A3 => n64979, A4 => 
                           n64980, ZN => n64966);
   U50772 : NAND4_X1 port map( A1 => n64944, A2 => n64945, A3 => n64946, A4 => 
                           n64947, ZN => n5387);
   U50773 : AOI221_X1 port map( B1 => n67476, B2 => n57875, C1 => n67470, C2 =>
                           n59035, A => n64962, ZN => n64944);
   U50774 : AOI221_X1 port map( B1 => n67500, B2 => n66319, C1 => n67494, C2 =>
                           n58124, A => n64961, ZN => n64945);
   U50775 : NOR4_X1 port map( A1 => n64957, A2 => n64958, A3 => n64959, A4 => 
                           n64960, ZN => n64946);
   U50776 : NAND4_X1 port map( A1 => n64924, A2 => n64925, A3 => n64926, A4 => 
                           n64927, ZN => n5389);
   U50777 : AOI221_X1 port map( B1 => n67476, B2 => n57851, C1 => n67470, C2 =>
                           n59036, A => n64942, ZN => n64924);
   U50778 : AOI221_X1 port map( B1 => n67500, B2 => n66320, C1 => n67494, C2 =>
                           n58126, A => n64941, ZN => n64925);
   U50779 : NOR4_X1 port map( A1 => n64937, A2 => n64938, A3 => n64939, A4 => 
                           n64940, ZN => n64926);
   U50780 : NAND4_X1 port map( A1 => n64904, A2 => n64905, A3 => n64906, A4 => 
                           n64907, ZN => n5391);
   U50781 : AOI221_X1 port map( B1 => n67476, B2 => n57827, C1 => n67470, C2 =>
                           n59037, A => n64922, ZN => n64904);
   U50782 : AOI221_X1 port map( B1 => n67500, B2 => n66321, C1 => n67494, C2 =>
                           n58128, A => n64921, ZN => n64905);
   U50783 : NOR4_X1 port map( A1 => n64917, A2 => n64918, A3 => n64919, A4 => 
                           n64920, ZN => n64906);
   U50784 : NAND4_X1 port map( A1 => n64884, A2 => n64885, A3 => n64886, A4 => 
                           n64887, ZN => n5393);
   U50785 : AOI221_X1 port map( B1 => n67476, B2 => n57803, C1 => n67470, C2 =>
                           n59038, A => n64902, ZN => n64884);
   U50786 : AOI221_X1 port map( B1 => n67500, B2 => n66322, C1 => n67494, C2 =>
                           n58130, A => n64901, ZN => n64885);
   U50787 : NOR4_X1 port map( A1 => n64897, A2 => n64898, A3 => n64899, A4 => 
                           n64900, ZN => n64886);
   U50788 : NAND4_X1 port map( A1 => n64864, A2 => n64865, A3 => n64866, A4 => 
                           n64867, ZN => n5395);
   U50789 : AOI221_X1 port map( B1 => n67476, B2 => n57779, C1 => n67470, C2 =>
                           n59039, A => n64882, ZN => n64864);
   U50790 : AOI221_X1 port map( B1 => n67500, B2 => n66323, C1 => n67494, C2 =>
                           n58132, A => n64881, ZN => n64865);
   U50791 : NOR4_X1 port map( A1 => n64877, A2 => n64878, A3 => n64879, A4 => 
                           n64880, ZN => n64866);
   U50792 : NAND4_X1 port map( A1 => n64844, A2 => n64845, A3 => n64846, A4 => 
                           n64847, ZN => n5397);
   U50793 : AOI221_X1 port map( B1 => n67476, B2 => n57755, C1 => n67470, C2 =>
                           n59040, A => n64862, ZN => n64844);
   U50794 : AOI221_X1 port map( B1 => n67500, B2 => n66324, C1 => n67494, C2 =>
                           n58134, A => n64861, ZN => n64845);
   U50795 : NOR4_X1 port map( A1 => n64857, A2 => n64858, A3 => n64859, A4 => 
                           n64860, ZN => n64846);
   U50796 : NAND4_X1 port map( A1 => n64824, A2 => n64825, A3 => n64826, A4 => 
                           n64827, ZN => n5399);
   U50797 : AOI221_X1 port map( B1 => n67477, B2 => n57731, C1 => n67471, C2 =>
                           n59041, A => n64842, ZN => n64824);
   U50798 : AOI221_X1 port map( B1 => n67501, B2 => n66325, C1 => n67495, C2 =>
                           n58135, A => n64841, ZN => n64825);
   U50799 : NOR4_X1 port map( A1 => n64837, A2 => n64838, A3 => n64839, A4 => 
                           n64840, ZN => n64826);
   U50800 : NAND4_X1 port map( A1 => n64804, A2 => n64805, A3 => n64806, A4 => 
                           n64807, ZN => n5401);
   U50801 : AOI221_X1 port map( B1 => n67477, B2 => n57707, C1 => n67471, C2 =>
                           n59042, A => n64822, ZN => n64804);
   U50802 : AOI221_X1 port map( B1 => n67501, B2 => n66326, C1 => n67495, C2 =>
                           n58137, A => n64821, ZN => n64805);
   U50803 : NOR4_X1 port map( A1 => n64817, A2 => n64818, A3 => n64819, A4 => 
                           n64820, ZN => n64806);
   U50804 : NAND4_X1 port map( A1 => n64784, A2 => n64785, A3 => n64786, A4 => 
                           n64787, ZN => n5403);
   U50805 : AOI221_X1 port map( B1 => n67477, B2 => n57683, C1 => n67471, C2 =>
                           n59043, A => n64802, ZN => n64784);
   U50806 : AOI221_X1 port map( B1 => n67501, B2 => n66327, C1 => n67495, C2 =>
                           n58139, A => n64801, ZN => n64785);
   U50807 : NOR4_X1 port map( A1 => n64797, A2 => n64798, A3 => n64799, A4 => 
                           n64800, ZN => n64786);
   U50808 : NAND4_X1 port map( A1 => n64764, A2 => n64765, A3 => n64766, A4 => 
                           n64767, ZN => n5405);
   U50809 : AOI221_X1 port map( B1 => n67477, B2 => n57659, C1 => n67471, C2 =>
                           n59044, A => n64782, ZN => n64764);
   U50810 : AOI221_X1 port map( B1 => n67501, B2 => n66328, C1 => n67495, C2 =>
                           n58141, A => n64781, ZN => n64765);
   U50811 : NOR4_X1 port map( A1 => n64777, A2 => n64778, A3 => n64779, A4 => 
                           n64780, ZN => n64766);
   U50812 : NAND4_X1 port map( A1 => n64744, A2 => n64745, A3 => n64746, A4 => 
                           n64747, ZN => n5407);
   U50813 : AOI221_X1 port map( B1 => n67477, B2 => n57635, C1 => n67471, C2 =>
                           n59045, A => n64762, ZN => n64744);
   U50814 : AOI221_X1 port map( B1 => n67501, B2 => n66329, C1 => n67495, C2 =>
                           n58143, A => n64761, ZN => n64745);
   U50815 : NOR4_X1 port map( A1 => n64757, A2 => n64758, A3 => n64759, A4 => 
                           n64760, ZN => n64746);
   U50816 : NAND4_X1 port map( A1 => n64724, A2 => n64725, A3 => n64726, A4 => 
                           n64727, ZN => n5409);
   U50817 : AOI221_X1 port map( B1 => n67477, B2 => n57611, C1 => n67471, C2 =>
                           n59046, A => n64742, ZN => n64724);
   U50818 : AOI221_X1 port map( B1 => n67501, B2 => n66330, C1 => n67495, C2 =>
                           n58145, A => n64741, ZN => n64725);
   U50819 : NOR4_X1 port map( A1 => n64737, A2 => n64738, A3 => n64739, A4 => 
                           n64740, ZN => n64726);
   U50820 : NAND4_X1 port map( A1 => n64704, A2 => n64705, A3 => n64706, A4 => 
                           n64707, ZN => n5411);
   U50821 : AOI221_X1 port map( B1 => n67477, B2 => n57587, C1 => n67471, C2 =>
                           n59047, A => n64722, ZN => n64704);
   U50822 : AOI221_X1 port map( B1 => n67501, B2 => n66331, C1 => n67495, C2 =>
                           n58147, A => n64721, ZN => n64705);
   U50823 : NOR4_X1 port map( A1 => n64717, A2 => n64718, A3 => n64719, A4 => 
                           n64720, ZN => n64706);
   U50824 : NAND4_X1 port map( A1 => n64684, A2 => n64685, A3 => n64686, A4 => 
                           n64687, ZN => n5413);
   U50825 : AOI221_X1 port map( B1 => n67477, B2 => n57563, C1 => n67471, C2 =>
                           n59048, A => n64702, ZN => n64684);
   U50826 : AOI221_X1 port map( B1 => n67501, B2 => n66332, C1 => n67495, C2 =>
                           n58149, A => n64701, ZN => n64685);
   U50827 : NOR4_X1 port map( A1 => n64697, A2 => n64698, A3 => n64699, A4 => 
                           n64700, ZN => n64686);
   U50828 : NAND4_X1 port map( A1 => n64664, A2 => n64665, A3 => n64666, A4 => 
                           n64667, ZN => n5415);
   U50829 : AOI221_X1 port map( B1 => n67477, B2 => n57539, C1 => n67471, C2 =>
                           n59049, A => n64682, ZN => n64664);
   U50830 : AOI221_X1 port map( B1 => n67501, B2 => n66333, C1 => n67495, C2 =>
                           n58151, A => n64681, ZN => n64665);
   U50831 : NOR4_X1 port map( A1 => n64677, A2 => n64678, A3 => n64679, A4 => 
                           n64680, ZN => n64666);
   U50832 : NAND4_X1 port map( A1 => n64644, A2 => n64645, A3 => n64646, A4 => 
                           n64647, ZN => n5417);
   U50833 : AOI221_X1 port map( B1 => n67477, B2 => n57515, C1 => n67471, C2 =>
                           n59050, A => n64662, ZN => n64644);
   U50834 : AOI221_X1 port map( B1 => n67501, B2 => n66334, C1 => n67495, C2 =>
                           n58153, A => n64661, ZN => n64645);
   U50835 : NOR4_X1 port map( A1 => n64657, A2 => n64658, A3 => n64659, A4 => 
                           n64660, ZN => n64646);
   U50836 : NAND4_X1 port map( A1 => n64624, A2 => n64625, A3 => n64626, A4 => 
                           n64627, ZN => n5419);
   U50837 : AOI221_X1 port map( B1 => n67477, B2 => n57491, C1 => n67471, C2 =>
                           n59051, A => n64642, ZN => n64624);
   U50838 : AOI221_X1 port map( B1 => n67501, B2 => n66335, C1 => n67495, C2 =>
                           n58155, A => n64641, ZN => n64625);
   U50839 : NOR4_X1 port map( A1 => n64637, A2 => n64638, A3 => n64639, A4 => 
                           n64640, ZN => n64626);
   U50840 : NAND4_X1 port map( A1 => n64604, A2 => n64605, A3 => n64606, A4 => 
                           n64607, ZN => n5421);
   U50841 : AOI221_X1 port map( B1 => n67477, B2 => n57467, C1 => n67471, C2 =>
                           n59052, A => n64622, ZN => n64604);
   U50842 : AOI221_X1 port map( B1 => n67501, B2 => n66336, C1 => n67495, C2 =>
                           n58157, A => n64621, ZN => n64605);
   U50843 : NOR4_X1 port map( A1 => n64617, A2 => n64618, A3 => n64619, A4 => 
                           n64620, ZN => n64606);
   U50844 : NAND4_X1 port map( A1 => n64584, A2 => n64585, A3 => n64586, A4 => 
                           n64587, ZN => n5423);
   U50845 : AOI221_X1 port map( B1 => n67478, B2 => n57443, C1 => n67472, C2 =>
                           n59053, A => n64602, ZN => n64584);
   U50846 : AOI221_X1 port map( B1 => n67502, B2 => n66337, C1 => n67496, C2 =>
                           n58159, A => n64601, ZN => n64585);
   U50847 : NOR4_X1 port map( A1 => n64597, A2 => n64598, A3 => n64599, A4 => 
                           n64600, ZN => n64586);
   U50848 : NAND4_X1 port map( A1 => n64564, A2 => n64565, A3 => n64566, A4 => 
                           n64567, ZN => n5425);
   U50849 : AOI221_X1 port map( B1 => n67478, B2 => n57419, C1 => n67472, C2 =>
                           n59054, A => n64582, ZN => n64564);
   U50850 : AOI221_X1 port map( B1 => n67502, B2 => n66338, C1 => n67496, C2 =>
                           n58161, A => n64581, ZN => n64565);
   U50851 : NOR4_X1 port map( A1 => n64577, A2 => n64578, A3 => n64579, A4 => 
                           n64580, ZN => n64566);
   U50852 : NAND4_X1 port map( A1 => n64544, A2 => n64545, A3 => n64546, A4 => 
                           n64547, ZN => n5427);
   U50853 : AOI221_X1 port map( B1 => n67478, B2 => n57395, C1 => n67472, C2 =>
                           n59055, A => n64562, ZN => n64544);
   U50854 : AOI221_X1 port map( B1 => n67502, B2 => n66339, C1 => n67496, C2 =>
                           n58163, A => n64561, ZN => n64545);
   U50855 : NOR4_X1 port map( A1 => n64557, A2 => n64558, A3 => n64559, A4 => 
                           n64560, ZN => n64546);
   U50856 : NAND4_X1 port map( A1 => n64524, A2 => n64525, A3 => n64526, A4 => 
                           n64527, ZN => n5429);
   U50857 : AOI221_X1 port map( B1 => n67478, B2 => n57371, C1 => n67472, C2 =>
                           n59056, A => n64542, ZN => n64524);
   U50858 : AOI221_X1 port map( B1 => n67502, B2 => n66340, C1 => n67496, C2 =>
                           n58165, A => n64541, ZN => n64525);
   U50859 : NOR4_X1 port map( A1 => n64537, A2 => n64538, A3 => n64539, A4 => 
                           n64540, ZN => n64526);
   U50860 : NAND4_X1 port map( A1 => n64504, A2 => n64505, A3 => n64506, A4 => 
                           n64507, ZN => n5431);
   U50861 : AOI221_X1 port map( B1 => n67478, B2 => n57347, C1 => n67472, C2 =>
                           n59057, A => n64522, ZN => n64504);
   U50862 : AOI221_X1 port map( B1 => n67502, B2 => n66341, C1 => n67496, C2 =>
                           n58167, A => n64521, ZN => n64505);
   U50863 : NOR4_X1 port map( A1 => n64517, A2 => n64518, A3 => n64519, A4 => 
                           n64520, ZN => n64506);
   U50864 : NAND4_X1 port map( A1 => n64484, A2 => n64485, A3 => n64486, A4 => 
                           n64487, ZN => n5433);
   U50865 : AOI221_X1 port map( B1 => n67478, B2 => n57323, C1 => n67472, C2 =>
                           n59058, A => n64502, ZN => n64484);
   U50866 : AOI221_X1 port map( B1 => n67502, B2 => n66342, C1 => n67496, C2 =>
                           n58169, A => n64501, ZN => n64485);
   U50867 : NOR4_X1 port map( A1 => n64497, A2 => n64498, A3 => n64499, A4 => 
                           n64500, ZN => n64486);
   U50868 : NAND4_X1 port map( A1 => n64464, A2 => n64465, A3 => n64466, A4 => 
                           n64467, ZN => n5435);
   U50869 : AOI221_X1 port map( B1 => n67478, B2 => n57299, C1 => n67472, C2 =>
                           n59059, A => n64482, ZN => n64464);
   U50870 : AOI221_X1 port map( B1 => n67502, B2 => n66343, C1 => n67496, C2 =>
                           n58171, A => n64481, ZN => n64465);
   U50871 : NOR4_X1 port map( A1 => n64477, A2 => n64478, A3 => n64479, A4 => 
                           n64480, ZN => n64466);
   U50872 : NAND4_X1 port map( A1 => n64444, A2 => n64445, A3 => n64446, A4 => 
                           n64447, ZN => n5437);
   U50873 : AOI221_X1 port map( B1 => n67478, B2 => n57275, C1 => n67472, C2 =>
                           n59060, A => n64462, ZN => n64444);
   U50874 : AOI221_X1 port map( B1 => n67502, B2 => n66344, C1 => n67496, C2 =>
                           n58173, A => n64461, ZN => n64445);
   U50875 : NOR4_X1 port map( A1 => n64457, A2 => n64458, A3 => n64459, A4 => 
                           n64460, ZN => n64446);
   U50876 : NAND4_X1 port map( A1 => n64424, A2 => n64425, A3 => n64426, A4 => 
                           n64427, ZN => n5439);
   U50877 : AOI221_X1 port map( B1 => n67478, B2 => n57251, C1 => n67472, C2 =>
                           n59061, A => n64442, ZN => n64424);
   U50878 : AOI221_X1 port map( B1 => n67502, B2 => n66345, C1 => n67496, C2 =>
                           n58175, A => n64441, ZN => n64425);
   U50879 : NOR4_X1 port map( A1 => n64437, A2 => n64438, A3 => n64439, A4 => 
                           n64440, ZN => n64426);
   U50880 : NAND4_X1 port map( A1 => n64404, A2 => n64405, A3 => n64406, A4 => 
                           n64407, ZN => n5441);
   U50881 : AOI221_X1 port map( B1 => n67478, B2 => n57227, C1 => n67472, C2 =>
                           n59062, A => n64422, ZN => n64404);
   U50882 : AOI221_X1 port map( B1 => n67502, B2 => n66346, C1 => n67496, C2 =>
                           n58177, A => n64421, ZN => n64405);
   U50883 : NOR4_X1 port map( A1 => n64417, A2 => n64418, A3 => n64419, A4 => 
                           n64420, ZN => n64406);
   U50884 : NAND4_X1 port map( A1 => n64384, A2 => n64385, A3 => n64386, A4 => 
                           n64387, ZN => n5443);
   U50885 : AOI221_X1 port map( B1 => n67478, B2 => n57203, C1 => n67472, C2 =>
                           n59063, A => n64402, ZN => n64384);
   U50886 : AOI221_X1 port map( B1 => n67502, B2 => n66347, C1 => n67496, C2 =>
                           n58179, A => n64401, ZN => n64385);
   U50887 : NOR4_X1 port map( A1 => n64397, A2 => n64398, A3 => n64399, A4 => 
                           n64400, ZN => n64386);
   U50888 : NAND4_X1 port map( A1 => n64364, A2 => n64365, A3 => n64366, A4 => 
                           n64367, ZN => n5445);
   U50889 : AOI221_X1 port map( B1 => n67478, B2 => n57179, C1 => n67472, C2 =>
                           n59064, A => n64382, ZN => n64364);
   U50890 : AOI221_X1 port map( B1 => n67502, B2 => n66348, C1 => n67496, C2 =>
                           n58181, A => n64381, ZN => n64365);
   U50891 : NOR4_X1 port map( A1 => n64377, A2 => n64378, A3 => n64379, A4 => 
                           n64380, ZN => n64366);
   U50892 : NAND4_X1 port map( A1 => n64344, A2 => n64345, A3 => n64346, A4 => 
                           n64347, ZN => n5447);
   U50893 : AOI221_X1 port map( B1 => n67479, B2 => n57155, C1 => n67473, C2 =>
                           n59065, A => n64362, ZN => n64344);
   U50894 : AOI221_X1 port map( B1 => n67503, B2 => n66349, C1 => n67497, C2 =>
                           n58183, A => n64361, ZN => n64345);
   U50895 : NOR4_X1 port map( A1 => n64357, A2 => n64358, A3 => n64359, A4 => 
                           n64360, ZN => n64346);
   U50896 : NAND4_X1 port map( A1 => n64324, A2 => n64325, A3 => n64326, A4 => 
                           n64327, ZN => n5449);
   U50897 : AOI221_X1 port map( B1 => n67479, B2 => n57131, C1 => n67473, C2 =>
                           n59066, A => n64342, ZN => n64324);
   U50898 : AOI221_X1 port map( B1 => n67503, B2 => n66350, C1 => n67497, C2 =>
                           n58185, A => n64341, ZN => n64325);
   U50899 : NOR4_X1 port map( A1 => n64337, A2 => n64338, A3 => n64339, A4 => 
                           n64340, ZN => n64326);
   U50900 : NAND4_X1 port map( A1 => n64304, A2 => n64305, A3 => n64306, A4 => 
                           n64307, ZN => n5451);
   U50901 : AOI221_X1 port map( B1 => n67479, B2 => n57107, C1 => n67473, C2 =>
                           n59067, A => n64322, ZN => n64304);
   U50902 : AOI221_X1 port map( B1 => n67503, B2 => n66351, C1 => n67497, C2 =>
                           n58187, A => n64321, ZN => n64305);
   U50903 : NOR4_X1 port map( A1 => n64317, A2 => n64318, A3 => n64319, A4 => 
                           n64320, ZN => n64306);
   U50904 : NAND4_X1 port map( A1 => n64284, A2 => n64285, A3 => n64286, A4 => 
                           n64287, ZN => n5453);
   U50905 : AOI221_X1 port map( B1 => n67479, B2 => n57083, C1 => n67473, C2 =>
                           n59068, A => n64302, ZN => n64284);
   U50906 : AOI221_X1 port map( B1 => n67503, B2 => n66352, C1 => n67497, C2 =>
                           n58189, A => n64301, ZN => n64285);
   U50907 : NOR4_X1 port map( A1 => n64297, A2 => n64298, A3 => n64299, A4 => 
                           n64300, ZN => n64286);
   U50908 : NAND4_X1 port map( A1 => n64264, A2 => n64265, A3 => n64266, A4 => 
                           n64267, ZN => n5455);
   U50909 : AOI221_X1 port map( B1 => n67479, B2 => n57059, C1 => n67473, C2 =>
                           n59069, A => n64282, ZN => n64264);
   U50910 : AOI221_X1 port map( B1 => n67503, B2 => n66353, C1 => n67497, C2 =>
                           n58191, A => n64281, ZN => n64265);
   U50911 : NOR4_X1 port map( A1 => n64277, A2 => n64278, A3 => n64279, A4 => 
                           n64280, ZN => n64266);
   U50912 : NAND4_X1 port map( A1 => n64244, A2 => n64245, A3 => n64246, A4 => 
                           n64247, ZN => n5457);
   U50913 : AOI221_X1 port map( B1 => n67479, B2 => n57035, C1 => n67473, C2 =>
                           n59070, A => n64262, ZN => n64244);
   U50914 : AOI221_X1 port map( B1 => n67503, B2 => n66354, C1 => n67497, C2 =>
                           n58193, A => n64261, ZN => n64245);
   U50915 : NOR4_X1 port map( A1 => n64257, A2 => n64258, A3 => n64259, A4 => 
                           n64260, ZN => n64246);
   U50916 : NAND4_X1 port map( A1 => n64224, A2 => n64225, A3 => n64226, A4 => 
                           n64227, ZN => n5459);
   U50917 : AOI221_X1 port map( B1 => n67479, B2 => n57011, C1 => n67473, C2 =>
                           n59071, A => n64242, ZN => n64224);
   U50918 : AOI221_X1 port map( B1 => n67503, B2 => n66355, C1 => n67497, C2 =>
                           n58195, A => n64241, ZN => n64225);
   U50919 : NOR4_X1 port map( A1 => n64237, A2 => n64238, A3 => n64239, A4 => 
                           n64240, ZN => n64226);
   U50920 : NAND4_X1 port map( A1 => n64204, A2 => n64205, A3 => n64206, A4 => 
                           n64207, ZN => n5461);
   U50921 : AOI221_X1 port map( B1 => n67479, B2 => n56987, C1 => n67473, C2 =>
                           n59072, A => n64222, ZN => n64204);
   U50922 : AOI221_X1 port map( B1 => n67503, B2 => n66356, C1 => n67497, C2 =>
                           n58197, A => n64221, ZN => n64205);
   U50923 : NOR4_X1 port map( A1 => n64217, A2 => n64218, A3 => n64219, A4 => 
                           n64220, ZN => n64206);
   U50924 : NAND4_X1 port map( A1 => n64184, A2 => n64185, A3 => n64186, A4 => 
                           n64187, ZN => n5463);
   U50925 : AOI221_X1 port map( B1 => n67479, B2 => n56963, C1 => n67473, C2 =>
                           n59073, A => n64202, ZN => n64184);
   U50926 : AOI221_X1 port map( B1 => n67503, B2 => n66357, C1 => n67497, C2 =>
                           n58199, A => n64201, ZN => n64185);
   U50927 : NOR4_X1 port map( A1 => n64197, A2 => n64198, A3 => n64199, A4 => 
                           n64200, ZN => n64186);
   U50928 : NAND4_X1 port map( A1 => n64164, A2 => n64165, A3 => n64166, A4 => 
                           n64167, ZN => n5465);
   U50929 : AOI221_X1 port map( B1 => n67479, B2 => n56939, C1 => n67473, C2 =>
                           n59074, A => n64182, ZN => n64164);
   U50930 : AOI221_X1 port map( B1 => n67503, B2 => n66358, C1 => n67497, C2 =>
                           n58201, A => n64181, ZN => n64165);
   U50931 : NOR4_X1 port map( A1 => n64177, A2 => n64178, A3 => n64179, A4 => 
                           n64180, ZN => n64166);
   U50932 : NAND4_X1 port map( A1 => n64144, A2 => n64145, A3 => n64146, A4 => 
                           n64147, ZN => n5467);
   U50933 : AOI221_X1 port map( B1 => n67479, B2 => n56915, C1 => n67473, C2 =>
                           n59075, A => n64162, ZN => n64144);
   U50934 : AOI221_X1 port map( B1 => n67503, B2 => n66359, C1 => n67497, C2 =>
                           n58203, A => n64161, ZN => n64145);
   U50935 : NOR4_X1 port map( A1 => n64157, A2 => n64158, A3 => n64159, A4 => 
                           n64160, ZN => n64146);
   U50936 : NAND4_X1 port map( A1 => n64124, A2 => n64125, A3 => n64126, A4 => 
                           n64127, ZN => n5469);
   U50937 : AOI221_X1 port map( B1 => n67479, B2 => n56891, C1 => n67473, C2 =>
                           n59076, A => n64142, ZN => n64124);
   U50938 : AOI221_X1 port map( B1 => n67503, B2 => n66360, C1 => n67497, C2 =>
                           n58205, A => n64141, ZN => n64125);
   U50939 : NOR4_X1 port map( A1 => n64137, A2 => n64138, A3 => n64139, A4 => 
                           n64140, ZN => n64126);
   U50940 : NAND4_X1 port map( A1 => n64104, A2 => n64105, A3 => n64106, A4 => 
                           n64107, ZN => n5471);
   U50941 : AOI221_X1 port map( B1 => n67480, B2 => n56867, C1 => n67474, C2 =>
                           n59077, A => n64122, ZN => n64104);
   U50942 : AOI221_X1 port map( B1 => n67504, B2 => n66361, C1 => n67498, C2 =>
                           n58207, A => n64121, ZN => n64105);
   U50943 : NOR4_X1 port map( A1 => n64117, A2 => n64118, A3 => n64119, A4 => 
                           n64120, ZN => n64106);
   U50944 : NAND4_X1 port map( A1 => n64084, A2 => n64085, A3 => n64086, A4 => 
                           n64087, ZN => n5473);
   U50945 : AOI221_X1 port map( B1 => n67480, B2 => n56843, C1 => n67474, C2 =>
                           n59078, A => n64102, ZN => n64084);
   U50946 : AOI221_X1 port map( B1 => n67504, B2 => n66362, C1 => n67498, C2 =>
                           n58209, A => n64101, ZN => n64085);
   U50947 : NOR4_X1 port map( A1 => n64097, A2 => n64098, A3 => n64099, A4 => 
                           n64100, ZN => n64086);
   U50948 : NAND4_X1 port map( A1 => n64064, A2 => n64065, A3 => n64066, A4 => 
                           n64067, ZN => n5475);
   U50949 : AOI221_X1 port map( B1 => n67480, B2 => n56819, C1 => n67474, C2 =>
                           n59079, A => n64082, ZN => n64064);
   U50950 : AOI221_X1 port map( B1 => n67504, B2 => n66363, C1 => n67498, C2 =>
                           n58211, A => n64081, ZN => n64065);
   U50951 : NOR4_X1 port map( A1 => n64077, A2 => n64078, A3 => n64079, A4 => 
                           n64080, ZN => n64066);
   U50952 : NAND4_X1 port map( A1 => n64044, A2 => n64045, A3 => n64046, A4 => 
                           n64047, ZN => n5477);
   U50953 : AOI221_X1 port map( B1 => n67480, B2 => n56795, C1 => n67474, C2 =>
                           n59080, A => n64062, ZN => n64044);
   U50954 : AOI221_X1 port map( B1 => n67504, B2 => n66364, C1 => n67498, C2 =>
                           n58213, A => n64061, ZN => n64045);
   U50955 : NOR4_X1 port map( A1 => n64057, A2 => n64058, A3 => n64059, A4 => 
                           n64060, ZN => n64046);
   U50956 : NAND4_X1 port map( A1 => n64024, A2 => n64025, A3 => n64026, A4 => 
                           n64027, ZN => n5479);
   U50957 : AOI221_X1 port map( B1 => n67480, B2 => n56771, C1 => n67474, C2 =>
                           n59081, A => n64042, ZN => n64024);
   U50958 : AOI221_X1 port map( B1 => n67504, B2 => n66365, C1 => n67498, C2 =>
                           n58215, A => n64041, ZN => n64025);
   U50959 : NOR4_X1 port map( A1 => n64037, A2 => n64038, A3 => n64039, A4 => 
                           n64040, ZN => n64026);
   U50960 : NAND4_X1 port map( A1 => n64004, A2 => n64005, A3 => n64006, A4 => 
                           n64007, ZN => n5481);
   U50961 : AOI221_X1 port map( B1 => n67480, B2 => n56747, C1 => n67474, C2 =>
                           n59082, A => n64022, ZN => n64004);
   U50962 : AOI221_X1 port map( B1 => n67504, B2 => n66366, C1 => n67498, C2 =>
                           n58217, A => n64021, ZN => n64005);
   U50963 : NOR4_X1 port map( A1 => n64017, A2 => n64018, A3 => n64019, A4 => 
                           n64020, ZN => n64006);
   U50964 : NAND4_X1 port map( A1 => n63984, A2 => n63985, A3 => n63986, A4 => 
                           n63987, ZN => n5483);
   U50965 : AOI221_X1 port map( B1 => n67480, B2 => n56723, C1 => n67474, C2 =>
                           n59083, A => n64002, ZN => n63984);
   U50966 : AOI221_X1 port map( B1 => n67504, B2 => n66367, C1 => n67498, C2 =>
                           n58219, A => n64001, ZN => n63985);
   U50967 : NOR4_X1 port map( A1 => n63997, A2 => n63998, A3 => n63999, A4 => 
                           n64000, ZN => n63986);
   U50968 : NAND4_X1 port map( A1 => n63964, A2 => n63965, A3 => n63966, A4 => 
                           n63967, ZN => n5485);
   U50969 : AOI221_X1 port map( B1 => n67480, B2 => n56699, C1 => n67474, C2 =>
                           n59084, A => n63982, ZN => n63964);
   U50970 : AOI221_X1 port map( B1 => n67504, B2 => n66368, C1 => n67498, C2 =>
                           n58221, A => n63981, ZN => n63965);
   U50971 : NOR4_X1 port map( A1 => n63977, A2 => n63978, A3 => n63979, A4 => 
                           n63980, ZN => n63966);
   U50972 : NAND4_X1 port map( A1 => n63944, A2 => n63945, A3 => n63946, A4 => 
                           n63947, ZN => n5487);
   U50973 : AOI221_X1 port map( B1 => n67480, B2 => n56675, C1 => n67474, C2 =>
                           n59085, A => n63962, ZN => n63944);
   U50974 : AOI221_X1 port map( B1 => n67504, B2 => n66369, C1 => n67498, C2 =>
                           n58223, A => n63961, ZN => n63945);
   U50975 : NOR4_X1 port map( A1 => n63957, A2 => n63958, A3 => n63959, A4 => 
                           n63960, ZN => n63946);
   U50976 : NAND4_X1 port map( A1 => n63924, A2 => n63925, A3 => n63926, A4 => 
                           n63927, ZN => n5489);
   U50977 : AOI221_X1 port map( B1 => n67480, B2 => n56651, C1 => n67474, C2 =>
                           n59086, A => n63942, ZN => n63924);
   U50978 : AOI221_X1 port map( B1 => n67504, B2 => n66370, C1 => n67498, C2 =>
                           n58225, A => n63941, ZN => n63925);
   U50979 : NOR4_X1 port map( A1 => n63937, A2 => n63938, A3 => n63939, A4 => 
                           n63940, ZN => n63926);
   U50980 : NAND4_X1 port map( A1 => n63904, A2 => n63905, A3 => n63906, A4 => 
                           n63907, ZN => n5491);
   U50981 : AOI221_X1 port map( B1 => n67480, B2 => n56627, C1 => n67474, C2 =>
                           n59087, A => n63922, ZN => n63904);
   U50982 : AOI221_X1 port map( B1 => n67504, B2 => n66371, C1 => n67498, C2 =>
                           n58227, A => n63921, ZN => n63905);
   U50983 : NOR4_X1 port map( A1 => n63917, A2 => n63918, A3 => n63919, A4 => 
                           n63920, ZN => n63906);
   U50984 : NAND4_X1 port map( A1 => n63884, A2 => n63885, A3 => n63886, A4 => 
                           n63887, ZN => n5493);
   U50985 : AOI221_X1 port map( B1 => n67480, B2 => n56603, C1 => n67474, C2 =>
                           n59088, A => n63902, ZN => n63884);
   U50986 : AOI221_X1 port map( B1 => n67504, B2 => n66372, C1 => n67498, C2 =>
                           n58229, A => n63901, ZN => n63885);
   U50987 : NOR4_X1 port map( A1 => n63897, A2 => n63898, A3 => n63899, A4 => 
                           n63900, ZN => n63886);
   U50988 : NAND4_X1 port map( A1 => n63863, A2 => n63864, A3 => n63865, A4 => 
                           n63866, ZN => n5495);
   U50989 : AOI221_X1 port map( B1 => n67481, B2 => n56579, C1 => n67475, C2 =>
                           n59089, A => n63882, ZN => n63863);
   U50990 : AOI221_X1 port map( B1 => n67505, B2 => n66305, C1 => n67499, C2 =>
                           n58231, A => n63881, ZN => n63864);
   U50991 : NOR4_X1 port map( A1 => n63867, A2 => n63868, A3 => n63869, A4 => 
                           n63870, ZN => n63866);
   U50992 : NAND4_X1 port map( A1 => n63842, A2 => n63843, A3 => n63844, A4 => 
                           n63845, ZN => n5497);
   U50993 : AOI221_X1 port map( B1 => n67481, B2 => n56555, C1 => n67475, C2 =>
                           n59090, A => n63861, ZN => n63842);
   U50994 : AOI221_X1 port map( B1 => n67505, B2 => n66306, C1 => n67499, C2 =>
                           n58232, A => n63860, ZN => n63843);
   U50995 : NOR4_X1 port map( A1 => n63846, A2 => n63847, A3 => n63848, A4 => 
                           n63849, ZN => n63845);
   U50996 : NAND4_X1 port map( A1 => n63821, A2 => n63822, A3 => n63823, A4 => 
                           n63824, ZN => n5499);
   U50997 : AOI221_X1 port map( B1 => n67481, B2 => n56531, C1 => n67475, C2 =>
                           n59091, A => n63840, ZN => n63821);
   U50998 : AOI221_X1 port map( B1 => n67505, B2 => n66307, C1 => n67499, C2 =>
                           n58233, A => n63839, ZN => n63822);
   U50999 : NOR4_X1 port map( A1 => n63825, A2 => n63826, A3 => n63827, A4 => 
                           n63828, ZN => n63824);
   U51000 : NAND4_X1 port map( A1 => n63767, A2 => n63768, A3 => n63769, A4 => 
                           n63770, ZN => n5501);
   U51001 : AOI221_X1 port map( B1 => n67481, B2 => n56490, C1 => n67475, C2 =>
                           n59092, A => n63817, ZN => n63767);
   U51002 : AOI221_X1 port map( B1 => n67505, B2 => n66308, C1 => n67499, C2 =>
                           n58234, A => n63812, ZN => n63768);
   U51003 : NOR4_X1 port map( A1 => n63771, A2 => n63772, A3 => n63773, A4 => 
                           n63774, ZN => n63770);
   U51004 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n63295);
   U51005 : INV_X1 port map( A => RESET, ZN => n62087);
   U51006 : INV_X1 port map( A => DATAIN(60), ZN => n61966);
   U51007 : INV_X1 port map( A => DATAIN(61), ZN => n61964);
   U51008 : INV_X1 port map( A => DATAIN(62), ZN => n61962);
   U51009 : INV_X1 port map( A => DATAIN(63), ZN => n61960);
   U51010 : INV_X1 port map( A => DATAIN(0), ZN => n62086);
   U51011 : INV_X1 port map( A => DATAIN(1), ZN => n62084);
   U51012 : INV_X1 port map( A => DATAIN(2), ZN => n62082);
   U51013 : INV_X1 port map( A => DATAIN(3), ZN => n62080);
   U51014 : INV_X1 port map( A => DATAIN(4), ZN => n62078);
   U51015 : INV_X1 port map( A => DATAIN(5), ZN => n62076);
   U51016 : INV_X1 port map( A => DATAIN(6), ZN => n62074);
   U51017 : INV_X1 port map( A => DATAIN(7), ZN => n62072);
   U51018 : INV_X1 port map( A => DATAIN(8), ZN => n62070);
   U51019 : INV_X1 port map( A => DATAIN(9), ZN => n62068);
   U51020 : INV_X1 port map( A => DATAIN(10), ZN => n62066);
   U51021 : INV_X1 port map( A => DATAIN(11), ZN => n62064);
   U51022 : INV_X1 port map( A => DATAIN(12), ZN => n62062);
   U51023 : INV_X1 port map( A => DATAIN(13), ZN => n62060);
   U51024 : INV_X1 port map( A => DATAIN(14), ZN => n62058);
   U51025 : INV_X1 port map( A => DATAIN(15), ZN => n62056);
   U51026 : INV_X1 port map( A => DATAIN(16), ZN => n62054);
   U51027 : INV_X1 port map( A => DATAIN(17), ZN => n62052);
   U51028 : INV_X1 port map( A => DATAIN(18), ZN => n62050);
   U51029 : INV_X1 port map( A => DATAIN(19), ZN => n62048);
   U51030 : INV_X1 port map( A => DATAIN(20), ZN => n62046);
   U51031 : INV_X1 port map( A => DATAIN(21), ZN => n62044);
   U51032 : INV_X1 port map( A => DATAIN(22), ZN => n62042);
   U51033 : INV_X1 port map( A => DATAIN(23), ZN => n62040);
   U51034 : INV_X1 port map( A => DATAIN(24), ZN => n62038);
   U51035 : INV_X1 port map( A => DATAIN(25), ZN => n62036);
   U51036 : INV_X1 port map( A => DATAIN(26), ZN => n62034);
   U51037 : INV_X1 port map( A => DATAIN(27), ZN => n62032);
   U51038 : INV_X1 port map( A => DATAIN(28), ZN => n62030);
   U51039 : INV_X1 port map( A => DATAIN(29), ZN => n62028);
   U51040 : INV_X1 port map( A => DATAIN(30), ZN => n62026);
   U51041 : INV_X1 port map( A => DATAIN(31), ZN => n62024);
   U51042 : INV_X1 port map( A => DATAIN(32), ZN => n62022);
   U51043 : INV_X1 port map( A => DATAIN(33), ZN => n62020);
   U51044 : INV_X1 port map( A => DATAIN(34), ZN => n62018);
   U51045 : INV_X1 port map( A => DATAIN(35), ZN => n62016);
   U51046 : INV_X1 port map( A => DATAIN(36), ZN => n62014);
   U51047 : INV_X1 port map( A => DATAIN(37), ZN => n62012);
   U51048 : INV_X1 port map( A => DATAIN(38), ZN => n62010);
   U51049 : INV_X1 port map( A => DATAIN(39), ZN => n62008);
   U51050 : INV_X1 port map( A => DATAIN(40), ZN => n62006);
   U51051 : INV_X1 port map( A => DATAIN(41), ZN => n62004);
   U51052 : INV_X1 port map( A => DATAIN(42), ZN => n62002);
   U51053 : INV_X1 port map( A => DATAIN(43), ZN => n62000);
   U51054 : INV_X1 port map( A => DATAIN(44), ZN => n61998);
   U51055 : INV_X1 port map( A => DATAIN(45), ZN => n61996);
   U51056 : INV_X1 port map( A => DATAIN(46), ZN => n61994);
   U51057 : INV_X1 port map( A => DATAIN(47), ZN => n61992);
   U51058 : INV_X1 port map( A => DATAIN(48), ZN => n61990);
   U51059 : INV_X1 port map( A => DATAIN(49), ZN => n61988);
   U51060 : INV_X1 port map( A => DATAIN(50), ZN => n61986);
   U51061 : INV_X1 port map( A => DATAIN(51), ZN => n61984);
   U51062 : INV_X1 port map( A => DATAIN(52), ZN => n61982);
   U51063 : INV_X1 port map( A => DATAIN(53), ZN => n61980);
   U51064 : INV_X1 port map( A => DATAIN(54), ZN => n61978);
   U51065 : INV_X1 port map( A => DATAIN(55), ZN => n61976);
   U51066 : INV_X1 port map( A => DATAIN(56), ZN => n61974);
   U51067 : INV_X1 port map( A => DATAIN(57), ZN => n61972);
   U51068 : INV_X1 port map( A => DATAIN(58), ZN => n61970);
   U51069 : INV_X1 port map( A => DATAIN(59), ZN => n61968);
   U51070 : INV_X1 port map( A => ADD_WR(3), ZN => n62491);
   U51071 : INV_X1 port map( A => ADD_WR(0), ZN => n62490);
   U51072 : INV_X1 port map( A => ADD_WR(1), ZN => n63497);
   U51073 : INV_X1 port map( A => ADD_RD2(2), ZN => n66299);
   U51074 : INV_X1 port map( A => ADD_RD2(1), ZN => n66301);
   U51075 : INV_X1 port map( A => ADD_WR(2), ZN => n63496);
   U51076 : INV_X1 port map( A => ADD_RD1(2), ZN => n65099);
   U51077 : AND3_X1 port map( A1 => ENABLE, A2 => n62958, A3 => WR, ZN => 
                           n62492);
   U51078 : INV_X1 port map( A => ADD_WR(4), ZN => n62958);
   U51079 : CLKBUF_X1 port map( A => n65150, Z => n67265);
   U51080 : CLKBUF_X1 port map( A => n65149, Z => n67271);
   U51081 : CLKBUF_X1 port map( A => n65147, Z => n67277);
   U51082 : CLKBUF_X1 port map( A => n65146, Z => n67283);
   U51083 : CLKBUF_X1 port map( A => n65145, Z => n67289);
   U51084 : CLKBUF_X1 port map( A => n65144, Z => n67295);
   U51085 : CLKBUF_X1 port map( A => n65142, Z => n67301);
   U51086 : CLKBUF_X1 port map( A => n65141, Z => n67307);
   U51087 : CLKBUF_X1 port map( A => n65140, Z => n67313);
   U51088 : CLKBUF_X1 port map( A => n65139, Z => n67319);
   U51089 : CLKBUF_X1 port map( A => n65138, Z => n67325);
   U51090 : CLKBUF_X1 port map( A => n65137, Z => n67331);
   U51091 : CLKBUF_X1 port map( A => n65136, Z => n67337);
   U51092 : CLKBUF_X1 port map( A => n65135, Z => n67343);
   U51093 : CLKBUF_X1 port map( A => n65134, Z => n67349);
   U51094 : CLKBUF_X1 port map( A => n65133, Z => n67355);
   U51095 : CLKBUF_X1 port map( A => n65132, Z => n67361);
   U51096 : CLKBUF_X1 port map( A => n65127, Z => n67367);
   U51097 : CLKBUF_X1 port map( A => n65126, Z => n67373);
   U51098 : CLKBUF_X1 port map( A => n65124, Z => n67379);
   U51099 : CLKBUF_X1 port map( A => n65123, Z => n67385);
   U51100 : CLKBUF_X1 port map( A => n65122, Z => n67391);
   U51101 : CLKBUF_X1 port map( A => n65121, Z => n67397);
   U51102 : CLKBUF_X1 port map( A => n65119, Z => n67403);
   U51103 : CLKBUF_X1 port map( A => n65118, Z => n67409);
   U51104 : CLKBUF_X1 port map( A => n65117, Z => n67415);
   U51105 : CLKBUF_X1 port map( A => n65116, Z => n67421);
   U51106 : CLKBUF_X1 port map( A => n65114, Z => n67427);
   U51107 : CLKBUF_X1 port map( A => n65113, Z => n67433);
   U51108 : CLKBUF_X1 port map( A => n65112, Z => n67439);
   U51109 : CLKBUF_X1 port map( A => n65111, Z => n67445);
   U51110 : CLKBUF_X1 port map( A => n65109, Z => n67451);
   U51111 : CLKBUF_X1 port map( A => n65108, Z => n67457);
   U51112 : CLKBUF_X1 port map( A => n63819, Z => n67463);
   U51113 : CLKBUF_X1 port map( A => n63818, Z => n67469);
   U51114 : CLKBUF_X1 port map( A => n63816, Z => n67475);
   U51115 : CLKBUF_X1 port map( A => n63815, Z => n67481);
   U51116 : CLKBUF_X1 port map( A => n63814, Z => n67487);
   U51117 : CLKBUF_X1 port map( A => n63813, Z => n67493);
   U51118 : CLKBUF_X1 port map( A => n63811, Z => n67499);
   U51119 : CLKBUF_X1 port map( A => n63810, Z => n67505);
   U51120 : CLKBUF_X1 port map( A => n63809, Z => n67511);
   U51121 : CLKBUF_X1 port map( A => n63808, Z => n67517);
   U51122 : CLKBUF_X1 port map( A => n63807, Z => n67523);
   U51123 : CLKBUF_X1 port map( A => n63806, Z => n67529);
   U51124 : CLKBUF_X1 port map( A => n63805, Z => n67535);
   U51125 : CLKBUF_X1 port map( A => n63804, Z => n67541);
   U51126 : CLKBUF_X1 port map( A => n63803, Z => n67547);
   U51127 : CLKBUF_X1 port map( A => n63802, Z => n67553);
   U51128 : CLKBUF_X1 port map( A => n63801, Z => n67559);
   U51129 : CLKBUF_X1 port map( A => n63795, Z => n67565);
   U51130 : CLKBUF_X1 port map( A => n63794, Z => n67571);
   U51131 : CLKBUF_X1 port map( A => n63792, Z => n67577);
   U51132 : CLKBUF_X1 port map( A => n63791, Z => n67583);
   U51133 : CLKBUF_X1 port map( A => n63790, Z => n67589);
   U51134 : CLKBUF_X1 port map( A => n63788, Z => n67595);
   U51135 : CLKBUF_X1 port map( A => n63786, Z => n67601);
   U51136 : CLKBUF_X1 port map( A => n63785, Z => n67607);
   U51137 : CLKBUF_X1 port map( A => n63784, Z => n67613);
   U51138 : CLKBUF_X1 port map( A => n63783, Z => n67619);
   U51139 : CLKBUF_X1 port map( A => n63781, Z => n67625);
   U51140 : CLKBUF_X1 port map( A => n63780, Z => n67631);
   U51141 : CLKBUF_X1 port map( A => n63778, Z => n67641);
   U51142 : CLKBUF_X1 port map( A => n63776, Z => n67647);
   U51143 : CLKBUF_X1 port map( A => n63775, Z => n67653);
   U51144 : CLKBUF_X1 port map( A => n63766, Z => n67659);
   U51145 : CLKBUF_X1 port map( A => n63700, Z => n67672);
   U51146 : CLKBUF_X1 port map( A => n63634, Z => n67685);
   U51147 : CLKBUF_X1 port map( A => n63568, Z => n67698);
   U51148 : CLKBUF_X1 port map( A => n63502, Z => n67711);
   U51149 : CLKBUF_X1 port map( A => n63499, Z => n67724);
   U51150 : CLKBUF_X1 port map( A => n63498, Z => n67730);
   U51151 : CLKBUF_X1 port map( A => n63431, Z => n67736);
   U51152 : CLKBUF_X1 port map( A => n63364, Z => n67749);
   U51153 : CLKBUF_X1 port map( A => n63298, Z => n67762);
   U51154 : CLKBUF_X1 port map( A => n63231, Z => n67775);
   U51155 : CLKBUF_X1 port map( A => n63228, Z => n67788);
   U51156 : CLKBUF_X1 port map( A => n63227, Z => n67794);
   U51157 : CLKBUF_X1 port map( A => n63163, Z => n67800);
   U51158 : CLKBUF_X1 port map( A => n63097, Z => n67813);
   U51159 : CLKBUF_X1 port map( A => n63094, Z => n67826);
   U51160 : CLKBUF_X1 port map( A => n63093, Z => n67832);
   U51161 : CLKBUF_X1 port map( A => n63028, Z => n67838);
   U51162 : CLKBUF_X1 port map( A => n62961, Z => n67851);
   U51163 : CLKBUF_X1 port map( A => n62894, Z => n67864);
   U51164 : CLKBUF_X1 port map( A => n62828, Z => n67877);
   U51165 : CLKBUF_X1 port map( A => n62765, Z => n67890);
   U51166 : CLKBUF_X1 port map( A => n62763, Z => n67903);
   U51167 : CLKBUF_X1 port map( A => n62762, Z => n67909);
   U51168 : CLKBUF_X1 port map( A => n62698, Z => n67915);
   U51169 : CLKBUF_X1 port map( A => n62695, Z => n67928);
   U51170 : CLKBUF_X1 port map( A => n62693, Z => n67934);
   U51171 : CLKBUF_X1 port map( A => n62628, Z => n67940);
   U51172 : CLKBUF_X1 port map( A => n62561, Z => n67953);
   U51173 : CLKBUF_X1 port map( A => n62495, Z => n67966);
   U51174 : CLKBUF_X1 port map( A => n62425, Z => n67979);
   U51175 : CLKBUF_X1 port map( A => n62359, Z => n67992);
   U51176 : CLKBUF_X1 port map( A => n62292, Z => n68005);
   U51177 : CLKBUF_X1 port map( A => n62226, Z => n68018);
   U51178 : CLKBUF_X1 port map( A => n62159, Z => n68031);
   U51179 : CLKBUF_X1 port map( A => n62092, Z => n68044);
   U51180 : CLKBUF_X1 port map( A => n62087, Z => n68057);
   U51181 : CLKBUF_X1 port map( A => n61959, Z => n68255);

end SYN_A;
